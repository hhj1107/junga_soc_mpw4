magic
tech sky130A
magscale 1 2
timestamp 1640332777
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 215938 700680 215944 700732
rect 215996 700720 216002 700732
rect 235166 700720 235172 700732
rect 215996 700692 235172 700720
rect 215996 700680 216002 700692
rect 235166 700680 235172 700692
rect 235224 700680 235230 700732
rect 209038 700612 209044 700664
rect 209096 700652 209102 700664
rect 267642 700652 267648 700664
rect 209096 700624 267648 700652
rect 209096 700612 209102 700624
rect 267642 700612 267648 700624
rect 267700 700612 267706 700664
rect 206370 700544 206376 700596
rect 206428 700584 206434 700596
rect 283834 700584 283840 700596
rect 206428 700556 283840 700584
rect 206428 700544 206434 700556
rect 283834 700544 283840 700556
rect 283892 700544 283898 700596
rect 385678 700544 385684 700596
rect 385736 700584 385742 700596
rect 397454 700584 397460 700596
rect 385736 700556 397460 700584
rect 385736 700544 385742 700556
rect 397454 700544 397460 700556
rect 397512 700544 397518 700596
rect 399478 700544 399484 700596
rect 399536 700584 399542 700596
rect 478506 700584 478512 700596
rect 399536 700556 478512 700584
rect 399536 700544 399542 700556
rect 478506 700544 478512 700556
rect 478564 700544 478570 700596
rect 206278 700476 206284 700528
rect 206336 700516 206342 700528
rect 300118 700516 300124 700528
rect 206336 700488 300124 700516
rect 206336 700476 206342 700488
rect 300118 700476 300124 700488
rect 300176 700476 300182 700528
rect 382918 700476 382924 700528
rect 382976 700516 382982 700528
rect 462314 700516 462320 700528
rect 382976 700488 462320 700516
rect 382976 700476 382982 700488
rect 462314 700476 462320 700488
rect 462372 700476 462378 700528
rect 204898 700408 204904 700460
rect 204956 700448 204962 700460
rect 332502 700448 332508 700460
rect 204956 700420 332508 700448
rect 204956 700408 204962 700420
rect 332502 700408 332508 700420
rect 332560 700408 332566 700460
rect 370498 700408 370504 700460
rect 370556 700448 370562 700460
rect 494790 700448 494796 700460
rect 370556 700420 494796 700448
rect 370556 700408 370562 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 170306 700340 170312 700392
rect 170364 700380 170370 700392
rect 196526 700380 196532 700392
rect 170364 700352 196532 700380
rect 170364 700340 170370 700352
rect 196526 700340 196532 700352
rect 196584 700340 196590 700392
rect 213178 700340 213184 700392
rect 213236 700380 213242 700392
rect 348786 700380 348792 700392
rect 213236 700352 348792 700380
rect 213236 700340 213242 700352
rect 348786 700340 348792 700352
rect 348844 700340 348850 700392
rect 381538 700340 381544 700392
rect 381596 700380 381602 700392
rect 527174 700380 527180 700392
rect 381596 700352 527180 700380
rect 381596 700340 381602 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 33778 700312 33784 700324
rect 24360 700284 33784 700312
rect 24360 700272 24366 700284
rect 33778 700272 33784 700284
rect 33836 700272 33842 700324
rect 58894 700272 58900 700324
rect 58952 700312 58958 700324
rect 72970 700312 72976 700324
rect 58952 700284 72976 700312
rect 58952 700272 58958 700284
rect 72970 700272 72976 700284
rect 73028 700272 73034 700324
rect 154114 700272 154120 700324
rect 154172 700312 154178 700324
rect 196618 700312 196624 700324
rect 154172 700284 196624 700312
rect 154172 700272 154178 700284
rect 196618 700272 196624 700284
rect 196676 700272 196682 700324
rect 197998 700272 198004 700324
rect 198056 700312 198062 700324
rect 364978 700312 364984 700324
rect 198056 700284 364984 700312
rect 198056 700272 198062 700284
rect 364978 700272 364984 700284
rect 365036 700272 365042 700324
rect 367738 700272 367744 700324
rect 367796 700312 367802 700324
rect 559650 700312 559656 700324
rect 367796 700284 559656 700312
rect 367796 700272 367802 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 88334 699660 88340 699712
rect 88392 699700 88398 699712
rect 89162 699700 89168 699712
rect 88392 699672 89168 699700
rect 88392 699660 88398 699672
rect 89162 699660 89168 699672
rect 89220 699660 89226 699712
rect 104894 699660 104900 699712
rect 104952 699700 104958 699712
rect 105446 699700 105452 699712
rect 104952 699672 105452 699700
rect 104952 699660 104958 699672
rect 105446 699660 105452 699672
rect 105504 699660 105510 699712
rect 210418 699660 210424 699712
rect 210476 699700 210482 699712
rect 218974 699700 218980 699712
rect 210476 699672 218980 699700
rect 210476 699660 210482 699672
rect 218974 699660 218980 699672
rect 219032 699660 219038 699712
rect 134150 698572 134156 698624
rect 134208 698612 134214 698624
rect 137830 698612 137836 698624
rect 134208 698584 137836 698612
rect 134208 698572 134214 698584
rect 137830 698572 137836 698584
rect 137888 698572 137894 698624
rect 134150 696980 134156 696992
rect 132466 696952 134156 696980
rect 128906 696872 128912 696924
rect 128964 696912 128970 696924
rect 132466 696912 132494 696952
rect 134150 696940 134156 696952
rect 134208 696940 134214 696992
rect 378778 696940 378784 696992
rect 378836 696980 378842 696992
rect 580166 696980 580172 696992
rect 378836 696952 580172 696980
rect 378836 696940 378842 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 128964 696884 132494 696912
rect 128964 696872 128970 696884
rect 126514 693744 126520 693796
rect 126572 693784 126578 693796
rect 128906 693784 128912 693796
rect 126572 693756 128912 693784
rect 126572 693744 126578 693756
rect 128906 693744 128912 693756
rect 128964 693744 128970 693796
rect 124582 690140 124588 690192
rect 124640 690180 124646 690192
rect 126514 690180 126520 690192
rect 124640 690152 126520 690180
rect 124640 690140 124646 690152
rect 126514 690140 126520 690152
rect 126572 690140 126578 690192
rect 121454 688644 121460 688696
rect 121512 688684 121518 688696
rect 124582 688684 124588 688696
rect 121512 688656 124588 688684
rect 121512 688644 121518 688656
rect 124582 688644 124588 688656
rect 124640 688644 124646 688696
rect 114554 684360 114560 684412
rect 114612 684400 114618 684412
rect 121454 684400 121460 684412
rect 114612 684372 121460 684400
rect 114612 684360 114618 684372
rect 121454 684360 121460 684372
rect 121512 684360 121518 684412
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 396718 683136 396724 683188
rect 396776 683176 396782 683188
rect 580166 683176 580172 683188
rect 396776 683148 580172 683176
rect 396776 683136 396782 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 114554 681748 114560 681760
rect 113146 681720 114560 681748
rect 106274 681640 106280 681692
rect 106332 681680 106338 681692
rect 113146 681680 113174 681720
rect 114554 681708 114560 681720
rect 114612 681708 114618 681760
rect 106332 681652 113174 681680
rect 106332 681640 106338 681652
rect 104250 674704 104256 674756
rect 104308 674744 104314 674756
rect 106182 674744 106188 674756
rect 104308 674716 106188 674744
rect 104308 674704 104314 674716
rect 106182 674704 106188 674716
rect 106240 674704 106246 674756
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 35158 670732 35164 670744
rect 3568 670704 35164 670732
rect 3568 670692 3574 670704
rect 35158 670692 35164 670704
rect 35216 670692 35222 670744
rect 363598 670692 363604 670744
rect 363656 670732 363662 670744
rect 580166 670732 580172 670744
rect 363656 670704 580172 670732
rect 363656 670692 363662 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 102778 667360 102784 667412
rect 102836 667400 102842 667412
rect 104250 667400 104256 667412
rect 102836 667372 104256 667400
rect 102836 667360 102842 667372
rect 104250 667360 104256 667372
rect 104308 667360 104314 667412
rect 100754 662396 100760 662448
rect 100812 662436 100818 662448
rect 102778 662436 102784 662448
rect 100812 662408 102784 662436
rect 100812 662396 100818 662408
rect 102778 662396 102784 662408
rect 102836 662396 102842 662448
rect 100754 659716 100760 659728
rect 96632 659688 100760 659716
rect 96522 659608 96528 659660
rect 96580 659648 96586 659660
rect 96632 659648 96660 659688
rect 100754 659676 100760 659688
rect 100812 659676 100818 659728
rect 96580 659620 96660 659648
rect 96580 659608 96586 659620
rect 94498 657976 94504 658028
rect 94556 658016 94562 658028
rect 96522 658016 96528 658028
rect 94556 657988 96528 658016
rect 94556 657976 94562 657988
rect 96522 657976 96528 657988
rect 96580 657976 96586 658028
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 21358 656928 21364 656940
rect 3476 656900 21364 656928
rect 3476 656888 3482 656900
rect 21358 656888 21364 656900
rect 21416 656888 21422 656940
rect 92474 650088 92480 650140
rect 92532 650128 92538 650140
rect 94498 650128 94504 650140
rect 92532 650100 94504 650128
rect 92532 650088 92538 650100
rect 94498 650088 94504 650100
rect 94556 650088 94562 650140
rect 77202 647844 77208 647896
rect 77260 647884 77266 647896
rect 92474 647884 92480 647896
rect 77260 647856 92480 647884
rect 77260 647844 77266 647856
rect 92474 647844 92480 647856
rect 92532 647844 92538 647896
rect 74534 645872 74540 645924
rect 74592 645912 74598 645924
rect 77202 645912 77208 645924
rect 74592 645884 77208 645912
rect 74592 645872 74598 645884
rect 77202 645872 77208 645884
rect 77260 645872 77266 645924
rect 377398 643084 377404 643136
rect 377456 643124 377462 643136
rect 580166 643124 580172 643136
rect 377456 643096 580172 643124
rect 377456 643084 377462 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 74534 638976 74540 638988
rect 74506 638936 74540 638976
rect 74592 638936 74598 638988
rect 71774 638868 71780 638920
rect 71832 638908 71838 638920
rect 74506 638908 74534 638936
rect 71832 638880 74534 638908
rect 71832 638868 71838 638880
rect 71774 636256 71780 636268
rect 70412 636228 71780 636256
rect 69014 636148 69020 636200
rect 69072 636188 69078 636200
rect 70412 636188 70440 636228
rect 71774 636216 71780 636228
rect 71832 636216 71838 636268
rect 69072 636160 70440 636188
rect 69072 636148 69078 636160
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 11698 632108 11704 632120
rect 3476 632080 11704 632108
rect 3476 632068 3482 632080
rect 11698 632068 11704 632080
rect 11756 632068 11762 632120
rect 69014 632108 69020 632120
rect 67652 632080 69020 632108
rect 65518 632000 65524 632052
rect 65576 632040 65582 632052
rect 67652 632040 67680 632080
rect 69014 632068 69020 632080
rect 69072 632068 69078 632120
rect 65576 632012 67680 632040
rect 65576 632000 65582 632012
rect 395338 630640 395344 630692
rect 395396 630680 395402 630692
rect 580166 630680 580172 630692
rect 395396 630652 580172 630680
rect 395396 630640 395402 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 36538 618304 36544 618316
rect 3200 618276 36544 618304
rect 3200 618264 3206 618276
rect 36538 618264 36544 618276
rect 36596 618264 36602 618316
rect 360838 616836 360844 616888
rect 360896 616876 360902 616888
rect 580166 616876 580172 616888
rect 360896 616848 580172 616876
rect 360896 616836 360902 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 22738 605860 22744 605872
rect 3292 605832 22744 605860
rect 3292 605820 3298 605832
rect 22738 605820 22744 605832
rect 22796 605820 22802 605872
rect 64138 604460 64144 604512
rect 64196 604500 64202 604512
rect 65518 604500 65524 604512
rect 64196 604472 65524 604500
rect 64196 604460 64202 604472
rect 65518 604460 65524 604472
rect 65576 604460 65582 604512
rect 558178 590656 558184 590708
rect 558236 590696 558242 590708
rect 579798 590696 579804 590708
rect 558236 590668 579804 590696
rect 558236 590656 558242 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 14458 579680 14464 579692
rect 3384 579652 14464 579680
rect 3384 579640 3390 579652
rect 14458 579640 14464 579652
rect 14516 579640 14522 579692
rect 393958 576852 393964 576904
rect 394016 576892 394022 576904
rect 580166 576892 580172 576904
rect 394016 576864 580172 576892
rect 394016 576852 394022 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 62758 572704 62764 572756
rect 62816 572744 62822 572756
rect 64138 572744 64144 572756
rect 62816 572716 64144 572744
rect 62816 572704 62822 572716
rect 64138 572704 64144 572716
rect 64196 572704 64202 572756
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 39298 565876 39304 565888
rect 3476 565848 39304 565876
rect 3476 565836 3482 565848
rect 39298 565836 39304 565848
rect 39356 565836 39362 565888
rect 358078 563048 358084 563100
rect 358136 563088 358142 563100
rect 579798 563088 579804 563100
rect 358136 563060 579804 563088
rect 358136 563048 358142 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 61378 561008 61384 561060
rect 61436 561048 61442 561060
rect 62758 561048 62764 561060
rect 61436 561020 62764 561048
rect 61436 561008 61442 561020
rect 62758 561008 62764 561020
rect 62816 561008 62822 561060
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 25498 553432 25504 553444
rect 3476 553404 25504 553432
rect 3476 553392 3482 553404
rect 25498 553392 25504 553404
rect 25556 553392 25562 553444
rect 59998 553392 60004 553444
rect 60056 553432 60062 553444
rect 61378 553432 61384 553444
rect 60056 553404 61384 553432
rect 60056 553392 60062 553404
rect 61378 553392 61384 553404
rect 61436 553392 61442 553444
rect 376018 536800 376024 536852
rect 376076 536840 376082 536852
rect 580166 536840 580172 536852
rect 376076 536812 580172 536840
rect 376076 536800 376082 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 15838 527184 15844 527196
rect 3476 527156 15844 527184
rect 3476 527144 3482 527156
rect 15838 527144 15844 527156
rect 15896 527144 15902 527196
rect 392578 524424 392584 524476
rect 392636 524464 392642 524476
rect 580166 524464 580172 524476
rect 392636 524436 580172 524464
rect 392636 524424 392642 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 43438 514808 43444 514820
rect 3476 514780 43444 514808
rect 3476 514768 3482 514780
rect 43438 514768 43444 514780
rect 43496 514768 43502 514820
rect 213362 510620 213368 510672
rect 213420 510660 213426 510672
rect 580166 510660 580172 510672
rect 213420 510632 580172 510660
rect 213420 510620 213426 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 29638 501004 29644 501016
rect 3108 500976 29644 501004
rect 3108 500964 3114 500976
rect 29638 500964 29644 500976
rect 29696 500964 29702 501016
rect 374638 484372 374644 484424
rect 374696 484412 374702 484424
rect 580166 484412 580172 484424
rect 374696 484384 580172 484412
rect 374696 484372 374702 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 17218 474756 17224 474768
rect 3476 474728 17224 474756
rect 3476 474716 3482 474728
rect 17218 474716 17224 474728
rect 17276 474716 17282 474768
rect 389818 470568 389824 470620
rect 389876 470608 389882 470620
rect 579982 470608 579988 470620
rect 389876 470580 579988 470608
rect 389876 470568 389882 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 47578 462380 47584 462392
rect 3292 462352 47584 462380
rect 3292 462340 3298 462352
rect 47578 462340 47584 462352
rect 47636 462340 47642 462392
rect 425698 456764 425704 456816
rect 425756 456804 425762 456816
rect 580166 456804 580172 456816
rect 425756 456776 580172 456804
rect 425756 456764 425762 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 32398 448576 32404 448588
rect 3200 448548 32404 448576
rect 3200 448536 3206 448548
rect 32398 448536 32404 448548
rect 32456 448536 32462 448588
rect 209222 430584 209228 430636
rect 209280 430624 209286 430636
rect 216674 430624 216680 430636
rect 209280 430596 216680 430624
rect 209280 430584 209286 430596
rect 216674 430584 216680 430596
rect 216732 430584 216738 430636
rect 388438 430584 388444 430636
rect 388496 430624 388502 430636
rect 580166 430624 580172 430636
rect 388496 430596 580172 430624
rect 388496 430584 388502 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 18598 422328 18604 422340
rect 3476 422300 18604 422328
rect 3476 422288 3482 422300
rect 18598 422288 18604 422300
rect 18656 422288 18662 422340
rect 214558 408348 214564 408400
rect 214616 408388 214622 408400
rect 216674 408388 216680 408400
rect 214616 408360 216680 408388
rect 214616 408348 214622 408360
rect 216674 408348 216680 408360
rect 216732 408348 216738 408400
rect 371878 404336 371884 404388
rect 371936 404376 371942 404388
rect 580166 404376 580172 404388
rect 371936 404348 580172 404376
rect 371936 404336 371942 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 218606 400052 218612 400104
rect 218664 400092 218670 400104
rect 218664 400064 226748 400092
rect 218664 400052 218670 400064
rect 226720 400036 226748 400064
rect 218146 399984 218152 400036
rect 218204 400024 218210 400036
rect 226334 400024 226340 400036
rect 218204 399996 226340 400024
rect 218204 399984 218210 399996
rect 226334 399984 226340 399996
rect 226392 399984 226398 400036
rect 226702 399984 226708 400036
rect 226760 399984 226766 400036
rect 218238 399916 218244 399968
rect 218296 399956 218302 399968
rect 226518 399956 226524 399968
rect 218296 399928 226524 399956
rect 218296 399916 218302 399928
rect 226518 399916 226524 399928
rect 226576 399916 226582 399968
rect 217594 399848 217600 399900
rect 217652 399888 217658 399900
rect 231854 399888 231860 399900
rect 217652 399860 231860 399888
rect 217652 399848 217658 399860
rect 231854 399848 231860 399860
rect 231912 399848 231918 399900
rect 58894 399780 58900 399832
rect 58952 399820 58958 399832
rect 121454 399820 121460 399832
rect 58952 399792 121460 399820
rect 58952 399780 58958 399792
rect 121454 399780 121460 399792
rect 121512 399780 121518 399832
rect 177942 399780 177948 399832
rect 178000 399820 178006 399832
rect 209222 399820 209228 399832
rect 178000 399792 209228 399820
rect 178000 399780 178006 399792
rect 209222 399780 209228 399792
rect 209280 399780 209286 399832
rect 217686 399780 217692 399832
rect 217744 399820 217750 399832
rect 232130 399820 232136 399832
rect 217744 399792 232136 399820
rect 217744 399780 217750 399792
rect 232130 399780 232136 399792
rect 232188 399780 232194 399832
rect 111702 399712 111708 399764
rect 111760 399752 111766 399764
rect 204898 399752 204904 399764
rect 111760 399724 204904 399752
rect 111760 399712 111766 399724
rect 204898 399712 204904 399724
rect 204956 399712 204962 399764
rect 217410 399712 217416 399764
rect 217468 399752 217474 399764
rect 233234 399752 233240 399764
rect 217468 399724 233240 399752
rect 217468 399712 217474 399724
rect 233234 399712 233240 399724
rect 233292 399712 233298 399764
rect 57054 399644 57060 399696
rect 57112 399684 57118 399696
rect 230750 399684 230756 399696
rect 57112 399656 230756 399684
rect 57112 399644 57118 399656
rect 230750 399644 230756 399656
rect 230808 399644 230814 399696
rect 57238 399576 57244 399628
rect 57296 399616 57302 399628
rect 232038 399616 232044 399628
rect 57296 399588 232044 399616
rect 57296 399576 57302 399588
rect 232038 399576 232044 399588
rect 232096 399576 232102 399628
rect 57146 399508 57152 399560
rect 57204 399548 57210 399560
rect 231946 399548 231952 399560
rect 57204 399520 231952 399548
rect 57204 399508 57210 399520
rect 231946 399508 231952 399520
rect 232004 399508 232010 399560
rect 244918 399508 244924 399560
rect 244976 399548 244982 399560
rect 358998 399548 359004 399560
rect 244976 399520 359004 399548
rect 244976 399508 244982 399520
rect 358998 399508 359004 399520
rect 359056 399508 359062 399560
rect 57330 399440 57336 399492
rect 57388 399480 57394 399492
rect 232222 399480 232228 399492
rect 57388 399452 232228 399480
rect 57388 399440 57394 399452
rect 232222 399440 232228 399452
rect 232280 399440 232286 399492
rect 242250 399440 242256 399492
rect 242308 399480 242314 399492
rect 359090 399480 359096 399492
rect 242308 399452 359096 399480
rect 242308 399440 242314 399452
rect 359090 399440 359096 399452
rect 359148 399440 359154 399492
rect 218422 399372 218428 399424
rect 218480 399412 218486 399424
rect 226426 399412 226432 399424
rect 218480 399384 226432 399412
rect 218480 399372 218486 399384
rect 226426 399372 226432 399384
rect 226484 399372 226490 399424
rect 59998 398828 60004 398880
rect 60056 398868 60062 398880
rect 62022 398868 62028 398880
rect 60056 398840 62028 398868
rect 60056 398828 60062 398840
rect 62022 398828 62028 398840
rect 62080 398828 62086 398880
rect 59354 398760 59360 398812
rect 59412 398800 59418 398812
rect 214558 398800 214564 398812
rect 59412 398772 214564 398800
rect 59412 398760 59418 398772
rect 214558 398760 214564 398772
rect 214616 398760 214622 398812
rect 219526 398692 219532 398744
rect 219584 398732 219590 398744
rect 224954 398732 224960 398744
rect 219584 398704 224960 398732
rect 219584 398692 219590 398704
rect 224954 398692 224960 398704
rect 225012 398692 225018 398744
rect 219618 398556 219624 398608
rect 219676 398596 219682 398608
rect 225230 398596 225236 398608
rect 219676 398568 225236 398596
rect 219676 398556 219682 398568
rect 225230 398556 225236 398568
rect 225288 398556 225294 398608
rect 219894 398488 219900 398540
rect 219952 398528 219958 398540
rect 226610 398528 226616 398540
rect 219952 398500 226616 398528
rect 219952 398488 219958 398500
rect 226610 398488 226616 398500
rect 226668 398488 226674 398540
rect 121362 398216 121368 398268
rect 121420 398256 121426 398268
rect 196618 398256 196624 398268
rect 121420 398228 196624 398256
rect 121420 398216 121426 398228
rect 196618 398216 196624 398228
rect 196676 398216 196682 398268
rect 225138 398256 225144 398268
rect 219406 398228 225144 398256
rect 115842 398148 115848 398200
rect 115900 398188 115906 398200
rect 206370 398188 206376 398200
rect 115900 398160 206376 398188
rect 115900 398148 115906 398160
rect 206370 398148 206376 398160
rect 206428 398148 206434 398200
rect 218054 398148 218060 398200
rect 218112 398188 218118 398200
rect 219406 398188 219434 398228
rect 225138 398216 225144 398228
rect 225196 398216 225202 398268
rect 218112 398160 219434 398188
rect 218112 398148 218118 398160
rect 219710 398148 219716 398200
rect 219768 398188 219774 398200
rect 225046 398188 225052 398200
rect 219768 398160 225052 398188
rect 219768 398148 219774 398160
rect 225046 398148 225052 398160
rect 225104 398148 225110 398200
rect 57882 398080 57888 398132
rect 57940 398120 57946 398132
rect 165614 398120 165620 398132
rect 57940 398092 165620 398120
rect 57940 398080 57946 398092
rect 165614 398080 165620 398092
rect 165672 398080 165678 398132
rect 217502 398080 217508 398132
rect 217560 398120 217566 398132
rect 232314 398120 232320 398132
rect 217560 398092 232320 398120
rect 217560 398080 217566 398092
rect 232314 398080 232320 398092
rect 232372 398080 232378 398132
rect 3510 397468 3516 397520
rect 3568 397508 3574 397520
rect 140774 397508 140780 397520
rect 3568 397480 140780 397508
rect 3568 397468 3574 397480
rect 140774 397468 140780 397480
rect 140832 397468 140838 397520
rect 216582 397332 216588 397384
rect 216640 397372 216646 397384
rect 275278 397372 275284 397384
rect 216640 397344 275284 397372
rect 216640 397332 216646 397344
rect 275278 397332 275284 397344
rect 275336 397332 275342 397384
rect 85482 397264 85488 397316
rect 85540 397304 85546 397316
rect 230566 397304 230572 397316
rect 85540 397276 230572 397304
rect 85540 397264 85546 397276
rect 230566 397264 230572 397276
rect 230624 397264 230630 397316
rect 304258 397264 304264 397316
rect 304316 397304 304322 397316
rect 308582 397304 308588 397316
rect 304316 397276 308588 397304
rect 304316 397264 304322 397276
rect 308582 397264 308588 397276
rect 308640 397264 308646 397316
rect 62942 397196 62948 397248
rect 63000 397236 63006 397248
rect 239214 397236 239220 397248
rect 63000 397208 239220 397236
rect 63000 397196 63006 397208
rect 239214 397196 239220 397208
rect 239272 397196 239278 397248
rect 79594 397128 79600 397180
rect 79652 397168 79658 397180
rect 230658 397168 230664 397180
rect 79652 397140 230664 397168
rect 79652 397128 79658 397140
rect 230658 397128 230664 397140
rect 230716 397128 230722 397180
rect 253290 397128 253296 397180
rect 253348 397168 253354 397180
rect 259454 397168 259460 397180
rect 253348 397140 259460 397168
rect 253348 397128 253354 397140
rect 259454 397128 259460 397140
rect 259512 397128 259518 397180
rect 89346 397060 89352 397112
rect 89404 397100 89410 397112
rect 94498 397100 94504 397112
rect 89404 397072 94504 397100
rect 89404 397060 89410 397072
rect 94498 397060 94504 397072
rect 94556 397060 94562 397112
rect 183462 397060 183468 397112
rect 183520 397100 183526 397112
rect 229278 397100 229284 397112
rect 183520 397072 229284 397100
rect 183520 397060 183526 397072
rect 229278 397060 229284 397072
rect 229336 397060 229342 397112
rect 62758 396992 62764 397044
rect 62816 397032 62822 397044
rect 113818 397032 113824 397044
rect 62816 397004 113824 397032
rect 62816 396992 62822 397004
rect 113818 396992 113824 397004
rect 113876 396992 113882 397044
rect 206922 396992 206928 397044
rect 206980 397032 206986 397044
rect 268654 397032 268660 397044
rect 206980 397004 268660 397032
rect 206980 396992 206986 397004
rect 268654 396992 268660 397004
rect 268712 396992 268718 397044
rect 61470 396924 61476 396976
rect 61528 396964 61534 396976
rect 109126 396964 109132 396976
rect 61528 396936 109132 396964
rect 61528 396924 61534 396936
rect 109126 396924 109132 396936
rect 109184 396924 109190 396976
rect 188338 396924 188344 396976
rect 188396 396964 188402 396976
rect 250070 396964 250076 396976
rect 188396 396936 250076 396964
rect 188396 396924 188402 396936
rect 250070 396924 250076 396936
rect 250128 396924 250134 396976
rect 82354 396856 82360 396908
rect 82412 396896 82418 396908
rect 162118 396896 162124 396908
rect 82412 396868 162124 396896
rect 82412 396856 82418 396868
rect 162118 396856 162124 396868
rect 162176 396856 162182 396908
rect 173158 396856 173164 396908
rect 173216 396896 173222 396908
rect 236178 396896 236184 396908
rect 173216 396868 236184 396896
rect 173216 396856 173222 396868
rect 236178 396856 236184 396868
rect 236236 396856 236242 396908
rect 78306 396788 78312 396840
rect 78364 396828 78370 396840
rect 168374 396828 168380 396840
rect 78364 396800 168380 396828
rect 78364 396788 78370 396800
rect 168374 396788 168380 396800
rect 168432 396788 168438 396840
rect 186958 396788 186964 396840
rect 187016 396828 187022 396840
rect 252738 396828 252744 396840
rect 187016 396800 252744 396828
rect 187016 396788 187022 396800
rect 252738 396788 252744 396800
rect 252796 396788 252802 396840
rect 113358 396720 113364 396772
rect 113416 396760 113422 396772
rect 230842 396760 230848 396772
rect 113416 396732 230848 396760
rect 113416 396720 113422 396732
rect 230842 396720 230848 396732
rect 230900 396720 230906 396772
rect 250438 396720 250444 396772
rect 250496 396760 250502 396772
rect 256878 396760 256884 396772
rect 250496 396732 256884 396760
rect 250496 396720 250502 396732
rect 256878 396720 256884 396732
rect 256936 396720 256942 396772
rect 262858 396720 262864 396772
rect 262916 396760 262922 396772
rect 265158 396760 265164 396772
rect 262916 396732 265164 396760
rect 262916 396720 262922 396732
rect 265158 396720 265164 396732
rect 265216 396720 265222 396772
rect 268470 396720 268476 396772
rect 268528 396760 268534 396772
rect 269390 396760 269396 396772
rect 268528 396732 269396 396760
rect 268528 396720 268534 396732
rect 269390 396720 269396 396732
rect 269448 396720 269454 396772
rect 282178 396720 282184 396772
rect 282236 396760 282242 396772
rect 283742 396760 283748 396772
rect 282236 396732 283748 396760
rect 282236 396720 282242 396732
rect 283742 396720 283748 396732
rect 283800 396720 283806 396772
rect 291838 396720 291844 396772
rect 291896 396760 291902 396772
rect 292666 396760 292672 396772
rect 291896 396732 292672 396760
rect 291896 396720 291902 396732
rect 292666 396720 292672 396732
rect 292724 396720 292730 396772
rect 112346 396652 112352 396704
rect 112404 396692 112410 396704
rect 230934 396692 230940 396704
rect 112404 396664 230940 396692
rect 112404 396652 112410 396664
rect 230934 396652 230940 396664
rect 230992 396652 230998 396704
rect 242158 396652 242164 396704
rect 242216 396692 242222 396704
rect 244550 396692 244556 396704
rect 242216 396664 244556 396692
rect 242216 396652 242222 396664
rect 244550 396652 244556 396664
rect 244608 396652 244614 396704
rect 249058 396652 249064 396704
rect 249116 396692 249122 396704
rect 251358 396692 251364 396704
rect 249116 396664 251364 396692
rect 249116 396652 249122 396664
rect 251358 396652 251364 396664
rect 251416 396652 251422 396704
rect 251910 396652 251916 396704
rect 251968 396692 251974 396704
rect 254118 396692 254124 396704
rect 251968 396664 254124 396692
rect 251968 396652 251974 396664
rect 254118 396652 254124 396664
rect 254176 396652 254182 396704
rect 268378 396652 268384 396704
rect 268436 396692 268442 396704
rect 273622 396692 273628 396704
rect 268436 396664 273628 396692
rect 268436 396652 268442 396664
rect 273622 396652 273628 396664
rect 273680 396652 273686 396704
rect 284938 396652 284944 396704
rect 284996 396692 285002 396704
rect 285950 396692 285956 396704
rect 284996 396664 285956 396692
rect 284996 396652 285002 396664
rect 285950 396652 285956 396664
rect 286008 396652 286014 396704
rect 58618 396584 58624 396636
rect 58676 396624 58682 396636
rect 95878 396624 95884 396636
rect 58676 396596 95884 396624
rect 58676 396584 58682 396596
rect 95878 396584 95884 396596
rect 95936 396584 95942 396636
rect 106918 396584 106924 396636
rect 106976 396624 106982 396636
rect 230474 396624 230480 396636
rect 106976 396596 230480 396624
rect 106976 396584 106982 396596
rect 230474 396584 230480 396596
rect 230532 396584 230538 396636
rect 61378 396516 61384 396568
rect 61436 396556 61442 396568
rect 98086 396556 98092 396568
rect 61436 396528 98092 396556
rect 61436 396516 61442 396528
rect 98086 396516 98092 396528
rect 98144 396516 98150 396568
rect 104802 396516 104808 396568
rect 104860 396556 104866 396568
rect 229370 396556 229376 396568
rect 104860 396528 229376 396556
rect 104860 396516 104866 396528
rect 229370 396516 229376 396528
rect 229428 396516 229434 396568
rect 95050 396448 95056 396500
rect 95108 396488 95114 396500
rect 229094 396488 229100 396500
rect 95108 396460 229100 396488
rect 95108 396448 95114 396460
rect 229094 396448 229100 396460
rect 229152 396448 229158 396500
rect 246298 396448 246304 396500
rect 246356 396488 246362 396500
rect 263594 396488 263600 396500
rect 246356 396460 263600 396488
rect 246356 396448 246362 396460
rect 263594 396448 263600 396460
rect 263652 396448 263658 396500
rect 90082 396380 90088 396432
rect 90140 396420 90146 396432
rect 227714 396420 227720 396432
rect 90140 396392 227720 396420
rect 90140 396380 90146 396392
rect 227714 396380 227720 396392
rect 227772 396380 227778 396432
rect 260098 396380 260104 396432
rect 260156 396420 260162 396432
rect 325878 396420 325884 396432
rect 260156 396392 325884 396420
rect 260156 396380 260162 396392
rect 325878 396380 325884 396392
rect 325936 396380 325942 396432
rect 59998 396312 60004 396364
rect 60056 396352 60062 396364
rect 76190 396352 76196 396364
rect 60056 396324 76196 396352
rect 60056 396312 60062 396324
rect 76190 396312 76196 396324
rect 76248 396312 76254 396364
rect 91462 396312 91468 396364
rect 91520 396352 91526 396364
rect 229186 396352 229192 396364
rect 91520 396324 229192 396352
rect 91520 396312 91526 396324
rect 229186 396312 229192 396324
rect 229244 396312 229250 396364
rect 235258 396312 235264 396364
rect 235316 396352 235322 396364
rect 272334 396352 272340 396364
rect 235316 396324 272340 396352
rect 235316 396312 235322 396324
rect 272334 396312 272340 396324
rect 272392 396312 272398 396364
rect 93486 396244 93492 396296
rect 93544 396284 93550 396296
rect 231026 396284 231032 396296
rect 93544 396256 231032 396284
rect 93544 396244 93550 396256
rect 231026 396244 231032 396256
rect 231084 396244 231090 396296
rect 233970 396244 233976 396296
rect 234028 396284 234034 396296
rect 247678 396284 247684 396296
rect 234028 396256 247684 396284
rect 234028 396244 234034 396256
rect 247678 396244 247684 396256
rect 247736 396244 247742 396296
rect 253198 396244 253204 396296
rect 253256 396284 253262 396296
rect 261938 396284 261944 396296
rect 253256 396256 261944 396284
rect 253256 396244 253262 396256
rect 261938 396244 261944 396256
rect 261996 396244 262002 396296
rect 269758 396244 269764 396296
rect 269816 396284 269822 396296
rect 315758 396284 315764 396296
rect 269816 396256 315764 396284
rect 269816 396244 269822 396256
rect 315758 396244 315764 396256
rect 315816 396244 315822 396296
rect 58894 396176 58900 396228
rect 58952 396216 58958 396228
rect 82998 396216 83004 396228
rect 58952 396188 83004 396216
rect 58952 396176 58958 396188
rect 82998 396176 83004 396188
rect 83056 396176 83062 396228
rect 222838 396176 222844 396228
rect 222896 396216 222902 396228
rect 277670 396216 277676 396228
rect 222896 396188 277676 396216
rect 222896 396176 222902 396188
rect 277670 396176 277676 396188
rect 277728 396176 277734 396228
rect 59906 396108 59912 396160
rect 59964 396148 59970 396160
rect 80422 396148 80428 396160
rect 59964 396120 80428 396148
rect 59964 396108 59970 396120
rect 80422 396108 80428 396120
rect 80480 396108 80486 396160
rect 106090 396108 106096 396160
rect 106148 396148 106154 396160
rect 115198 396148 115204 396160
rect 106148 396120 115204 396148
rect 106148 396108 106154 396120
rect 115198 396108 115204 396120
rect 115256 396108 115262 396160
rect 237466 396108 237472 396160
rect 237524 396148 237530 396160
rect 248598 396148 248604 396160
rect 237524 396120 248604 396148
rect 237524 396108 237530 396120
rect 248598 396108 248604 396120
rect 248656 396108 248662 396160
rect 255958 396108 255964 396160
rect 256016 396148 256022 396160
rect 260926 396148 260932 396160
rect 256016 396120 260932 396148
rect 256016 396108 256022 396120
rect 260926 396108 260932 396120
rect 260984 396108 260990 396160
rect 316678 396108 316684 396160
rect 316736 396148 316742 396160
rect 342622 396148 342628 396160
rect 316736 396120 342628 396148
rect 316736 396108 316742 396120
rect 342622 396108 342628 396120
rect 342680 396108 342686 396160
rect 102778 396040 102784 396092
rect 102836 396080 102842 396092
rect 106918 396080 106924 396092
rect 102836 396052 106924 396080
rect 102836 396040 102842 396052
rect 106918 396040 106924 396052
rect 106976 396040 106982 396092
rect 108850 396040 108856 396092
rect 108908 396080 108914 396092
rect 119338 396080 119344 396092
rect 108908 396052 119344 396080
rect 108908 396040 108914 396052
rect 119338 396040 119344 396052
rect 119396 396040 119402 396092
rect 163866 395972 163872 396024
rect 163924 396012 163930 396024
rect 219434 396012 219440 396024
rect 163924 395984 219440 396012
rect 163924 395972 163930 395984
rect 219434 395972 219440 395984
rect 219492 395972 219498 396024
rect 251818 395972 251824 396024
rect 251876 396012 251882 396024
rect 256142 396012 256148 396024
rect 251876 395984 256148 396012
rect 251876 395972 251882 395984
rect 256142 395972 256148 395984
rect 256200 395972 256206 396024
rect 118602 395904 118608 395956
rect 118660 395944 118666 395956
rect 189074 395944 189080 395956
rect 118660 395916 189080 395944
rect 118660 395904 118666 395916
rect 189074 395904 189080 395916
rect 189132 395904 189138 395956
rect 113634 395836 113640 395888
rect 113692 395876 113698 395888
rect 184934 395876 184940 395888
rect 113692 395848 184940 395876
rect 113692 395836 113698 395848
rect 184934 395836 184940 395848
rect 184992 395836 184998 395888
rect 195882 395836 195888 395888
rect 195940 395876 195946 395888
rect 262306 395876 262312 395888
rect 195940 395848 262312 395876
rect 195940 395836 195946 395848
rect 262306 395836 262312 395848
rect 262364 395836 262370 395888
rect 154114 395768 154120 395820
rect 154172 395808 154178 395820
rect 227990 395808 227996 395820
rect 154172 395780 227996 395808
rect 154172 395768 154178 395780
rect 227990 395768 227996 395780
rect 228048 395768 228054 395820
rect 171042 395700 171048 395752
rect 171100 395740 171106 395752
rect 250346 395740 250352 395752
rect 171100 395712 250352 395740
rect 171100 395700 171106 395712
rect 250346 395700 250352 395712
rect 250404 395700 250410 395752
rect 184842 395632 184848 395684
rect 184900 395672 184906 395684
rect 268286 395672 268292 395684
rect 184900 395644 268292 395672
rect 184900 395632 184906 395644
rect 268286 395632 268292 395644
rect 268344 395632 268350 395684
rect 136450 395564 136456 395616
rect 136508 395604 136514 395616
rect 227806 395604 227812 395616
rect 136508 395576 227812 395604
rect 136508 395564 136514 395576
rect 227806 395564 227812 395576
rect 227864 395564 227870 395616
rect 118234 395496 118240 395548
rect 118292 395536 118298 395548
rect 224862 395536 224868 395548
rect 118292 395508 224868 395536
rect 118292 395496 118298 395508
rect 224862 395496 224868 395508
rect 224920 395496 224926 395548
rect 233878 395496 233884 395548
rect 233936 395536 233942 395548
rect 247954 395536 247960 395548
rect 233936 395508 247960 395536
rect 233936 395496 233942 395508
rect 247954 395496 247960 395508
rect 248012 395496 248018 395548
rect 61562 395428 61568 395480
rect 61620 395468 61626 395480
rect 278866 395468 278872 395480
rect 61620 395440 278872 395468
rect 61620 395428 61626 395440
rect 278866 395428 278872 395440
rect 278924 395428 278930 395480
rect 56502 395360 56508 395412
rect 56560 395400 56566 395412
rect 290182 395400 290188 395412
rect 56560 395372 290188 395400
rect 56560 395360 56566 395372
rect 290182 395360 290188 395372
rect 290240 395360 290246 395412
rect 54570 395292 54576 395344
rect 54628 395332 54634 395344
rect 298462 395332 298468 395344
rect 54628 395304 298468 395332
rect 54628 395292 54634 395304
rect 298462 395292 298468 395304
rect 298520 395292 298526 395344
rect 62114 394680 62120 394732
rect 62172 394720 62178 394732
rect 62172 394692 64874 394720
rect 62172 394680 62178 394692
rect 64846 394652 64874 394692
rect 66254 394652 66260 394664
rect 64846 394624 66260 394652
rect 66254 394612 66260 394624
rect 66312 394612 66318 394664
rect 238018 394000 238024 394052
rect 238076 394040 238082 394052
rect 251174 394040 251180 394052
rect 238076 394012 251180 394040
rect 238076 394000 238082 394012
rect 251174 394000 251180 394012
rect 251232 394000 251238 394052
rect 177850 393932 177856 393984
rect 177908 393972 177914 393984
rect 237466 393972 237472 393984
rect 177908 393944 237472 393972
rect 177908 393932 177914 393944
rect 237466 393932 237472 393944
rect 237524 393932 237530 393984
rect 240778 392640 240784 392692
rect 240836 392680 240842 392692
rect 258166 392680 258172 392692
rect 240836 392652 258172 392680
rect 240836 392640 240842 392652
rect 258166 392640 258172 392652
rect 258224 392640 258230 392692
rect 193122 392572 193128 392624
rect 193180 392612 193186 392624
rect 253290 392612 253296 392624
rect 193180 392584 253296 392612
rect 193180 392572 193186 392584
rect 253290 392572 253296 392584
rect 253348 392572 253354 392624
rect 258718 392572 258724 392624
rect 258776 392612 258782 392624
rect 277486 392612 277492 392624
rect 258776 392584 277492 392612
rect 258776 392572 258782 392584
rect 277486 392572 277492 392584
rect 277544 392572 277550 392624
rect 66254 389172 66260 389224
rect 66312 389212 66318 389224
rect 68278 389212 68284 389224
rect 66312 389184 68284 389212
rect 66312 389172 66318 389184
rect 68278 389172 68284 389184
rect 68336 389172 68342 389224
rect 84102 378156 84108 378208
rect 84160 378196 84166 378208
rect 580166 378196 580172 378208
rect 84160 378168 580172 378196
rect 84160 378156 84166 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 68278 378088 68284 378140
rect 68336 378128 68342 378140
rect 69658 378128 69664 378140
rect 68336 378100 69664 378128
rect 68336 378088 68342 378100
rect 69658 378088 69664 378100
rect 69716 378088 69722 378140
rect 43438 373396 43444 373448
rect 43496 373436 43502 373448
rect 136634 373436 136640 373448
rect 43496 373408 136640 373436
rect 43496 373396 43502 373408
rect 136634 373396 136640 373408
rect 136692 373396 136698 373448
rect 39298 373328 39304 373380
rect 39356 373368 39362 373380
rect 133874 373368 133880 373380
rect 39356 373340 133880 373368
rect 39356 373328 39362 373340
rect 133874 373328 133880 373340
rect 133932 373328 133938 373380
rect 3418 373260 3424 373312
rect 3476 373300 3482 373312
rect 142154 373300 142160 373312
rect 3476 373272 142160 373300
rect 3476 373260 3482 373272
rect 142154 373260 142160 373272
rect 142212 373260 142218 373312
rect 195790 373260 195796 373312
rect 195848 373300 195854 373312
rect 287054 373300 287060 373312
rect 195848 373272 287060 373300
rect 195848 373260 195854 373272
rect 287054 373260 287060 373272
rect 287112 373260 287118 373312
rect 69658 372852 69664 372904
rect 69716 372892 69722 372904
rect 70394 372892 70400 372904
rect 69716 372864 70400 372892
rect 69716 372852 69722 372864
rect 70394 372852 70400 372864
rect 70452 372852 70458 372904
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 143534 371260 143540 371272
rect 3476 371232 143540 371260
rect 3476 371220 3482 371232
rect 143534 371220 143540 371232
rect 143592 371220 143598 371272
rect 70394 369792 70400 369844
rect 70452 369832 70458 369844
rect 75178 369832 75184 369844
rect 70452 369804 75184 369832
rect 70452 369792 70458 369804
rect 75178 369792 75184 369804
rect 75236 369792 75242 369844
rect 85482 364352 85488 364404
rect 85540 364392 85546 364404
rect 579614 364392 579620 364404
rect 85540 364364 579620 364392
rect 85540 364352 85546 364364
rect 579614 364352 579620 364364
rect 579672 364352 579678 364404
rect 75178 358708 75184 358760
rect 75236 358748 75242 358760
rect 76650 358748 76656 358760
rect 75236 358720 76656 358748
rect 75236 358708 75242 358720
rect 76650 358708 76656 358720
rect 76708 358708 76714 358760
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 144914 357456 144920 357468
rect 3200 357428 144920 357456
rect 3200 357416 3206 357428
rect 144914 357416 144920 357428
rect 144972 357416 144978 357468
rect 76650 357348 76656 357400
rect 76708 357388 76714 357400
rect 78030 357388 78036 357400
rect 76708 357360 78036 357388
rect 76708 357348 76714 357360
rect 78030 357348 78036 357360
rect 78088 357348 78094 357400
rect 56318 356668 56324 356720
rect 56376 356708 56382 356720
rect 145006 356708 145012 356720
rect 56376 356680 145012 356708
rect 56376 356668 56382 356680
rect 145006 356668 145012 356680
rect 145064 356668 145070 356720
rect 78030 353268 78036 353320
rect 78088 353308 78094 353320
rect 80698 353308 80704 353320
rect 78088 353280 80704 353308
rect 78088 353268 78094 353280
rect 80698 353268 80704 353280
rect 80756 353268 80762 353320
rect 82722 351908 82728 351960
rect 82780 351948 82786 351960
rect 580166 351948 580172 351960
rect 82780 351920 580172 351948
rect 82780 351908 82786 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 143626 345080 143632 345092
rect 3384 345052 143632 345080
rect 3384 345040 3390 345052
rect 143626 345040 143632 345052
rect 143684 345040 143690 345092
rect 80698 335996 80704 336048
rect 80756 336036 80762 336048
rect 84194 336036 84200 336048
rect 80756 336008 84200 336036
rect 80756 335996 80762 336008
rect 84194 335996 84200 336008
rect 84252 335996 84258 336048
rect 84194 329740 84200 329792
rect 84252 329780 84258 329792
rect 86218 329780 86224 329792
rect 84252 329752 86224 329780
rect 84252 329740 84258 329752
rect 86218 329740 86224 329752
rect 86276 329740 86282 329792
rect 86218 324572 86224 324624
rect 86276 324612 86282 324624
rect 87966 324612 87972 324624
rect 86276 324584 87972 324612
rect 86276 324572 86282 324584
rect 87966 324572 87972 324584
rect 88024 324572 88030 324624
rect 81342 324300 81348 324352
rect 81400 324340 81406 324352
rect 580166 324340 580172 324352
rect 81400 324312 580172 324340
rect 81400 324300 81406 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 87966 322940 87972 322992
rect 88024 322980 88030 322992
rect 88024 322952 89760 322980
rect 88024 322940 88030 322952
rect 89732 322912 89760 322952
rect 91738 322912 91744 322924
rect 89732 322884 91744 322912
rect 91738 322872 91744 322884
rect 91796 322872 91802 322924
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 146294 318832 146300 318844
rect 3476 318804 146300 318832
rect 3476 318792 3482 318804
rect 146294 318792 146300 318804
rect 146352 318792 146358 318844
rect 91738 314236 91744 314288
rect 91796 314276 91802 314288
rect 94590 314276 94596 314288
rect 91796 314248 94596 314276
rect 91796 314236 91802 314248
rect 94590 314236 94596 314248
rect 94648 314236 94654 314288
rect 82630 311856 82636 311908
rect 82688 311896 82694 311908
rect 579982 311896 579988 311908
rect 82688 311868 579988 311896
rect 82688 311856 82694 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 113082 305600 113088 305652
rect 113140 305640 113146 305652
rect 213178 305640 213184 305652
rect 113140 305612 213184 305640
rect 113140 305600 113146 305612
rect 213178 305600 213184 305612
rect 213236 305600 213242 305652
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 147674 305028 147680 305040
rect 3292 305000 147680 305028
rect 3292 304988 3298 305000
rect 147674 304988 147680 305000
rect 147732 304988 147738 305040
rect 79962 298120 79968 298172
rect 80020 298160 80026 298172
rect 580166 298160 580172 298172
rect 80020 298132 580172 298160
rect 80020 298120 80026 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 94590 295332 94596 295384
rect 94648 295372 94654 295384
rect 97258 295372 97264 295384
rect 94648 295344 97264 295372
rect 94648 295332 94654 295344
rect 97258 295332 97264 295344
rect 97316 295332 97322 295384
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 146386 292584 146392 292596
rect 3476 292556 146392 292584
rect 3476 292544 3482 292556
rect 146386 292544 146392 292556
rect 146444 292544 146450 292596
rect 97258 282888 97264 282940
rect 97316 282928 97322 282940
rect 97316 282900 98040 282928
rect 97316 282888 97322 282900
rect 98012 282860 98040 282900
rect 99466 282860 99472 282872
rect 98012 282832 99472 282860
rect 99466 282820 99472 282832
rect 99524 282820 99530 282872
rect 99466 278672 99472 278724
rect 99524 278712 99530 278724
rect 101490 278712 101496 278724
rect 99524 278684 101496 278712
rect 99524 278672 99530 278684
rect 101490 278672 101496 278684
rect 101548 278672 101554 278724
rect 101490 275204 101496 275256
rect 101548 275244 101554 275256
rect 102134 275244 102140 275256
rect 101548 275216 102140 275244
rect 101548 275204 101554 275216
rect 102134 275204 102140 275216
rect 102192 275204 102198 275256
rect 78582 271872 78588 271924
rect 78640 271912 78646 271924
rect 580166 271912 580172 271924
rect 78640 271884 580172 271912
rect 78640 271872 78646 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 102134 269084 102140 269136
rect 102192 269124 102198 269136
rect 104158 269124 104164 269136
rect 102192 269096 104164 269124
rect 102192 269084 102198 269096
rect 104158 269084 104164 269096
rect 104216 269084 104222 269136
rect 77202 266976 77208 267028
rect 77260 267016 77266 267028
rect 168466 267016 168472 267028
rect 77260 266988 168472 267016
rect 77260 266976 77266 266988
rect 168466 266976 168472 266988
rect 168524 266976 168530 267028
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 149054 266404 149060 266416
rect 3108 266376 149060 266404
rect 3108 266364 3114 266376
rect 149054 266364 149060 266376
rect 149112 266364 149118 266416
rect 106918 266296 106924 266348
rect 106976 266336 106982 266348
rect 195974 266336 195980 266348
rect 106976 266308 195980 266336
rect 106976 266296 106982 266308
rect 195974 266296 195980 266308
rect 196032 266296 196038 266348
rect 101950 266228 101956 266280
rect 102008 266268 102014 266280
rect 193214 266268 193220 266280
rect 102008 266240 193220 266268
rect 102008 266228 102014 266240
rect 193214 266228 193220 266240
rect 193272 266228 193278 266280
rect 107470 266160 107476 266212
rect 107528 266200 107534 266212
rect 202874 266200 202880 266212
rect 107528 266172 202880 266200
rect 107528 266160 107534 266172
rect 202874 266160 202880 266172
rect 202932 266160 202938 266212
rect 92290 266092 92296 266144
rect 92348 266132 92354 266144
rect 225874 266132 225880 266144
rect 92348 266104 225880 266132
rect 92348 266092 92354 266104
rect 225874 266092 225880 266104
rect 225932 266092 225938 266144
rect 86862 266024 86868 266076
rect 86920 266064 86926 266076
rect 225598 266064 225604 266076
rect 86920 266036 225604 266064
rect 86920 266024 86926 266036
rect 225598 266024 225604 266036
rect 225656 266024 225662 266076
rect 85390 265956 85396 266008
rect 85448 265996 85454 266008
rect 231118 265996 231124 266008
rect 85448 265968 231124 265996
rect 85448 265956 85454 265968
rect 231118 265956 231124 265968
rect 231176 265956 231182 266008
rect 88242 265888 88248 265940
rect 88300 265928 88306 265940
rect 175274 265928 175280 265940
rect 88300 265900 175280 265928
rect 88300 265888 88306 265900
rect 175274 265888 175280 265900
rect 175332 265888 175338 265940
rect 182082 265888 182088 265940
rect 182140 265928 182146 265940
rect 358906 265928 358912 265940
rect 182140 265900 358912 265928
rect 182140 265888 182146 265900
rect 358906 265888 358912 265900
rect 358964 265888 358970 265940
rect 53190 265820 53196 265872
rect 53248 265860 53254 265872
rect 259546 265860 259552 265872
rect 53248 265832 259552 265860
rect 53248 265820 53254 265832
rect 259546 265820 259552 265832
rect 259604 265820 259610 265872
rect 54294 265752 54300 265804
rect 54352 265792 54358 265804
rect 313274 265792 313280 265804
rect 54352 265764 313280 265792
rect 54352 265752 54358 265764
rect 313274 265752 313280 265764
rect 313332 265752 313338 265804
rect 54202 265684 54208 265736
rect 54260 265724 54266 265736
rect 317414 265724 317420 265736
rect 54260 265696 317420 265724
rect 54260 265684 54266 265696
rect 317414 265684 317420 265696
rect 317472 265684 317478 265736
rect 88242 265616 88248 265668
rect 88300 265656 88306 265668
rect 580258 265656 580264 265668
rect 88300 265628 580264 265656
rect 88300 265616 88306 265628
rect 580258 265616 580264 265628
rect 580316 265616 580322 265668
rect 115198 265548 115204 265600
rect 115256 265588 115262 265600
rect 200114 265588 200120 265600
rect 115256 265560 200120 265588
rect 115256 265548 115262 265560
rect 200114 265548 200120 265560
rect 200172 265548 200178 265600
rect 94498 265480 94504 265532
rect 94556 265520 94562 265532
rect 178034 265520 178040 265532
rect 94556 265492 178040 265520
rect 94556 265480 94562 265492
rect 178034 265480 178040 265492
rect 178092 265480 178098 265532
rect 187602 265480 187608 265532
rect 187660 265520 187666 265532
rect 251910 265520 251916 265532
rect 187660 265492 251916 265520
rect 187660 265480 187666 265492
rect 251910 265480 251916 265492
rect 251968 265480 251974 265532
rect 184750 264936 184756 264988
rect 184808 264976 184814 264988
rect 186958 264976 186964 264988
rect 184808 264948 186964 264976
rect 184808 264936 184814 264948
rect 186958 264936 186964 264948
rect 187016 264936 187022 264988
rect 36538 264868 36544 264920
rect 36596 264908 36602 264920
rect 131114 264908 131120 264920
rect 36596 264880 131120 264908
rect 36596 264868 36602 264880
rect 131114 264868 131120 264880
rect 131172 264868 131178 264920
rect 133782 264868 133788 264920
rect 133840 264908 133846 264920
rect 198090 264908 198096 264920
rect 133840 264880 198096 264908
rect 133840 264868 133846 264880
rect 198090 264868 198096 264880
rect 198148 264868 198154 264920
rect 209590 264868 209596 264920
rect 209648 264908 209654 264920
rect 268470 264908 268476 264920
rect 209648 264880 268476 264908
rect 209648 264868 209654 264880
rect 268470 264868 268476 264880
rect 268528 264868 268534 264920
rect 55858 264800 55864 264852
rect 55916 264840 55922 264852
rect 155954 264840 155960 264852
rect 55916 264812 155960 264840
rect 55916 264800 55922 264812
rect 155954 264800 155960 264812
rect 156012 264800 156018 264852
rect 173802 264800 173808 264852
rect 173860 264840 173866 264852
rect 252554 264840 252560 264852
rect 173860 264812 252560 264840
rect 173860 264800 173866 264812
rect 252554 264800 252560 264812
rect 252612 264800 252618 264852
rect 119982 264732 119988 264784
rect 120040 264772 120046 264784
rect 223666 264772 223672 264784
rect 120040 264744 223672 264772
rect 120040 264732 120046 264744
rect 223666 264732 223672 264744
rect 223724 264732 223730 264784
rect 8202 264664 8208 264716
rect 8260 264704 8266 264716
rect 124214 264704 124220 264716
rect 8260 264676 124220 264704
rect 8260 264664 8266 264676
rect 124214 264664 124220 264676
rect 124272 264664 124278 264716
rect 131022 264664 131028 264716
rect 131080 264704 131086 264716
rect 228542 264704 228548 264716
rect 131080 264676 228548 264704
rect 131080 264664 131086 264676
rect 228542 264664 228548 264676
rect 228600 264664 228606 264716
rect 111518 264596 111524 264648
rect 111576 264636 111582 264648
rect 229462 264636 229468 264648
rect 111576 264608 229468 264636
rect 111576 264596 111582 264608
rect 229462 264596 229468 264608
rect 229520 264596 229526 264648
rect 100662 264528 100668 264580
rect 100720 264568 100726 264580
rect 231302 264568 231308 264580
rect 100720 264540 231308 264568
rect 100720 264528 100726 264540
rect 231302 264528 231308 264540
rect 231360 264528 231366 264580
rect 90910 264460 90916 264512
rect 90968 264500 90974 264512
rect 227898 264500 227904 264512
rect 90968 264472 227904 264500
rect 90968 264460 90974 264472
rect 227898 264460 227904 264472
rect 227956 264460 227962 264512
rect 59538 264392 59544 264444
rect 59596 264432 59602 264444
rect 273346 264432 273352 264444
rect 59596 264404 273352 264432
rect 59596 264392 59602 264404
rect 273346 264392 273352 264404
rect 273404 264392 273410 264444
rect 54386 264324 54392 264376
rect 54444 264364 54450 264376
rect 276106 264364 276112 264376
rect 54444 264336 276112 264364
rect 54444 264324 54450 264336
rect 276106 264324 276112 264336
rect 276164 264324 276170 264376
rect 107562 264256 107568 264308
rect 107620 264296 107626 264308
rect 399478 264296 399484 264308
rect 107620 264268 399484 264296
rect 107620 264256 107626 264268
rect 399478 264256 399484 264268
rect 399536 264256 399542 264308
rect 104802 264188 104808 264240
rect 104860 264228 104866 264240
rect 542354 264228 542360 264240
rect 104860 264200 542360 264228
rect 104860 264188 104866 264200
rect 542354 264188 542360 264200
rect 542412 264188 542418 264240
rect 35158 264120 35164 264172
rect 35216 264160 35222 264172
rect 128354 264160 128360 264172
rect 35216 264132 128360 264160
rect 35216 264120 35222 264132
rect 128354 264120 128360 264132
rect 128412 264120 128418 264172
rect 139302 264120 139308 264172
rect 139360 264160 139366 264172
rect 201586 264160 201592 264172
rect 139360 264132 201592 264160
rect 139360 264120 139366 264132
rect 201586 264120 201592 264132
rect 201644 264120 201650 264172
rect 223482 264120 223488 264172
rect 223540 264160 223546 264172
rect 260098 264160 260104 264172
rect 223540 264132 260104 264160
rect 223540 264120 223546 264132
rect 260098 264120 260104 264132
rect 260156 264120 260162 264172
rect 33778 264052 33784 264104
rect 33836 264092 33842 264104
rect 125594 264092 125600 264104
rect 33836 264064 125600 264092
rect 33836 264052 33842 264064
rect 125594 264052 125600 264064
rect 125652 264052 125658 264104
rect 161382 264052 161388 264104
rect 161440 264092 161446 264104
rect 216398 264092 216404 264104
rect 161440 264064 216404 264092
rect 161440 264052 161446 264064
rect 216398 264052 216404 264064
rect 216456 264052 216462 264104
rect 47578 263984 47584 264036
rect 47636 264024 47642 264036
rect 139394 264024 139400 264036
rect 47636 263996 139400 264024
rect 47636 263984 47642 263996
rect 139394 263984 139400 263996
rect 139452 263984 139458 264036
rect 201402 263984 201408 264036
rect 201460 264024 201466 264036
rect 246298 264024 246304 264036
rect 201460 263996 246304 264024
rect 201460 263984 201466 263996
rect 246298 263984 246304 263996
rect 246356 263984 246362 264036
rect 119338 263916 119344 263968
rect 119396 263956 119402 263968
rect 205634 263956 205640 263968
rect 119396 263928 205640 263956
rect 119396 263916 119402 263928
rect 205634 263916 205640 263928
rect 205692 263916 205698 263968
rect 119982 263848 119988 263900
rect 120040 263888 120046 263900
rect 196526 263888 196532 263900
rect 120040 263860 196532 263888
rect 120040 263848 120046 263860
rect 196526 263848 196532 263860
rect 196584 263848 196590 263900
rect 89530 263780 89536 263832
rect 89588 263820 89594 263832
rect 165706 263820 165712 263832
rect 89588 263792 165712 263820
rect 89588 263780 89594 263792
rect 165706 263780 165712 263792
rect 165764 263780 165770 263832
rect 99282 263508 99288 263560
rect 99340 263548 99346 263560
rect 228358 263548 228364 263560
rect 99340 263520 228364 263548
rect 99340 263508 99346 263520
rect 228358 263508 228364 263520
rect 228416 263508 228422 263560
rect 231394 263508 231400 263560
rect 231452 263548 231458 263560
rect 310514 263548 310520 263560
rect 231452 263520 310520 263548
rect 231452 263508 231458 263520
rect 310514 263508 310520 263520
rect 310572 263508 310578 263560
rect 108942 263440 108948 263492
rect 109000 263480 109006 263492
rect 385678 263480 385684 263492
rect 109000 263452 385684 263480
rect 109000 263440 109006 263452
rect 385678 263440 385684 263452
rect 385736 263440 385742 263492
rect 106090 263372 106096 263424
rect 106148 263412 106154 263424
rect 382918 263412 382924 263424
rect 106148 263384 382924 263412
rect 106148 263372 106154 263384
rect 382918 263372 382924 263384
rect 382976 263372 382982 263424
rect 103422 263304 103428 263356
rect 103480 263344 103486 263356
rect 381538 263344 381544 263356
rect 103480 263316 381544 263344
rect 103480 263304 103486 263316
rect 381538 263304 381544 263316
rect 381596 263304 381602 263356
rect 97810 263236 97816 263288
rect 97868 263276 97874 263288
rect 377398 263276 377404 263288
rect 97868 263248 377404 263276
rect 97868 263236 97874 263248
rect 377398 263236 377404 263248
rect 377456 263236 377462 263288
rect 101950 263168 101956 263220
rect 102008 263208 102014 263220
rect 396718 263208 396724 263220
rect 102008 263180 396724 263208
rect 102008 263168 102014 263180
rect 396718 263168 396724 263180
rect 396776 263168 396782 263220
rect 99282 263100 99288 263152
rect 99340 263140 99346 263152
rect 395338 263140 395344 263152
rect 99340 263112 395344 263140
rect 99340 263100 99346 263112
rect 395338 263100 395344 263112
rect 395396 263100 395402 263152
rect 91002 263032 91008 263084
rect 91060 263072 91066 263084
rect 389818 263072 389824 263084
rect 91060 263044 389824 263072
rect 91060 263032 91066 263044
rect 389818 263032 389824 263044
rect 389876 263032 389882 263084
rect 93762 262964 93768 263016
rect 93820 263004 93826 263016
rect 392578 263004 392584 263016
rect 93820 262976 392584 263004
rect 93820 262964 93826 262976
rect 392578 262964 392584 262976
rect 392636 262964 392642 263016
rect 86862 262896 86868 262948
rect 86920 262936 86926 262948
rect 388438 262936 388444 262948
rect 86920 262908 388444 262936
rect 86920 262896 86926 262908
rect 388438 262896 388444 262908
rect 388496 262896 388502 262948
rect 110322 262828 110328 262880
rect 110380 262868 110386 262880
rect 412634 262868 412640 262880
rect 110380 262840 412640 262868
rect 110380 262828 110386 262840
rect 412634 262828 412640 262840
rect 412692 262828 412698 262880
rect 56042 262760 56048 262812
rect 56100 262800 56106 262812
rect 115934 262800 115940 262812
rect 56100 262772 115940 262800
rect 56100 262760 56106 262772
rect 115934 262760 115940 262772
rect 115992 262760 115998 262812
rect 117222 262760 117228 262812
rect 117280 262800 117286 262812
rect 225506 262800 225512 262812
rect 117280 262772 225512 262800
rect 117280 262760 117286 262772
rect 225506 262760 225512 262772
rect 225564 262760 225570 262812
rect 234246 262760 234252 262812
rect 234304 262800 234310 262812
rect 266446 262800 266452 262812
rect 234304 262772 266452 262800
rect 234304 262760 234310 262772
rect 266446 262760 266452 262772
rect 266504 262760 266510 262812
rect 22738 262692 22744 262744
rect 22796 262732 22802 262744
rect 129734 262732 129740 262744
rect 22796 262704 129740 262732
rect 22796 262692 22802 262704
rect 129734 262692 129740 262704
rect 129792 262692 129798 262744
rect 162118 262692 162124 262744
rect 162176 262732 162182 262744
rect 173894 262732 173900 262744
rect 162176 262704 173900 262732
rect 162176 262692 162182 262704
rect 173894 262692 173900 262704
rect 173952 262692 173958 262744
rect 181990 262692 181996 262744
rect 182048 262732 182054 262744
rect 188338 262732 188344 262744
rect 182048 262704 188344 262732
rect 182048 262692 182054 262704
rect 188338 262692 188344 262704
rect 188396 262692 188402 262744
rect 198550 262692 198556 262744
rect 198608 262732 198614 262744
rect 291838 262732 291844 262744
rect 198608 262704 291844 262732
rect 198608 262692 198614 262704
rect 291838 262692 291844 262704
rect 291896 262692 291902 262744
rect 25498 262624 25504 262676
rect 25556 262664 25562 262676
rect 132494 262664 132500 262676
rect 25556 262636 132500 262664
rect 25556 262624 25562 262636
rect 132494 262624 132500 262636
rect 132552 262624 132558 262676
rect 151722 262624 151728 262676
rect 151780 262664 151786 262676
rect 212534 262664 212540 262676
rect 151780 262636 212540 262664
rect 151780 262624 151786 262636
rect 212534 262624 212540 262636
rect 212592 262624 212598 262676
rect 21358 262556 21364 262608
rect 21416 262596 21422 262608
rect 126974 262596 126980 262608
rect 21416 262568 126980 262596
rect 21416 262556 21422 262568
rect 126974 262556 126980 262568
rect 127032 262556 127038 262608
rect 32398 262488 32404 262540
rect 32456 262528 32462 262540
rect 138014 262528 138020 262540
rect 32456 262500 138020 262528
rect 32456 262488 32462 262500
rect 138014 262488 138020 262500
rect 138072 262488 138078 262540
rect 117222 262420 117228 262472
rect 117280 262460 117286 262472
rect 201494 262460 201500 262472
rect 117280 262432 201500 262460
rect 117280 262420 117286 262432
rect 201494 262420 201500 262432
rect 201552 262420 201558 262472
rect 4798 262148 4804 262200
rect 4856 262188 4862 262200
rect 127066 262188 127072 262200
rect 4856 262160 127072 262188
rect 4856 262148 4862 262160
rect 127066 262148 127072 262160
rect 127124 262148 127130 262200
rect 144822 262148 144828 262200
rect 144880 262188 144886 262200
rect 202966 262188 202972 262200
rect 144880 262160 202972 262188
rect 144880 262148 144886 262160
rect 202966 262148 202972 262160
rect 203024 262148 203030 262200
rect 211062 262148 211068 262200
rect 211120 262188 211126 262200
rect 304258 262188 304264 262200
rect 211120 262160 304264 262188
rect 211120 262148 211126 262160
rect 304258 262148 304264 262160
rect 304316 262148 304322 262200
rect 97902 262080 97908 262132
rect 97960 262120 97966 262132
rect 229646 262120 229652 262132
rect 97960 262092 229652 262120
rect 97960 262080 97966 262092
rect 229646 262080 229652 262092
rect 229704 262080 229710 262132
rect 235442 262080 235448 262132
rect 235500 262120 235506 262132
rect 280154 262120 280160 262132
rect 235500 262092 280160 262120
rect 235500 262080 235506 262092
rect 280154 262080 280160 262092
rect 280212 262080 280218 262132
rect 59446 262012 59452 262064
rect 59504 262052 59510 262064
rect 265066 262052 265072 262064
rect 59504 262024 265072 262052
rect 59504 262012 59510 262024
rect 265066 262012 265072 262024
rect 265124 262012 265130 262064
rect 101858 261944 101864 261996
rect 101916 261984 101922 261996
rect 367738 261984 367744 261996
rect 101916 261956 367744 261984
rect 101916 261944 101922 261956
rect 367738 261944 367744 261956
rect 367796 261944 367802 261996
rect 104710 261876 104716 261928
rect 104768 261916 104774 261928
rect 370498 261916 370504 261928
rect 104768 261888 370504 261916
rect 104768 261876 104774 261888
rect 370498 261876 370504 261888
rect 370556 261876 370562 261928
rect 100662 261808 100668 261860
rect 100720 261848 100726 261860
rect 378778 261848 378784 261860
rect 100720 261820 378784 261848
rect 100720 261808 100726 261820
rect 378778 261808 378784 261820
rect 378836 261808 378842 261860
rect 92382 261740 92388 261792
rect 92440 261780 92446 261792
rect 376018 261780 376024 261792
rect 92440 261752 376024 261780
rect 92440 261740 92446 261752
rect 376018 261740 376024 261752
rect 376076 261740 376082 261792
rect 89622 261672 89628 261724
rect 89680 261712 89686 261724
rect 374638 261712 374644 261724
rect 89680 261684 374644 261712
rect 89680 261672 89686 261684
rect 374638 261672 374644 261684
rect 374696 261672 374702 261724
rect 96430 261604 96436 261656
rect 96488 261644 96494 261656
rect 393958 261644 393964 261656
rect 96488 261616 393964 261644
rect 96488 261604 96494 261616
rect 393958 261604 393964 261616
rect 394016 261604 394022 261656
rect 108850 261536 108856 261588
rect 108908 261576 108914 261588
rect 429194 261576 429200 261588
rect 108908 261548 429200 261576
rect 108908 261536 108914 261548
rect 429194 261536 429200 261548
rect 429252 261536 429258 261588
rect 95142 261468 95148 261520
rect 95200 261508 95206 261520
rect 558178 261508 558184 261520
rect 95200 261480 558184 261508
rect 95200 261468 95206 261480
rect 558178 261468 558184 261480
rect 558236 261468 558242 261520
rect 18598 261400 18604 261452
rect 18656 261440 18662 261452
rect 140866 261440 140872 261452
rect 18656 261412 140872 261440
rect 18656 261400 18662 261412
rect 140866 261400 140872 261412
rect 140924 261400 140930 261452
rect 193030 261400 193036 261452
rect 193088 261440 193094 261452
rect 284938 261440 284944 261452
rect 193088 261412 284944 261440
rect 193088 261400 193094 261412
rect 284938 261400 284944 261412
rect 284996 261400 285002 261452
rect 17218 261332 17224 261384
rect 17276 261372 17282 261384
rect 138106 261372 138112 261384
rect 17276 261344 138112 261372
rect 17276 261332 17282 261344
rect 138106 261332 138112 261344
rect 138164 261332 138170 261384
rect 190362 261332 190368 261384
rect 190420 261372 190426 261384
rect 282178 261372 282184 261384
rect 190420 261344 282184 261372
rect 190420 261332 190426 261344
rect 282178 261332 282184 261344
rect 282236 261332 282242 261384
rect 14458 261264 14464 261316
rect 14516 261304 14522 261316
rect 132586 261304 132592 261316
rect 14516 261276 132592 261304
rect 14516 261264 14522 261276
rect 132586 261264 132592 261276
rect 132644 261264 132650 261316
rect 142062 261264 142068 261316
rect 142120 261304 142126 261316
rect 228634 261304 228640 261316
rect 142120 261276 228640 261304
rect 142120 261264 142126 261276
rect 228634 261264 228640 261276
rect 228692 261264 228698 261316
rect 232498 261264 232504 261316
rect 232556 261304 232562 261316
rect 273438 261304 273444 261316
rect 232556 261276 273444 261304
rect 232556 261264 232562 261276
rect 273438 261264 273444 261276
rect 273496 261264 273502 261316
rect 11698 261196 11704 261248
rect 11756 261236 11762 261248
rect 129826 261236 129832 261248
rect 11756 261208 129832 261236
rect 11756 261196 11762 261208
rect 129826 261196 129832 261208
rect 129884 261196 129890 261248
rect 148962 261196 148968 261248
rect 149020 261236 149026 261248
rect 211246 261236 211252 261248
rect 149020 261208 211252 261236
rect 149020 261196 149026 261208
rect 211246 261196 211252 261208
rect 211304 261196 211310 261248
rect 238202 261196 238208 261248
rect 238260 261236 238266 261248
rect 258074 261236 258080 261248
rect 238260 261208 258080 261236
rect 238260 261196 238266 261208
rect 258074 261196 258080 261208
rect 258132 261196 258138 261248
rect 29638 261128 29644 261180
rect 29696 261168 29702 261180
rect 135254 261168 135260 261180
rect 29696 261140 135260 261168
rect 29696 261128 29702 261140
rect 135254 261128 135260 261140
rect 135312 261128 135318 261180
rect 200850 261128 200856 261180
rect 200908 261168 200914 261180
rect 224770 261168 224776 261180
rect 200908 261140 224776 261168
rect 200908 261128 200914 261140
rect 224770 261128 224776 261140
rect 224828 261128 224834 261180
rect 117130 261060 117136 261112
rect 117188 261100 117194 261112
rect 215938 261100 215944 261112
rect 117188 261072 215944 261100
rect 117188 261060 117194 261072
rect 215938 261060 215944 261072
rect 215996 261060 216002 261112
rect 118602 260992 118608 261044
rect 118660 261032 118666 261044
rect 210418 261032 210424 261044
rect 118660 261004 210424 261032
rect 118660 260992 118666 261004
rect 210418 260992 210424 261004
rect 210476 260992 210482 261044
rect 111518 260924 111524 260976
rect 111576 260964 111582 260976
rect 197998 260964 198004 260976
rect 111576 260936 198004 260964
rect 111576 260924 111582 260936
rect 197998 260924 198004 260936
rect 198056 260924 198062 260976
rect 41322 260856 41328 260908
rect 41380 260896 41386 260908
rect 124306 260896 124312 260908
rect 41380 260868 124312 260896
rect 41380 260856 41386 260868
rect 124306 260856 124312 260868
rect 124364 260856 124370 260908
rect 104158 260788 104164 260840
rect 104216 260828 104222 260840
rect 106642 260828 106648 260840
rect 104216 260800 106648 260828
rect 104216 260788 104222 260800
rect 106642 260788 106648 260800
rect 106700 260788 106706 260840
rect 172422 260788 172428 260840
rect 172480 260828 172486 260840
rect 173158 260828 173164 260840
rect 172480 260800 173164 260828
rect 172480 260788 172486 260800
rect 173158 260788 173164 260800
rect 173216 260788 173222 260840
rect 199654 260788 199660 260840
rect 199712 260828 199718 260840
rect 229554 260828 229560 260840
rect 199712 260800 229560 260828
rect 199712 260788 199718 260800
rect 229554 260788 229560 260800
rect 229612 260788 229618 260840
rect 114462 260720 114468 260772
rect 114520 260760 114526 260772
rect 206278 260760 206284 260772
rect 114520 260732 206284 260760
rect 114520 260720 114526 260732
rect 206278 260720 206284 260732
rect 206336 260720 206342 260772
rect 56134 260652 56140 260704
rect 56192 260692 56198 260704
rect 103514 260692 103520 260704
rect 56192 260664 103520 260692
rect 56192 260652 56198 260664
rect 103514 260652 103520 260664
rect 103572 260652 103578 260704
rect 114370 260652 114376 260704
rect 114428 260692 114434 260704
rect 209038 260692 209044 260704
rect 114428 260664 209044 260692
rect 114428 260652 114434 260664
rect 209038 260652 209044 260664
rect 209096 260652 209102 260704
rect 15838 260584 15844 260636
rect 15896 260624 15902 260636
rect 135346 260624 135352 260636
rect 15896 260596 135352 260624
rect 15896 260584 15902 260596
rect 135346 260584 135352 260596
rect 135404 260584 135410 260636
rect 208302 260584 208308 260636
rect 208360 260624 208366 260636
rect 304994 260624 305000 260636
rect 208360 260596 305000 260624
rect 208360 260584 208366 260596
rect 304994 260584 305000 260596
rect 305052 260584 305058 260636
rect 90910 260516 90916 260568
rect 90968 260556 90974 260568
rect 213362 260556 213368 260568
rect 90968 260528 213368 260556
rect 90968 260516 90974 260528
rect 213362 260516 213368 260528
rect 213420 260516 213426 260568
rect 213638 260516 213644 260568
rect 213696 260556 213702 260568
rect 226886 260556 226892 260568
rect 213696 260528 226892 260556
rect 213696 260516 213702 260528
rect 226886 260516 226892 260528
rect 226944 260516 226950 260568
rect 238294 260516 238300 260568
rect 238352 260556 238358 260568
rect 270586 260556 270592 260568
rect 238352 260528 270592 260556
rect 238352 260516 238358 260528
rect 270586 260516 270592 260528
rect 270644 260516 270650 260568
rect 102042 260448 102048 260500
rect 102100 260488 102106 260500
rect 228450 260488 228456 260500
rect 102100 260460 228456 260488
rect 102100 260448 102106 260460
rect 228450 260448 228456 260460
rect 228508 260448 228514 260500
rect 234154 260448 234160 260500
rect 234212 260488 234218 260500
rect 295334 260488 295340 260500
rect 234212 260460 295340 260488
rect 234212 260448 234218 260460
rect 295334 260448 295340 260460
rect 295392 260448 295398 260500
rect 99190 260380 99196 260432
rect 99248 260420 99254 260432
rect 363598 260420 363604 260432
rect 99248 260392 363604 260420
rect 99248 260380 99254 260392
rect 363598 260380 363604 260392
rect 363656 260380 363662 260432
rect 93670 260312 93676 260364
rect 93728 260352 93734 260364
rect 358078 260352 358084 260364
rect 93728 260324 358084 260352
rect 93728 260312 93734 260324
rect 358078 260312 358084 260324
rect 358136 260312 358142 260364
rect 96338 260244 96344 260296
rect 96396 260284 96402 260296
rect 360838 260284 360844 260296
rect 96396 260256 360844 260284
rect 96396 260244 96402 260256
rect 360838 260244 360844 260256
rect 360896 260244 360902 260296
rect 85390 260176 85396 260228
rect 85448 260216 85454 260228
rect 371878 260216 371884 260228
rect 85448 260188 371884 260216
rect 85448 260176 85454 260188
rect 371878 260176 371884 260188
rect 371936 260176 371942 260228
rect 88150 260108 88156 260160
rect 88208 260148 88214 260160
rect 425698 260148 425704 260160
rect 88208 260120 425704 260148
rect 88208 260108 88214 260120
rect 425698 260108 425704 260120
rect 425756 260108 425762 260160
rect 260742 245556 260748 245608
rect 260800 245596 260806 245608
rect 580166 245596 580172 245608
rect 260800 245568 580172 245596
rect 260800 245556 260806 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 55766 229100 55772 229152
rect 55824 229140 55830 229152
rect 59814 229140 59820 229152
rect 55824 229112 59820 229140
rect 55824 229100 55830 229112
rect 59814 229100 59820 229112
rect 59872 229100 59878 229152
rect 57422 218016 57428 218068
rect 57480 218056 57486 218068
rect 58526 218056 58532 218068
rect 57480 218028 58532 218056
rect 57480 218016 57486 218028
rect 58526 218016 58532 218028
rect 58584 218016 58590 218068
rect 3050 215228 3056 215280
rect 3108 215268 3114 215280
rect 11698 215268 11704 215280
rect 3108 215240 11704 215268
rect 3108 215228 3114 215240
rect 11698 215228 11704 215240
rect 11756 215228 11762 215280
rect 54202 213868 54208 213920
rect 54260 213908 54266 213920
rect 57514 213908 57520 213920
rect 54260 213880 57520 213908
rect 54260 213868 54266 213880
rect 57514 213868 57520 213880
rect 57572 213868 57578 213920
rect 54294 197276 54300 197328
rect 54352 197316 54358 197328
rect 57514 197316 57520 197328
rect 54352 197288 57520 197316
rect 54352 197276 54358 197288
rect 57514 197276 57520 197288
rect 57572 197276 57578 197328
rect 54662 194488 54668 194540
rect 54720 194528 54726 194540
rect 57514 194528 57520 194540
rect 54720 194500 57520 194528
rect 54720 194488 54726 194500
rect 57514 194488 57520 194500
rect 57572 194488 57578 194540
rect 271138 193128 271144 193180
rect 271196 193168 271202 193180
rect 580166 193168 580172 193180
rect 271196 193140 580172 193168
rect 271196 193128 271202 193140
rect 580166 193128 580172 193140
rect 580224 193128 580230 193180
rect 53282 191768 53288 191820
rect 53340 191808 53346 191820
rect 57514 191808 57520 191820
rect 53340 191780 57520 191808
rect 53340 191768 53346 191780
rect 57514 191768 57520 191780
rect 57572 191768 57578 191820
rect 3326 188844 3332 188896
rect 3384 188884 3390 188896
rect 7558 188884 7564 188896
rect 3384 188856 7564 188884
rect 3384 188844 3390 188856
rect 7558 188844 7564 188856
rect 7616 188844 7622 188896
rect 54754 182112 54760 182164
rect 54812 182152 54818 182164
rect 57514 182152 57520 182164
rect 54812 182124 57520 182152
rect 54812 182112 54818 182124
rect 57514 182112 57520 182124
rect 57572 182112 57578 182164
rect 53374 177964 53380 178016
rect 53432 178004 53438 178016
rect 57514 178004 57520 178016
rect 53432 177976 57520 178004
rect 53432 177964 53438 177976
rect 57514 177964 57520 177976
rect 57572 177964 57578 178016
rect 54570 175176 54576 175228
rect 54628 175216 54634 175228
rect 57514 175216 57520 175228
rect 54628 175188 57520 175216
rect 54628 175176 54634 175188
rect 57514 175176 57520 175188
rect 57572 175176 57578 175228
rect 3050 164160 3056 164212
rect 3108 164200 3114 164212
rect 14458 164200 14464 164212
rect 3108 164172 14464 164200
rect 3108 164160 3114 164172
rect 14458 164160 14464 164172
rect 14516 164160 14522 164212
rect 53466 160012 53472 160064
rect 53524 160052 53530 160064
rect 57422 160052 57428 160064
rect 53524 160024 57428 160052
rect 53524 160012 53530 160024
rect 57422 160012 57428 160024
rect 57480 160012 57486 160064
rect 53190 155864 53196 155916
rect 53248 155904 53254 155916
rect 57514 155904 57520 155916
rect 53248 155876 57520 155904
rect 53248 155864 53254 155876
rect 57514 155864 57520 155876
rect 57572 155864 57578 155916
rect 54846 153144 54852 153196
rect 54904 153184 54910 153196
rect 57514 153184 57520 153196
rect 54904 153156 57520 153184
rect 54904 153144 54910 153156
rect 57514 153144 57520 153156
rect 57572 153144 57578 153196
rect 53558 147568 53564 147620
rect 53616 147608 53622 147620
rect 57422 147608 57428 147620
rect 53616 147580 57428 147608
rect 53616 147568 53622 147580
rect 57422 147568 57428 147580
rect 57480 147568 57486 147620
rect 53650 143488 53656 143540
rect 53708 143528 53714 143540
rect 57514 143528 57520 143540
rect 53708 143500 57520 143528
rect 53708 143488 53714 143500
rect 57514 143488 57520 143500
rect 57572 143488 57578 143540
rect 3050 137912 3056 137964
rect 3108 137952 3114 137964
rect 17218 137952 17224 137964
rect 3108 137924 17224 137952
rect 3108 137912 3114 137924
rect 17218 137912 17224 137924
rect 17276 137912 17282 137964
rect 57514 136552 57520 136604
rect 57572 136592 57578 136604
rect 59814 136592 59820 136604
rect 57572 136564 59820 136592
rect 57572 136552 57578 136564
rect 59814 136552 59820 136564
rect 59872 136552 59878 136604
rect 54386 134716 54392 134768
rect 54444 134756 54450 134768
rect 57422 134756 57428 134768
rect 54444 134728 57428 134756
rect 54444 134716 54450 134728
rect 57422 134716 57428 134728
rect 57480 134716 57486 134768
rect 53742 131044 53748 131096
rect 53800 131084 53806 131096
rect 57606 131084 57612 131096
rect 53800 131056 57612 131084
rect 53800 131044 53806 131056
rect 57606 131044 57612 131056
rect 57664 131044 57670 131096
rect 57698 127916 57704 127968
rect 57756 127956 57762 127968
rect 58710 127956 58716 127968
rect 57756 127928 58716 127956
rect 57756 127916 57762 127928
rect 58710 127916 58716 127928
rect 58768 127916 58774 127968
rect 54938 118600 54944 118652
rect 54996 118640 55002 118652
rect 57606 118640 57612 118652
rect 54996 118612 57612 118640
rect 54996 118600 55002 118612
rect 57606 118600 57612 118612
rect 57664 118600 57670 118652
rect 55030 113092 55036 113144
rect 55088 113132 55094 113144
rect 57606 113132 57612 113144
rect 55088 113104 57612 113132
rect 55088 113092 55094 113104
rect 57606 113092 57612 113104
rect 57664 113092 57670 113144
rect 3326 111732 3332 111784
rect 3384 111772 3390 111784
rect 15838 111772 15844 111784
rect 3384 111744 15844 111772
rect 3384 111732 3390 111744
rect 15838 111732 15844 111744
rect 15896 111732 15902 111784
rect 57698 106224 57704 106276
rect 57756 106264 57762 106276
rect 59814 106264 59820 106276
rect 57756 106236 59820 106264
rect 57756 106224 57762 106236
rect 59814 106224 59820 106236
rect 59872 106224 59878 106276
rect 410518 100648 410524 100700
rect 410576 100688 410582 100700
rect 580166 100688 580172 100700
rect 410576 100660 580172 100688
rect 410576 100648 410582 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 3234 97928 3240 97980
rect 3292 97968 3298 97980
rect 18598 97968 18604 97980
rect 3292 97940 18604 97968
rect 3292 97928 3298 97940
rect 18598 97928 18604 97940
rect 18656 97928 18662 97980
rect 2958 85484 2964 85536
rect 3016 85524 3022 85536
rect 32398 85524 32404 85536
rect 3016 85496 32404 85524
rect 3016 85484 3022 85496
rect 32398 85484 32404 85496
rect 32456 85484 32462 85536
rect 3326 71680 3332 71732
rect 3384 71720 3390 71732
rect 29638 71720 29644 71732
rect 3384 71692 29644 71720
rect 3384 71680 3390 71692
rect 29638 71680 29644 71692
rect 29696 71680 29702 71732
rect 54478 71680 54484 71732
rect 54536 71720 54542 71732
rect 57606 71720 57612 71732
rect 54536 71692 57612 71720
rect 54536 71680 54542 71692
rect 57606 71680 57612 71692
rect 57664 71680 57670 71732
rect 55122 62024 55128 62076
rect 55180 62064 55186 62076
rect 57054 62064 57060 62076
rect 55180 62036 57060 62064
rect 55180 62024 55186 62036
rect 57054 62024 57060 62036
rect 57112 62024 57118 62076
rect 580166 59956 580172 59968
rect 240888 59928 580172 59956
rect 240888 59900 240916 59928
rect 580166 59916 580172 59928
rect 580224 59916 580230 59968
rect 222102 59848 222108 59900
rect 222160 59888 222166 59900
rect 222160 59860 240824 59888
rect 222160 59848 222166 59860
rect 222562 59780 222568 59832
rect 222620 59820 222626 59832
rect 224126 59820 224132 59832
rect 222620 59792 224132 59820
rect 222620 59780 222626 59792
rect 224126 59780 224132 59792
rect 224184 59780 224190 59832
rect 224310 59780 224316 59832
rect 224368 59820 224374 59832
rect 224368 59792 238754 59820
rect 224368 59780 224374 59792
rect 224218 59712 224224 59764
rect 224276 59752 224282 59764
rect 224770 59752 224776 59764
rect 224276 59724 224776 59752
rect 224276 59712 224282 59724
rect 224770 59712 224776 59724
rect 224828 59712 224834 59764
rect 238726 59684 238754 59792
rect 240796 59752 240824 59860
rect 240870 59848 240876 59900
rect 240928 59848 240934 59900
rect 302234 59888 302240 59900
rect 241072 59860 302240 59888
rect 241072 59752 241100 59860
rect 302234 59848 302240 59860
rect 302292 59848 302298 59900
rect 263686 59820 263692 59832
rect 240796 59724 241100 59752
rect 248386 59792 263692 59820
rect 248386 59684 248414 59792
rect 263686 59780 263692 59792
rect 263744 59780 263750 59832
rect 238726 59656 248414 59684
rect 223574 59440 223580 59492
rect 223632 59480 223638 59492
rect 268378 59480 268384 59492
rect 223632 59452 268384 59480
rect 223632 59440 223638 59452
rect 268378 59440 268384 59452
rect 268436 59440 268442 59492
rect 224494 59372 224500 59424
rect 224552 59412 224558 59424
rect 276014 59412 276020 59424
rect 224552 59384 276020 59412
rect 224552 59372 224558 59384
rect 276014 59372 276020 59384
rect 276072 59372 276078 59424
rect 57790 59304 57796 59356
rect 57848 59344 57854 59356
rect 217042 59344 217048 59356
rect 57848 59316 217048 59344
rect 57848 59304 57854 59316
rect 217042 59304 217048 59316
rect 217100 59304 217106 59356
rect 217962 59304 217968 59356
rect 218020 59344 218026 59356
rect 229094 59344 229100 59356
rect 218020 59316 229100 59344
rect 218020 59304 218026 59316
rect 229094 59304 229100 59316
rect 229152 59304 229158 59356
rect 220906 59236 220912 59288
rect 220964 59276 220970 59288
rect 229370 59276 229376 59288
rect 220964 59248 229376 59276
rect 220964 59236 220970 59248
rect 229370 59236 229376 59248
rect 229428 59236 229434 59288
rect 221550 59168 221556 59220
rect 221608 59208 221614 59220
rect 230474 59208 230480 59220
rect 221608 59180 230480 59208
rect 221608 59168 221614 59180
rect 230474 59168 230480 59180
rect 230532 59168 230538 59220
rect 209866 59100 209872 59152
rect 209924 59140 209930 59152
rect 230658 59140 230664 59152
rect 209924 59112 230664 59140
rect 209924 59100 209930 59112
rect 230658 59100 230664 59112
rect 230716 59100 230722 59152
rect 150618 59032 150624 59084
rect 150676 59072 150682 59084
rect 151446 59072 151452 59084
rect 150676 59044 151452 59072
rect 150676 59032 150682 59044
rect 151446 59032 151452 59044
rect 151504 59032 151510 59084
rect 216766 59032 216772 59084
rect 216824 59072 216830 59084
rect 229278 59072 229284 59084
rect 216824 59044 229284 59072
rect 216824 59032 216830 59044
rect 229278 59032 229284 59044
rect 229336 59032 229342 59084
rect 149422 58964 149428 59016
rect 149480 59004 149486 59016
rect 150250 59004 150256 59016
rect 149480 58976 150256 59004
rect 149480 58964 149486 58976
rect 150250 58964 150256 58976
rect 150308 58964 150314 59016
rect 150710 58964 150716 59016
rect 150768 59004 150774 59016
rect 151722 59004 151728 59016
rect 150768 58976 151728 59004
rect 150768 58964 150774 58976
rect 151722 58964 151728 58976
rect 151780 58964 151786 59016
rect 215846 58964 215852 59016
rect 215904 59004 215910 59016
rect 229186 59004 229192 59016
rect 215904 58976 229192 59004
rect 215904 58964 215910 58976
rect 229186 58964 229192 58976
rect 229244 58964 229250 59016
rect 219158 58896 219164 58948
rect 219216 58936 219222 58948
rect 250438 58936 250444 58948
rect 219216 58908 250444 58936
rect 219216 58896 219222 58908
rect 250438 58896 250444 58908
rect 250496 58896 250502 58948
rect 211338 58828 211344 58880
rect 211396 58868 211402 58880
rect 240134 58868 240140 58880
rect 211396 58840 240140 58868
rect 211396 58828 211402 58840
rect 240134 58828 240140 58840
rect 240192 58828 240198 58880
rect 209222 58760 209228 58812
rect 209280 58800 209286 58812
rect 237374 58800 237380 58812
rect 209280 58772 237380 58800
rect 209280 58760 209286 58772
rect 237374 58760 237380 58772
rect 237432 58760 237438 58812
rect 214374 58692 214380 58744
rect 214432 58732 214438 58744
rect 227714 58732 227720 58744
rect 214432 58704 227720 58732
rect 214432 58692 214438 58704
rect 227714 58692 227720 58704
rect 227772 58692 227778 58744
rect 212258 58624 212264 58676
rect 212316 58664 212322 58676
rect 245654 58664 245660 58676
rect 212316 58636 245660 58664
rect 212316 58624 212322 58636
rect 245654 58624 245660 58636
rect 245712 58624 245718 58676
rect 210694 58556 210700 58608
rect 210752 58596 210758 58608
rect 230566 58596 230572 58608
rect 210752 58568 230572 58596
rect 210752 58556 210758 58568
rect 230566 58556 230572 58568
rect 230624 58556 230630 58608
rect 208946 58488 208952 58540
rect 209004 58528 209010 58540
rect 235994 58528 236000 58540
rect 209004 58500 236000 58528
rect 209004 58488 209010 58500
rect 235994 58488 236000 58500
rect 236052 58488 236058 58540
rect 214926 58420 214932 58472
rect 214984 58460 214990 58472
rect 262858 58460 262864 58472
rect 214984 58432 262864 58460
rect 214984 58420 214990 58432
rect 262858 58420 262864 58432
rect 262916 58420 262922 58472
rect 209498 58352 209504 58404
rect 209556 58392 209562 58404
rect 244366 58392 244372 58404
rect 209556 58364 244372 58392
rect 209556 58352 209562 58364
rect 244366 58352 244372 58364
rect 244424 58352 244430 58404
rect 216398 58284 216404 58336
rect 216456 58324 216462 58336
rect 342346 58324 342352 58336
rect 216456 58296 342352 58324
rect 216456 58284 216462 58296
rect 342346 58284 342352 58296
rect 342404 58284 342410 58336
rect 218514 58216 218520 58268
rect 218572 58256 218578 58268
rect 255406 58256 255412 58268
rect 218572 58228 255412 58256
rect 218572 58216 218578 58228
rect 255406 58216 255412 58228
rect 255464 58216 255470 58268
rect 220630 58148 220636 58200
rect 220688 58188 220694 58200
rect 253198 58188 253204 58200
rect 220688 58160 253204 58188
rect 220688 58148 220694 58160
rect 253198 58148 253204 58160
rect 253256 58148 253262 58200
rect 215570 58080 215576 58132
rect 215628 58120 215634 58132
rect 316678 58120 316684 58132
rect 215628 58092 316684 58120
rect 215628 58080 215634 58092
rect 316678 58080 316684 58092
rect 316736 58080 316742 58132
rect 180794 58012 180800 58064
rect 180852 58052 180858 58064
rect 181162 58052 181168 58064
rect 180852 58024 181168 58052
rect 180852 58012 180858 58024
rect 181162 58012 181168 58024
rect 181220 58012 181226 58064
rect 208670 58012 208676 58064
rect 208728 58052 208734 58064
rect 224954 58052 224960 58064
rect 208728 58024 224960 58052
rect 208728 58012 208734 58024
rect 224954 58012 224960 58024
rect 225012 58012 225018 58064
rect 180702 57944 180708 57996
rect 180760 57984 180766 57996
rect 181714 57984 181720 57996
rect 180760 57956 181720 57984
rect 180760 57944 180766 57956
rect 181714 57944 181720 57956
rect 181772 57944 181778 57996
rect 207750 57944 207756 57996
rect 207808 57984 207814 57996
rect 208302 57984 208308 57996
rect 207808 57956 208308 57984
rect 207808 57944 207814 57956
rect 208302 57944 208308 57956
rect 208360 57944 208366 57996
rect 216582 57944 216588 57996
rect 216640 57984 216646 57996
rect 216640 57956 219020 57984
rect 216640 57944 216646 57956
rect 218992 57928 219020 57956
rect 39942 57876 39948 57928
rect 40000 57916 40006 57928
rect 69934 57916 69940 57928
rect 40000 57888 69940 57916
rect 40000 57876 40006 57888
rect 69934 57876 69940 57888
rect 69992 57876 69998 57928
rect 76834 57916 76840 57928
rect 74506 57888 76840 57916
rect 34422 57808 34428 57860
rect 34480 57848 34486 57860
rect 68462 57848 68468 57860
rect 34480 57820 68468 57848
rect 34480 57808 34486 57820
rect 68462 57808 68468 57820
rect 68520 57808 68526 57860
rect 30282 57740 30288 57792
rect 30340 57780 30346 57792
rect 67542 57780 67548 57792
rect 30340 57752 67548 57780
rect 30340 57740 30346 57752
rect 67542 57740 67548 57752
rect 67600 57740 67606 57792
rect 74506 57780 74534 57888
rect 76834 57876 76840 57888
rect 76892 57876 76898 57928
rect 87874 57876 87880 57928
rect 87932 57916 87938 57928
rect 95326 57916 95332 57928
rect 87932 57888 95332 57916
rect 87932 57876 87938 57888
rect 95326 57876 95332 57888
rect 95384 57876 95390 57928
rect 95418 57876 95424 57928
rect 95476 57916 95482 57928
rect 103974 57916 103980 57928
rect 95476 57888 103980 57916
rect 95476 57876 95482 57888
rect 103974 57876 103980 57888
rect 104032 57876 104038 57928
rect 107102 57876 107108 57928
rect 107160 57916 107166 57928
rect 107160 57888 133184 57916
rect 107160 57876 107166 57888
rect 75086 57808 75092 57860
rect 75144 57848 75150 57860
rect 77386 57848 77392 57860
rect 75144 57820 77392 57848
rect 75144 57808 75150 57820
rect 77386 57808 77392 57820
rect 77444 57808 77450 57860
rect 91830 57808 91836 57860
rect 91888 57848 91894 57860
rect 113726 57848 113732 57860
rect 91888 57820 113732 57848
rect 91888 57808 91894 57820
rect 113726 57808 113732 57820
rect 113784 57808 113790 57860
rect 118142 57808 118148 57860
rect 118200 57848 118206 57860
rect 118602 57848 118608 57860
rect 118200 57820 118608 57848
rect 118200 57808 118206 57820
rect 118602 57808 118608 57820
rect 118660 57808 118666 57860
rect 120902 57808 120908 57860
rect 120960 57848 120966 57860
rect 120960 57820 126376 57848
rect 120960 57808 120966 57820
rect 78306 57780 78312 57792
rect 68296 57752 74534 57780
rect 75104 57752 78312 57780
rect 33042 57672 33048 57724
rect 33100 57712 33106 57724
rect 68094 57712 68100 57724
rect 33100 57684 68100 57712
rect 33100 57672 33106 57684
rect 68094 57672 68100 57684
rect 68152 57672 68158 57724
rect 28902 57604 28908 57656
rect 28960 57644 28966 57656
rect 66898 57644 66904 57656
rect 28960 57616 66904 57644
rect 28960 57604 28966 57616
rect 66898 57604 66904 57616
rect 66956 57604 66962 57656
rect 67542 57604 67548 57656
rect 67600 57644 67606 57656
rect 68296 57644 68324 57752
rect 73062 57672 73068 57724
rect 73120 57712 73126 57724
rect 73120 57684 74948 57712
rect 73120 57672 73126 57684
rect 67600 57616 68324 57644
rect 74920 57644 74948 57684
rect 75104 57644 75132 57752
rect 78306 57740 78312 57752
rect 78364 57740 78370 57792
rect 84286 57740 84292 57792
rect 84344 57780 84350 57792
rect 88978 57780 88984 57792
rect 84344 57752 88984 57780
rect 84344 57740 84350 57752
rect 88978 57740 88984 57752
rect 89036 57740 89042 57792
rect 92658 57740 92664 57792
rect 92716 57780 92722 57792
rect 126238 57780 126244 57792
rect 92716 57752 126244 57780
rect 92716 57740 92722 57752
rect 126238 57740 126244 57752
rect 126296 57740 126302 57792
rect 126348 57780 126376 57820
rect 126422 57808 126428 57860
rect 126480 57848 126486 57860
rect 133156 57848 133184 57888
rect 133782 57876 133788 57928
rect 133840 57916 133846 57928
rect 139486 57916 139492 57928
rect 133840 57888 139492 57916
rect 133840 57876 133846 57888
rect 139486 57876 139492 57888
rect 139544 57876 139550 57928
rect 141786 57876 141792 57928
rect 141844 57916 141850 57928
rect 218882 57916 218888 57928
rect 141844 57888 218888 57916
rect 141844 57876 141850 57888
rect 218882 57876 218888 57888
rect 218940 57876 218946 57928
rect 218974 57876 218980 57928
rect 219032 57876 219038 57928
rect 220354 57876 220360 57928
rect 220412 57916 220418 57928
rect 225322 57916 225328 57928
rect 220412 57888 225328 57916
rect 220412 57876 220418 57888
rect 225322 57876 225328 57888
rect 225380 57876 225386 57928
rect 226978 57876 226984 57928
rect 227036 57916 227042 57928
rect 300118 57916 300124 57928
rect 227036 57888 300124 57916
rect 227036 57876 227042 57888
rect 300118 57876 300124 57888
rect 300176 57876 300182 57928
rect 136266 57848 136272 57860
rect 126480 57820 128584 57848
rect 133156 57820 136272 57848
rect 126480 57808 126486 57820
rect 128446 57780 128452 57792
rect 126348 57752 128452 57780
rect 128446 57740 128452 57752
rect 128504 57740 128510 57792
rect 128556 57780 128584 57820
rect 136266 57808 136272 57820
rect 136324 57808 136330 57860
rect 137370 57808 137376 57860
rect 137428 57848 137434 57860
rect 137428 57820 218376 57848
rect 137428 57808 137434 57820
rect 142522 57780 142528 57792
rect 128556 57752 142528 57780
rect 142522 57740 142528 57752
rect 142580 57740 142586 57792
rect 216582 57780 216588 57792
rect 142816 57752 216588 57780
rect 77754 57712 77760 57724
rect 74920 57616 75132 57644
rect 75748 57684 77760 57712
rect 67600 57604 67606 57616
rect 27522 57536 27528 57588
rect 27580 57576 27586 57588
rect 66622 57576 66628 57588
rect 27580 57548 66628 57576
rect 27580 57536 27586 57548
rect 66622 57536 66628 57548
rect 66680 57536 66686 57588
rect 70302 57536 70308 57588
rect 70360 57576 70366 57588
rect 75748 57576 75776 57684
rect 77754 57672 77760 57684
rect 77812 57672 77818 57724
rect 84654 57672 84660 57724
rect 84712 57712 84718 57724
rect 86310 57712 86316 57724
rect 84712 57684 86316 57712
rect 84712 57672 84718 57684
rect 86310 57672 86316 57684
rect 86368 57672 86374 57724
rect 88794 57672 88800 57724
rect 88852 57712 88858 57724
rect 103882 57712 103888 57724
rect 88852 57684 103888 57712
rect 88852 57672 88858 57684
rect 103882 57672 103888 57684
rect 103940 57672 103946 57724
rect 113818 57672 113824 57724
rect 113876 57712 113882 57724
rect 113876 57684 128354 57712
rect 113876 57672 113882 57684
rect 80698 57604 80704 57656
rect 80756 57644 80762 57656
rect 81250 57644 81256 57656
rect 80756 57616 81256 57644
rect 80756 57604 80762 57616
rect 81250 57604 81256 57616
rect 81308 57604 81314 57656
rect 82170 57604 82176 57656
rect 82228 57644 82234 57656
rect 82630 57644 82636 57656
rect 82228 57616 82636 57644
rect 82228 57604 82234 57616
rect 82630 57604 82636 57616
rect 82688 57604 82694 57656
rect 83090 57604 83096 57656
rect 83148 57644 83154 57656
rect 84102 57644 84108 57656
rect 83148 57616 84108 57644
rect 83148 57604 83154 57616
rect 84102 57604 84108 57616
rect 84160 57604 84166 57656
rect 85206 57604 85212 57656
rect 85264 57644 85270 57656
rect 86218 57644 86224 57656
rect 85264 57616 86224 57644
rect 85264 57604 85270 57616
rect 86218 57604 86224 57616
rect 86276 57604 86282 57656
rect 86402 57604 86408 57656
rect 86460 57644 86466 57656
rect 86862 57644 86868 57656
rect 86460 57616 86868 57644
rect 86460 57604 86466 57616
rect 86862 57604 86868 57616
rect 86920 57604 86926 57656
rect 89990 57604 89996 57656
rect 90048 57644 90054 57656
rect 90726 57644 90732 57656
rect 90048 57616 90732 57644
rect 90048 57604 90054 57616
rect 90726 57604 90732 57616
rect 90784 57604 90790 57656
rect 91462 57604 91468 57656
rect 91520 57644 91526 57656
rect 92382 57644 92388 57656
rect 91520 57616 92388 57644
rect 91520 57604 91526 57616
rect 92382 57604 92388 57616
rect 92440 57604 92446 57656
rect 93302 57604 93308 57656
rect 93360 57644 93366 57656
rect 127894 57644 127900 57656
rect 93360 57616 127900 57644
rect 93360 57604 93366 57616
rect 127894 57604 127900 57616
rect 127952 57604 127958 57656
rect 127986 57604 127992 57656
rect 128044 57644 128050 57656
rect 128170 57644 128176 57656
rect 128044 57616 128176 57644
rect 128044 57604 128050 57616
rect 128170 57604 128176 57616
rect 128228 57604 128234 57656
rect 128326 57644 128354 57684
rect 135530 57672 135536 57724
rect 135588 57712 135594 57724
rect 142816 57712 142844 57752
rect 216582 57740 216588 57752
rect 216640 57740 216646 57792
rect 216674 57740 216680 57792
rect 216732 57780 216738 57792
rect 218238 57780 218244 57792
rect 216732 57752 218244 57780
rect 216732 57740 216738 57752
rect 218238 57740 218244 57752
rect 218296 57740 218302 57792
rect 161842 57712 161848 57724
rect 135588 57684 142844 57712
rect 147646 57684 161848 57712
rect 135588 57672 135594 57684
rect 137186 57644 137192 57656
rect 128326 57616 137192 57644
rect 137186 57604 137192 57616
rect 137244 57604 137250 57656
rect 138658 57644 138664 57656
rect 137296 57616 138664 57644
rect 70360 57548 75776 57576
rect 70360 57536 70366 57548
rect 75822 57536 75828 57588
rect 75880 57576 75886 57588
rect 78950 57576 78956 57588
rect 75880 57548 78956 57576
rect 75880 57536 75886 57548
rect 78950 57536 78956 57548
rect 79008 57536 79014 57588
rect 81894 57536 81900 57588
rect 81952 57576 81958 57588
rect 82722 57576 82728 57588
rect 81952 57548 82728 57576
rect 81952 57536 81958 57548
rect 82722 57536 82728 57548
rect 82780 57536 82786 57588
rect 85850 57536 85856 57588
rect 85908 57576 85914 57588
rect 86770 57576 86776 57588
rect 85908 57548 86776 57576
rect 85908 57536 85914 57548
rect 86770 57536 86776 57548
rect 86828 57536 86834 57588
rect 89714 57536 89720 57588
rect 89772 57576 89778 57588
rect 91002 57576 91008 57588
rect 89772 57548 91008 57576
rect 89772 57536 89778 57548
rect 91002 57536 91008 57548
rect 91060 57536 91066 57588
rect 94498 57536 94504 57588
rect 94556 57576 94562 57588
rect 95142 57576 95148 57588
rect 94556 57548 95148 57576
rect 94556 57536 94562 57548
rect 95142 57536 95148 57548
rect 95200 57536 95206 57588
rect 95970 57536 95976 57588
rect 96028 57576 96034 57588
rect 96522 57576 96528 57588
rect 96028 57548 96528 57576
rect 96028 57536 96034 57548
rect 96522 57536 96528 57548
rect 96580 57536 96586 57588
rect 97166 57536 97172 57588
rect 97224 57576 97230 57588
rect 97718 57576 97724 57588
rect 97224 57548 97724 57576
rect 97224 57536 97230 57548
rect 97718 57536 97724 57548
rect 97776 57536 97782 57588
rect 98914 57536 98920 57588
rect 98972 57576 98978 57588
rect 99282 57576 99288 57588
rect 98972 57548 99288 57576
rect 98972 57536 98978 57548
rect 99282 57536 99288 57548
rect 99340 57536 99346 57588
rect 104250 57536 104256 57588
rect 104308 57576 104314 57588
rect 131850 57576 131856 57588
rect 104308 57548 131856 57576
rect 104308 57536 104314 57548
rect 131850 57536 131856 57548
rect 131908 57536 131914 57588
rect 132034 57536 132040 57588
rect 132092 57576 132098 57588
rect 137296 57576 137324 57616
rect 138658 57604 138664 57616
rect 138716 57604 138722 57656
rect 142706 57604 142712 57656
rect 142764 57644 142770 57656
rect 147646 57644 147674 57684
rect 161842 57672 161848 57684
rect 161900 57672 161906 57724
rect 167638 57672 167644 57724
rect 167696 57712 167702 57724
rect 168098 57712 168104 57724
rect 167696 57684 168104 57712
rect 167696 57672 167702 57684
rect 168098 57672 168104 57684
rect 168156 57672 168162 57724
rect 169294 57672 169300 57724
rect 169352 57712 169358 57724
rect 169662 57712 169668 57724
rect 169352 57684 169668 57712
rect 169352 57672 169358 57684
rect 169662 57672 169668 57684
rect 169720 57672 169726 57724
rect 171226 57672 171232 57724
rect 171284 57712 171290 57724
rect 172238 57712 172244 57724
rect 171284 57684 172244 57712
rect 171284 57672 171290 57684
rect 172238 57672 172244 57684
rect 172296 57672 172302 57724
rect 172698 57672 172704 57724
rect 172756 57712 172762 57724
rect 173802 57712 173808 57724
rect 172756 57684 173808 57712
rect 172756 57672 172762 57684
rect 173802 57672 173808 57684
rect 173860 57672 173866 57724
rect 174446 57672 174452 57724
rect 174504 57712 174510 57724
rect 175182 57712 175188 57724
rect 174504 57684 175188 57712
rect 174504 57672 174510 57684
rect 175182 57672 175188 57684
rect 175240 57672 175246 57724
rect 175550 57672 175556 57724
rect 175608 57712 175614 57724
rect 176562 57712 176568 57724
rect 175608 57684 176568 57712
rect 175608 57672 175614 57684
rect 176562 57672 176568 57684
rect 176620 57672 176626 57724
rect 177206 57672 177212 57724
rect 177264 57712 177270 57724
rect 177942 57712 177948 57724
rect 177264 57684 177948 57712
rect 177264 57672 177270 57684
rect 177942 57672 177948 57684
rect 178000 57672 178006 57724
rect 178034 57672 178040 57724
rect 178092 57712 178098 57724
rect 179322 57712 179328 57724
rect 178092 57684 179328 57712
rect 178092 57672 178098 57684
rect 179322 57672 179328 57684
rect 179380 57672 179386 57724
rect 180702 57672 180708 57724
rect 180760 57712 180766 57724
rect 180978 57712 180984 57724
rect 180760 57684 180984 57712
rect 180760 57672 180766 57684
rect 180978 57672 180984 57684
rect 181036 57672 181042 57724
rect 181070 57672 181076 57724
rect 181128 57712 181134 57724
rect 181714 57712 181720 57724
rect 181128 57684 181720 57712
rect 181128 57672 181134 57684
rect 181714 57672 181720 57684
rect 181772 57672 181778 57724
rect 182542 57672 182548 57724
rect 182600 57712 182606 57724
rect 183094 57712 183100 57724
rect 182600 57684 183100 57712
rect 182600 57672 182606 57684
rect 183094 57672 183100 57684
rect 183152 57672 183158 57724
rect 183738 57672 183744 57724
rect 183796 57712 183802 57724
rect 184750 57712 184756 57724
rect 183796 57684 184756 57712
rect 183796 57672 183802 57684
rect 184750 57672 184756 57684
rect 184808 57672 184814 57724
rect 186774 57672 186780 57724
rect 186832 57712 186838 57724
rect 187418 57712 187424 57724
rect 186832 57684 187424 57712
rect 186832 57672 186838 57684
rect 187418 57672 187424 57684
rect 187476 57672 187482 57724
rect 187694 57672 187700 57724
rect 187752 57712 187758 57724
rect 188890 57712 188896 57724
rect 187752 57684 188896 57712
rect 187752 57672 187758 57684
rect 188890 57672 188896 57684
rect 188948 57672 188954 57724
rect 189074 57672 189080 57724
rect 189132 57712 189138 57724
rect 190086 57712 190092 57724
rect 189132 57684 190092 57712
rect 189132 57672 189138 57684
rect 190086 57672 190092 57684
rect 190144 57672 190150 57724
rect 190638 57672 190644 57724
rect 190696 57712 190702 57724
rect 191650 57712 191656 57724
rect 190696 57684 191656 57712
rect 190696 57672 190702 57684
rect 191650 57672 191656 57684
rect 191708 57672 191714 57724
rect 192018 57672 192024 57724
rect 192076 57712 192082 57724
rect 192754 57712 192760 57724
rect 192076 57684 192760 57712
rect 192076 57672 192082 57684
rect 192754 57672 192760 57684
rect 192812 57672 192818 57724
rect 194870 57672 194876 57724
rect 194928 57712 194934 57724
rect 195698 57712 195704 57724
rect 194928 57684 195704 57712
rect 194928 57672 194934 57684
rect 195698 57672 195704 57684
rect 195756 57672 195762 57724
rect 196342 57672 196348 57724
rect 196400 57712 196406 57724
rect 196986 57712 196992 57724
rect 196400 57684 196992 57712
rect 196400 57672 196406 57684
rect 196986 57672 196992 57684
rect 197044 57672 197050 57724
rect 197630 57672 197636 57724
rect 197688 57712 197694 57724
rect 198458 57712 198464 57724
rect 197688 57684 198464 57712
rect 197688 57672 197694 57684
rect 198458 57672 198464 57684
rect 198516 57672 198522 57724
rect 199010 57672 199016 57724
rect 199068 57712 199074 57724
rect 199746 57712 199752 57724
rect 199068 57684 199752 57712
rect 199068 57672 199074 57684
rect 199746 57672 199752 57684
rect 199804 57672 199810 57724
rect 200850 57672 200856 57724
rect 200908 57712 200914 57724
rect 201310 57712 201316 57724
rect 200908 57684 201316 57712
rect 200908 57672 200914 57684
rect 201310 57672 201316 57684
rect 201368 57672 201374 57724
rect 201770 57672 201776 57724
rect 201828 57712 201834 57724
rect 202506 57712 202512 57724
rect 201828 57684 202512 57712
rect 201828 57672 201834 57684
rect 202506 57672 202512 57684
rect 202564 57672 202570 57724
rect 203518 57672 203524 57724
rect 203576 57712 203582 57724
rect 203978 57712 203984 57724
rect 203576 57684 203984 57712
rect 203576 57672 203582 57684
rect 203978 57672 203984 57684
rect 204036 57672 204042 57724
rect 205082 57672 205088 57724
rect 205140 57712 205146 57724
rect 205542 57712 205548 57724
rect 205140 57684 205548 57712
rect 205140 57672 205146 57684
rect 205542 57672 205548 57684
rect 205600 57672 205606 57724
rect 206278 57672 206284 57724
rect 206336 57712 206342 57724
rect 206830 57712 206836 57724
rect 206336 57684 206836 57712
rect 206336 57672 206342 57684
rect 206830 57672 206836 57684
rect 206888 57672 206894 57724
rect 207106 57672 207112 57724
rect 207164 57712 207170 57724
rect 208210 57712 208216 57724
rect 207164 57684 208216 57712
rect 207164 57672 207170 57684
rect 208210 57672 208216 57684
rect 208268 57672 208274 57724
rect 208302 57672 208308 57724
rect 208360 57712 208366 57724
rect 216858 57712 216864 57724
rect 208360 57684 216864 57712
rect 208360 57672 208366 57684
rect 216858 57672 216864 57684
rect 216916 57672 216922 57724
rect 218348 57712 218376 57820
rect 219434 57808 219440 57860
rect 219492 57848 219498 57860
rect 225414 57848 225420 57860
rect 219492 57820 225420 57848
rect 219492 57808 219498 57820
rect 225414 57808 225420 57820
rect 225472 57808 225478 57860
rect 269758 57848 269764 57860
rect 231826 57820 269764 57848
rect 218422 57740 218428 57792
rect 218480 57780 218486 57792
rect 221642 57780 221648 57792
rect 218480 57752 221648 57780
rect 218480 57740 218486 57752
rect 221642 57740 221648 57752
rect 221700 57740 221706 57792
rect 223298 57740 223304 57792
rect 223356 57780 223362 57792
rect 231826 57780 231854 57820
rect 269758 57808 269764 57820
rect 269816 57808 269822 57860
rect 223356 57752 231854 57780
rect 223356 57740 223362 57752
rect 221458 57712 221464 57724
rect 218348 57684 221464 57712
rect 221458 57672 221464 57684
rect 221516 57672 221522 57724
rect 221826 57672 221832 57724
rect 221884 57712 221890 57724
rect 226978 57712 226984 57724
rect 221884 57684 226984 57712
rect 221884 57672 221890 57684
rect 226978 57672 226984 57684
rect 227036 57672 227042 57724
rect 142764 57616 147674 57644
rect 142764 57604 142770 57616
rect 148686 57604 148692 57656
rect 148744 57644 148750 57656
rect 347130 57644 347136 57656
rect 148744 57616 347136 57644
rect 148744 57604 148750 57616
rect 347130 57604 347136 57616
rect 347188 57604 347194 57656
rect 132092 57548 137324 57576
rect 132092 57536 132098 57548
rect 140958 57536 140964 57588
rect 141016 57576 141022 57588
rect 141016 57548 147674 57576
rect 141016 57536 141022 57548
rect 24762 57468 24768 57520
rect 24820 57508 24826 57520
rect 66070 57508 66076 57520
rect 24820 57480 66076 57508
rect 24820 57468 24826 57480
rect 66070 57468 66076 57480
rect 66128 57468 66134 57520
rect 66162 57468 66168 57520
rect 66220 57508 66226 57520
rect 76558 57508 76564 57520
rect 66220 57480 76564 57508
rect 66220 57468 66226 57480
rect 76558 57468 76564 57480
rect 76616 57468 76622 57520
rect 82814 57468 82820 57520
rect 82872 57508 82878 57520
rect 84010 57508 84016 57520
rect 82872 57480 84016 57508
rect 82872 57468 82878 57480
rect 84010 57468 84016 57480
rect 84068 57468 84074 57520
rect 87322 57468 87328 57520
rect 87380 57508 87386 57520
rect 88150 57508 88156 57520
rect 87380 57480 88156 57508
rect 87380 57468 87386 57480
rect 88150 57468 88156 57480
rect 88208 57468 88214 57520
rect 88518 57468 88524 57520
rect 88576 57508 88582 57520
rect 89530 57508 89536 57520
rect 88576 57480 89536 57508
rect 88576 57468 88582 57480
rect 89530 57468 89536 57480
rect 89588 57468 89594 57520
rect 90634 57468 90640 57520
rect 90692 57508 90698 57520
rect 90910 57508 90916 57520
rect 90692 57480 90916 57508
rect 90692 57468 90698 57480
rect 90910 57468 90916 57480
rect 90968 57468 90974 57520
rect 93026 57468 93032 57520
rect 93084 57508 93090 57520
rect 93670 57508 93676 57520
rect 93084 57480 93676 57508
rect 93084 57468 93090 57480
rect 93670 57468 93676 57480
rect 93728 57468 93734 57520
rect 93854 57468 93860 57520
rect 93912 57508 93918 57520
rect 95050 57508 95056 57520
rect 93912 57480 95056 57508
rect 93912 57468 93918 57480
rect 95050 57468 95056 57480
rect 95108 57468 95114 57520
rect 95694 57468 95700 57520
rect 95752 57508 95758 57520
rect 96338 57508 96344 57520
rect 95752 57480 96344 57508
rect 95752 57468 95758 57480
rect 96338 57468 96344 57480
rect 96396 57468 96402 57520
rect 96614 57468 96620 57520
rect 96672 57508 96678 57520
rect 97626 57508 97632 57520
rect 96672 57480 97632 57508
rect 96672 57468 96678 57480
rect 97626 57468 97632 57480
rect 97684 57468 97690 57520
rect 104158 57468 104164 57520
rect 104216 57508 104222 57520
rect 104216 57480 132172 57508
rect 104216 57468 104222 57480
rect 26142 57400 26148 57452
rect 26200 57440 26206 57452
rect 66346 57440 66352 57452
rect 26200 57412 66352 57440
rect 26200 57400 26206 57412
rect 66346 57400 66352 57412
rect 66404 57400 66410 57452
rect 70210 57400 70216 57452
rect 70268 57440 70274 57452
rect 75086 57440 75092 57452
rect 70268 57412 75092 57440
rect 70268 57400 70274 57412
rect 75086 57400 75092 57412
rect 75144 57400 75150 57452
rect 75178 57400 75184 57452
rect 75236 57440 75242 57452
rect 78582 57440 78588 57452
rect 75236 57412 78588 57440
rect 75236 57400 75242 57412
rect 78582 57400 78588 57412
rect 78640 57400 78646 57452
rect 81618 57400 81624 57452
rect 81676 57440 81682 57452
rect 82446 57440 82452 57452
rect 81676 57412 82452 57440
rect 81676 57400 81682 57412
rect 82446 57400 82452 57412
rect 82504 57400 82510 57452
rect 87598 57400 87604 57452
rect 87656 57440 87662 57452
rect 88242 57440 88248 57452
rect 87656 57412 88248 57440
rect 87656 57400 87662 57412
rect 88242 57400 88248 57412
rect 88300 57400 88306 57452
rect 96890 57400 96896 57452
rect 96948 57440 96954 57452
rect 97810 57440 97816 57452
rect 96948 57412 97816 57440
rect 96948 57400 96954 57412
rect 97810 57400 97816 57412
rect 97868 57400 97874 57452
rect 98086 57400 98092 57452
rect 98144 57440 98150 57452
rect 99282 57440 99288 57452
rect 98144 57412 99288 57440
rect 98144 57400 98150 57412
rect 99282 57400 99288 57412
rect 99340 57400 99346 57452
rect 103974 57400 103980 57452
rect 104032 57440 104038 57452
rect 132034 57440 132040 57452
rect 104032 57412 132040 57440
rect 104032 57400 104038 57412
rect 132034 57400 132040 57412
rect 132092 57400 132098 57452
rect 132144 57440 132172 57480
rect 132954 57468 132960 57520
rect 133012 57508 133018 57520
rect 137278 57508 137284 57520
rect 133012 57480 137284 57508
rect 133012 57468 133018 57480
rect 137278 57468 137284 57480
rect 137336 57468 137342 57520
rect 137370 57468 137376 57520
rect 137428 57508 137434 57520
rect 141602 57508 141608 57520
rect 137428 57480 141608 57508
rect 137428 57468 137434 57480
rect 141602 57468 141608 57480
rect 141660 57468 141666 57520
rect 142522 57468 142528 57520
rect 142580 57508 142586 57520
rect 146846 57508 146852 57520
rect 142580 57480 146852 57508
rect 142580 57468 142586 57480
rect 146846 57468 146852 57480
rect 146904 57468 146910 57520
rect 147646 57508 147674 57548
rect 148410 57536 148416 57588
rect 148468 57576 148474 57588
rect 347038 57576 347044 57588
rect 148468 57548 347044 57576
rect 148468 57536 148474 57548
rect 347038 57536 347044 57548
rect 347096 57536 347102 57588
rect 148318 57508 148324 57520
rect 147646 57480 148324 57508
rect 148318 57468 148324 57480
rect 148376 57468 148382 57520
rect 149606 57468 149612 57520
rect 149664 57508 149670 57520
rect 353294 57508 353300 57520
rect 149664 57480 353300 57508
rect 149664 57468 149670 57480
rect 353294 57468 353300 57480
rect 353352 57468 353358 57520
rect 138014 57440 138020 57452
rect 132144 57412 138020 57440
rect 138014 57400 138020 57412
rect 138072 57400 138078 57452
rect 143626 57400 143632 57452
rect 143684 57440 143690 57452
rect 165706 57440 165712 57452
rect 143684 57412 165712 57440
rect 143684 57400 143690 57412
rect 165706 57400 165712 57412
rect 165764 57400 165770 57452
rect 167178 57400 167184 57452
rect 167236 57440 167242 57452
rect 168190 57440 168196 57452
rect 167236 57412 168196 57440
rect 167236 57400 167242 57412
rect 168190 57400 168196 57412
rect 168248 57400 168254 57452
rect 168834 57400 168840 57452
rect 168892 57440 168898 57452
rect 169570 57440 169576 57452
rect 168892 57412 169576 57440
rect 168892 57400 168898 57412
rect 169570 57400 169576 57412
rect 169628 57400 169634 57452
rect 174170 57400 174176 57452
rect 174228 57440 174234 57452
rect 175090 57440 175096 57452
rect 174228 57412 175096 57440
rect 174228 57400 174234 57412
rect 175090 57400 175096 57412
rect 175148 57400 175154 57452
rect 175366 57400 175372 57452
rect 175424 57440 175430 57452
rect 176470 57440 176476 57452
rect 175424 57412 176476 57440
rect 175424 57400 175430 57412
rect 176470 57400 176476 57412
rect 176528 57400 176534 57452
rect 178126 57400 178132 57452
rect 178184 57440 178190 57452
rect 179230 57440 179236 57452
rect 178184 57412 179236 57440
rect 178184 57400 178190 57412
rect 179230 57400 179236 57412
rect 179288 57400 179294 57452
rect 179708 57412 185716 57440
rect 17862 57332 17868 57384
rect 17920 57372 17926 57384
rect 17920 57344 57744 57372
rect 17920 57332 17926 57344
rect 6822 57264 6828 57316
rect 6880 57304 6886 57316
rect 57606 57304 57612 57316
rect 6880 57276 57612 57304
rect 6880 57264 6886 57276
rect 57606 57264 57612 57276
rect 57664 57264 57670 57316
rect 57716 57304 57744 57344
rect 57790 57332 57796 57384
rect 57848 57372 57854 57384
rect 61562 57372 61568 57384
rect 57848 57344 61568 57372
rect 57848 57332 57854 57344
rect 61562 57332 61568 57344
rect 61620 57332 61626 57384
rect 64230 57372 64236 57384
rect 61672 57344 64236 57372
rect 61672 57304 61700 57344
rect 64230 57332 64236 57344
rect 64288 57332 64294 57384
rect 64782 57332 64788 57384
rect 64840 57372 64846 57384
rect 76190 57372 76196 57384
rect 64840 57344 76196 57372
rect 64840 57332 64846 57344
rect 76190 57332 76196 57344
rect 76248 57332 76254 57384
rect 83366 57332 83372 57384
rect 83424 57372 83430 57384
rect 92658 57372 92664 57384
rect 83424 57344 92664 57372
rect 83424 57332 83430 57344
rect 92658 57332 92664 57344
rect 92716 57332 92722 57384
rect 97534 57332 97540 57384
rect 97592 57372 97598 57384
rect 147766 57372 147772 57384
rect 97592 57344 147772 57372
rect 97592 57332 97598 57344
rect 147766 57332 147772 57344
rect 147824 57332 147830 57384
rect 148134 57332 148140 57384
rect 148192 57372 148198 57384
rect 152550 57372 152556 57384
rect 148192 57344 152556 57372
rect 148192 57332 148198 57344
rect 152550 57332 152556 57344
rect 152608 57332 152614 57384
rect 152642 57332 152648 57384
rect 152700 57372 152706 57384
rect 153102 57372 153108 57384
rect 152700 57344 153108 57372
rect 152700 57332 152706 57344
rect 153102 57332 153108 57344
rect 153160 57332 153166 57384
rect 153838 57332 153844 57384
rect 153896 57372 153902 57384
rect 154298 57372 154304 57384
rect 153896 57344 154304 57372
rect 153896 57332 153902 57344
rect 154298 57332 154304 57344
rect 154356 57332 154362 57384
rect 155034 57332 155040 57384
rect 155092 57372 155098 57384
rect 155678 57372 155684 57384
rect 155092 57344 155684 57372
rect 155092 57332 155098 57344
rect 155678 57332 155684 57344
rect 155736 57332 155742 57384
rect 156506 57332 156512 57384
rect 156564 57372 156570 57384
rect 157058 57372 157064 57384
rect 156564 57344 157064 57372
rect 156564 57332 156570 57344
rect 157058 57332 157064 57344
rect 157116 57332 157122 57384
rect 157306 57344 168328 57372
rect 57716 57276 61700 57304
rect 62022 57264 62028 57316
rect 62080 57304 62086 57316
rect 75638 57304 75644 57316
rect 62080 57276 75644 57304
rect 62080 57264 62086 57276
rect 75638 57264 75644 57276
rect 75696 57264 75702 57316
rect 86126 57264 86132 57316
rect 86184 57304 86190 57316
rect 101306 57304 101312 57316
rect 86184 57276 101312 57304
rect 86184 57264 86190 57276
rect 101306 57264 101312 57276
rect 101364 57264 101370 57316
rect 102594 57264 102600 57316
rect 102652 57304 102658 57316
rect 157306 57304 157334 57344
rect 102652 57276 157334 57304
rect 102652 57264 102658 57276
rect 166994 57264 167000 57316
rect 167052 57304 167058 57316
rect 168190 57304 168196 57316
rect 167052 57276 168196 57304
rect 167052 57264 167058 57276
rect 168190 57264 168196 57276
rect 168248 57264 168254 57316
rect 168300 57304 168328 57344
rect 168466 57332 168472 57384
rect 168524 57372 168530 57384
rect 169478 57372 169484 57384
rect 168524 57344 169484 57372
rect 168524 57332 168530 57344
rect 169478 57332 169484 57344
rect 169536 57332 169542 57384
rect 178678 57332 178684 57384
rect 178736 57372 178742 57384
rect 179708 57372 179736 57412
rect 178736 57344 179736 57372
rect 178736 57332 178742 57344
rect 180334 57332 180340 57384
rect 180392 57372 180398 57384
rect 180392 57344 185440 57372
rect 180392 57332 180398 57344
rect 168742 57304 168748 57316
rect 168300 57276 168748 57304
rect 168742 57264 168748 57276
rect 168800 57264 168806 57316
rect 179598 57264 179604 57316
rect 179656 57304 179662 57316
rect 180702 57304 180708 57316
rect 179656 57276 180708 57304
rect 179656 57264 179662 57276
rect 180702 57264 180708 57276
rect 180760 57264 180766 57316
rect 180794 57264 180800 57316
rect 180852 57304 180858 57316
rect 183554 57304 183560 57316
rect 180852 57276 183560 57304
rect 180852 57264 180858 57276
rect 183554 57264 183560 57276
rect 183612 57264 183618 57316
rect 3970 57196 3976 57248
rect 4028 57236 4034 57248
rect 60642 57236 60648 57248
rect 4028 57208 60648 57236
rect 4028 57196 4034 57208
rect 60642 57196 60648 57208
rect 60700 57196 60706 57248
rect 60826 57196 60832 57248
rect 60884 57236 60890 57248
rect 74994 57236 75000 57248
rect 60884 57208 75000 57236
rect 60884 57196 60890 57208
rect 74994 57196 75000 57208
rect 75052 57196 75058 57248
rect 77110 57236 77116 57248
rect 75840 57208 77116 57236
rect 35802 57128 35808 57180
rect 35860 57168 35866 57180
rect 68738 57168 68744 57180
rect 35860 57140 68744 57168
rect 35860 57128 35866 57140
rect 68738 57128 68744 57140
rect 68796 57128 68802 57180
rect 68922 57128 68928 57180
rect 68980 57168 68986 57180
rect 75840 57168 75868 57208
rect 77110 57196 77116 57208
rect 77168 57196 77174 57248
rect 87046 57196 87052 57248
rect 87104 57236 87110 57248
rect 102962 57236 102968 57248
rect 87104 57208 102968 57236
rect 87104 57196 87110 57208
rect 102962 57196 102968 57208
rect 103020 57196 103026 57248
rect 171594 57236 171600 57248
rect 114020 57208 171600 57236
rect 68980 57140 75868 57168
rect 68980 57128 68986 57140
rect 76558 57128 76564 57180
rect 76616 57168 76622 57180
rect 78030 57168 78036 57180
rect 76616 57140 78036 57168
rect 76616 57128 76622 57140
rect 78030 57128 78036 57140
rect 78088 57128 78094 57180
rect 91186 57128 91192 57180
rect 91244 57168 91250 57180
rect 97258 57168 97264 57180
rect 91244 57140 97264 57168
rect 91244 57128 91250 57140
rect 97258 57128 97264 57140
rect 97316 57128 97322 57180
rect 98362 57128 98368 57180
rect 98420 57168 98426 57180
rect 99006 57168 99012 57180
rect 98420 57140 99012 57168
rect 98420 57128 98426 57140
rect 99006 57128 99012 57140
rect 99064 57128 99070 57180
rect 103514 57128 103520 57180
rect 103572 57168 103578 57180
rect 103572 57140 106136 57168
rect 103572 57128 103578 57140
rect 41322 57060 41328 57112
rect 41380 57100 41386 57112
rect 70118 57100 70124 57112
rect 41380 57072 70124 57100
rect 41380 57060 41386 57072
rect 70118 57060 70124 57072
rect 70176 57060 70182 57112
rect 94958 57060 94964 57112
rect 95016 57100 95022 57112
rect 104158 57100 104164 57112
rect 95016 57072 104164 57100
rect 95016 57060 95022 57072
rect 104158 57060 104164 57072
rect 104216 57060 104222 57112
rect 43438 56992 43444 57044
rect 43496 57032 43502 57044
rect 70486 57032 70492 57044
rect 43496 57004 70492 57032
rect 43496 56992 43502 57004
rect 70486 56992 70492 57004
rect 70544 56992 70550 57044
rect 74718 57032 74724 57044
rect 74506 57004 74724 57032
rect 46842 56924 46848 56976
rect 46900 56964 46906 56976
rect 71682 56964 71688 56976
rect 46900 56936 71688 56964
rect 46900 56924 46906 56936
rect 71682 56924 71688 56936
rect 71740 56924 71746 56976
rect 48222 56856 48228 56908
rect 48280 56896 48286 56908
rect 72050 56896 72056 56908
rect 48280 56868 72056 56896
rect 48280 56856 48286 56868
rect 72050 56856 72056 56868
rect 72108 56856 72114 56908
rect 72142 56856 72148 56908
rect 72200 56896 72206 56908
rect 74166 56896 74172 56908
rect 72200 56868 74172 56896
rect 72200 56856 72206 56868
rect 74166 56856 74172 56868
rect 74224 56856 74230 56908
rect 53742 56788 53748 56840
rect 53800 56828 53806 56840
rect 73522 56828 73528 56840
rect 53800 56800 73528 56828
rect 53800 56788 53806 56800
rect 73522 56788 73528 56800
rect 73580 56788 73586 56840
rect 55122 56720 55128 56772
rect 55180 56760 55186 56772
rect 73798 56760 73804 56772
rect 55180 56732 73804 56760
rect 55180 56720 55186 56732
rect 73798 56720 73804 56732
rect 73856 56720 73862 56772
rect 59262 56652 59268 56704
rect 59320 56692 59326 56704
rect 74506 56692 74534 57004
rect 74718 56992 74724 57004
rect 74776 56992 74782 57044
rect 77202 56992 77208 57044
rect 77260 57032 77266 57044
rect 79226 57032 79232 57044
rect 77260 57004 79232 57032
rect 77260 56992 77266 57004
rect 79226 56992 79232 57004
rect 79284 56992 79290 57044
rect 84930 56992 84936 57044
rect 84988 57032 84994 57044
rect 87598 57032 87604 57044
rect 84988 57004 87604 57032
rect 84988 56992 84994 57004
rect 87598 56992 87604 57004
rect 87656 56992 87662 57044
rect 92290 56992 92296 57044
rect 92348 57032 92354 57044
rect 106108 57032 106136 57140
rect 106182 57060 106188 57112
rect 106240 57100 106246 57112
rect 113818 57100 113824 57112
rect 106240 57072 113824 57100
rect 106240 57060 106246 57072
rect 113818 57060 113824 57072
rect 113876 57060 113882 57112
rect 114020 57032 114048 57208
rect 171594 57196 171600 57208
rect 171652 57196 171658 57248
rect 176838 57196 176844 57248
rect 176896 57236 176902 57248
rect 180426 57236 180432 57248
rect 176896 57208 180432 57236
rect 176896 57196 176902 57208
rect 180426 57196 180432 57208
rect 180484 57196 180490 57248
rect 181346 57196 181352 57248
rect 181404 57236 181410 57248
rect 181990 57236 181996 57248
rect 181404 57208 181996 57236
rect 181404 57196 181410 57208
rect 181990 57196 181996 57208
rect 182048 57196 182054 57248
rect 182266 57196 182272 57248
rect 182324 57236 182330 57248
rect 183278 57236 183284 57248
rect 182324 57208 183284 57236
rect 182324 57196 182330 57208
rect 183278 57196 183284 57208
rect 183336 57196 183342 57248
rect 185412 57236 185440 57344
rect 185688 57304 185716 57412
rect 186498 57400 186504 57452
rect 186556 57440 186562 57452
rect 187510 57440 187516 57452
rect 186556 57412 187516 57440
rect 186556 57400 186562 57412
rect 187510 57400 187516 57412
rect 187568 57400 187574 57452
rect 187602 57400 187608 57452
rect 187660 57440 187666 57452
rect 187660 57412 190224 57440
rect 187660 57400 187666 57412
rect 190196 57372 190224 57412
rect 190362 57400 190368 57452
rect 190420 57440 190426 57452
rect 411898 57440 411904 57452
rect 190420 57412 411904 57440
rect 190420 57400 190426 57412
rect 411898 57400 411904 57412
rect 411956 57400 411962 57452
rect 418798 57372 418804 57384
rect 190196 57344 418804 57372
rect 418798 57332 418804 57344
rect 418856 57332 418862 57384
rect 425698 57304 425704 57316
rect 185688 57276 425704 57304
rect 425698 57264 425704 57276
rect 425756 57264 425762 57316
rect 429838 57236 429844 57248
rect 185412 57208 429844 57236
rect 429838 57196 429844 57208
rect 429896 57196 429902 57248
rect 114278 57128 114284 57180
rect 114336 57168 114342 57180
rect 146386 57168 146392 57180
rect 114336 57140 146392 57168
rect 114336 57128 114342 57140
rect 146386 57128 146392 57140
rect 146444 57128 146450 57180
rect 151998 57128 152004 57180
rect 152056 57168 152062 57180
rect 153010 57168 153016 57180
rect 152056 57140 153016 57168
rect 152056 57128 152062 57140
rect 153010 57128 153016 57140
rect 153068 57128 153074 57180
rect 153470 57128 153476 57180
rect 153528 57168 153534 57180
rect 154206 57168 154212 57180
rect 153528 57140 154212 57168
rect 153528 57128 153534 57140
rect 154206 57128 154212 57140
rect 154264 57128 154270 57180
rect 154758 57128 154764 57180
rect 154816 57168 154822 57180
rect 155862 57168 155868 57180
rect 154816 57140 155868 57168
rect 154816 57128 154822 57140
rect 155862 57128 155868 57140
rect 155920 57128 155926 57180
rect 155954 57128 155960 57180
rect 156012 57168 156018 57180
rect 156874 57168 156880 57180
rect 156012 57140 156880 57168
rect 156012 57128 156018 57140
rect 156874 57128 156880 57140
rect 156932 57128 156938 57180
rect 157334 57128 157340 57180
rect 157392 57168 157398 57180
rect 216674 57168 216680 57180
rect 157392 57140 216680 57168
rect 157392 57128 157398 57140
rect 216674 57128 216680 57140
rect 216732 57128 216738 57180
rect 218698 57168 218704 57180
rect 216784 57140 218704 57168
rect 117590 57060 117596 57112
rect 117648 57100 117654 57112
rect 118510 57100 118516 57112
rect 117648 57072 118516 57100
rect 117648 57060 117654 57072
rect 118510 57060 118516 57072
rect 118568 57060 118574 57112
rect 143534 57100 143540 57112
rect 118666 57072 143540 57100
rect 92348 57004 104204 57032
rect 106108 57004 114048 57032
rect 92348 56992 92354 57004
rect 95326 56924 95332 56976
rect 95384 56964 95390 56976
rect 102778 56964 102784 56976
rect 95384 56936 102784 56964
rect 95384 56924 95390 56936
rect 102778 56924 102784 56936
rect 102836 56924 102842 56976
rect 104176 56964 104204 57004
rect 104176 56936 109034 56964
rect 94222 56856 94228 56908
rect 94280 56896 94286 56908
rect 104250 56896 104256 56908
rect 94280 56868 104256 56896
rect 94280 56856 94286 56868
rect 104250 56856 104256 56868
rect 104308 56856 104314 56908
rect 80974 56788 80980 56840
rect 81032 56828 81038 56840
rect 83090 56828 83096 56840
rect 81032 56800 83096 56828
rect 81032 56788 81038 56800
rect 83090 56788 83096 56800
rect 83148 56788 83154 56840
rect 105262 56720 105268 56772
rect 105320 56760 105326 56772
rect 106182 56760 106188 56772
rect 105320 56732 106188 56760
rect 105320 56720 105326 56732
rect 106182 56720 106188 56732
rect 106240 56720 106246 56772
rect 59320 56664 74534 56692
rect 59320 56652 59326 56664
rect 99558 56652 99564 56704
rect 99616 56692 99622 56704
rect 100662 56692 100668 56704
rect 99616 56664 100668 56692
rect 99616 56652 99622 56664
rect 100662 56652 100668 56664
rect 100720 56652 100726 56704
rect 101122 56652 101128 56704
rect 101180 56692 101186 56704
rect 101858 56692 101864 56704
rect 101180 56664 101864 56692
rect 101180 56652 101186 56664
rect 101858 56652 101864 56664
rect 101916 56652 101922 56704
rect 102318 56652 102324 56704
rect 102376 56692 102382 56704
rect 103054 56692 103060 56704
rect 102376 56664 103060 56692
rect 102376 56652 102382 56664
rect 103054 56652 103060 56664
rect 103112 56652 103118 56704
rect 104342 56652 104348 56704
rect 104400 56692 104406 56704
rect 104802 56692 104808 56704
rect 104400 56664 104808 56692
rect 104400 56652 104406 56664
rect 104802 56652 104808 56664
rect 104860 56652 104866 56704
rect 104986 56652 104992 56704
rect 105044 56692 105050 56704
rect 105814 56692 105820 56704
rect 105044 56664 105820 56692
rect 105044 56652 105050 56664
rect 105814 56652 105820 56664
rect 105872 56652 105878 56704
rect 106458 56652 106464 56704
rect 106516 56692 106522 56704
rect 107562 56692 107568 56704
rect 106516 56664 107568 56692
rect 106516 56652 106522 56664
rect 107562 56652 107568 56664
rect 107620 56652 107626 56704
rect 57238 56584 57244 56636
rect 57296 56624 57302 56636
rect 72142 56624 72148 56636
rect 57296 56596 72148 56624
rect 57296 56584 57302 56596
rect 72142 56584 72148 56596
rect 72200 56584 72206 56636
rect 72418 56584 72424 56636
rect 72476 56624 72482 56636
rect 75914 56624 75920 56636
rect 72476 56596 75920 56624
rect 72476 56584 72482 56596
rect 75914 56584 75920 56596
rect 75972 56584 75978 56636
rect 98730 56584 98736 56636
rect 98788 56624 98794 56636
rect 99190 56624 99196 56636
rect 98788 56596 99196 56624
rect 98788 56584 98794 56596
rect 99190 56584 99196 56596
rect 99248 56584 99254 56636
rect 99926 56584 99932 56636
rect 99984 56624 99990 56636
rect 100386 56624 100392 56636
rect 99984 56596 100392 56624
rect 99984 56584 99990 56596
rect 100386 56584 100392 56596
rect 100444 56584 100450 56636
rect 101674 56584 101680 56636
rect 101732 56624 101738 56636
rect 102042 56624 102048 56636
rect 101732 56596 102048 56624
rect 101732 56584 101738 56596
rect 102042 56584 102048 56596
rect 102100 56584 102106 56636
rect 102870 56584 102876 56636
rect 102928 56624 102934 56636
rect 103422 56624 103428 56636
rect 102928 56596 103428 56624
rect 102928 56584 102934 56596
rect 103422 56584 103428 56596
rect 103480 56584 103486 56636
rect 104066 56584 104072 56636
rect 104124 56624 104130 56636
rect 104526 56624 104532 56636
rect 104124 56596 104532 56624
rect 104124 56584 104130 56596
rect 104526 56584 104532 56596
rect 104584 56584 104590 56636
rect 105538 56584 105544 56636
rect 105596 56624 105602 56636
rect 106090 56624 106096 56636
rect 105596 56596 106096 56624
rect 105596 56584 105602 56596
rect 106090 56584 106096 56596
rect 106148 56584 106154 56636
rect 106734 56584 106740 56636
rect 106792 56624 106798 56636
rect 107470 56624 107476 56636
rect 106792 56596 107476 56624
rect 106792 56584 106798 56596
rect 107470 56584 107476 56596
rect 107528 56584 107534 56636
rect 107654 56584 107660 56636
rect 107712 56624 107718 56636
rect 108482 56624 108488 56636
rect 107712 56596 108488 56624
rect 107712 56584 107718 56596
rect 108482 56584 108488 56596
rect 108540 56584 108546 56636
rect 109006 56624 109034 56936
rect 113358 56924 113364 56976
rect 113416 56964 113422 56976
rect 113416 56936 118464 56964
rect 113416 56924 113422 56936
rect 115474 56856 115480 56908
rect 115532 56896 115538 56908
rect 115842 56896 115848 56908
rect 115532 56868 115848 56896
rect 115532 56856 115538 56868
rect 115842 56856 115848 56868
rect 115900 56856 115906 56908
rect 118436 56896 118464 56936
rect 118666 56896 118694 57072
rect 143534 57060 143540 57072
rect 143592 57060 143598 57112
rect 146294 57060 146300 57112
rect 146352 57100 146358 57112
rect 155126 57100 155132 57112
rect 146352 57072 155132 57100
rect 146352 57060 146358 57072
rect 155126 57060 155132 57072
rect 155184 57060 155190 57112
rect 156230 57060 156236 57112
rect 156288 57100 156294 57112
rect 157242 57100 157248 57112
rect 156288 57072 157248 57100
rect 156288 57060 156294 57072
rect 157242 57060 157248 57072
rect 157300 57060 157306 57112
rect 216784 57100 216812 57140
rect 218698 57128 218704 57140
rect 218756 57128 218762 57180
rect 218974 57128 218980 57180
rect 219032 57168 219038 57180
rect 221550 57168 221556 57180
rect 219032 57140 221556 57168
rect 219032 57128 219038 57140
rect 221550 57128 221556 57140
rect 221608 57128 221614 57180
rect 162136 57072 216812 57100
rect 121730 56992 121736 57044
rect 121788 57032 121794 57044
rect 127710 57032 127716 57044
rect 121788 57004 127716 57032
rect 121788 56992 121794 57004
rect 127710 56992 127716 57004
rect 127768 56992 127774 57044
rect 128446 56992 128452 57044
rect 128504 57032 128510 57044
rect 136634 57032 136640 57044
rect 128504 57004 136640 57032
rect 128504 56992 128510 57004
rect 136634 56992 136640 57004
rect 136692 56992 136698 57044
rect 140038 56992 140044 57044
rect 140096 57032 140102 57044
rect 140096 57004 147674 57032
rect 140096 56992 140102 57004
rect 122650 56924 122656 56976
rect 122708 56964 122714 56976
rect 127802 56964 127808 56976
rect 122708 56936 127808 56964
rect 122708 56924 122714 56936
rect 127802 56924 127808 56936
rect 127860 56924 127866 56976
rect 144178 56964 144184 56976
rect 128188 56936 144184 56964
rect 124858 56896 124864 56908
rect 118436 56868 118694 56896
rect 120092 56868 124864 56896
rect 109494 56788 109500 56840
rect 109552 56828 109558 56840
rect 110230 56828 110236 56840
rect 109552 56800 110236 56828
rect 109552 56788 109558 56800
rect 110230 56788 110236 56800
rect 110288 56788 110294 56840
rect 110690 56788 110696 56840
rect 110748 56828 110754 56840
rect 111702 56828 111708 56840
rect 110748 56800 111708 56828
rect 110748 56788 110754 56800
rect 111702 56788 111708 56800
rect 111760 56788 111766 56840
rect 111886 56788 111892 56840
rect 111944 56828 111950 56840
rect 112898 56828 112904 56840
rect 111944 56800 112904 56828
rect 111944 56788 111950 56800
rect 112898 56788 112904 56800
rect 112956 56788 112962 56840
rect 113726 56788 113732 56840
rect 113784 56828 113790 56840
rect 120092 56828 120120 56868
rect 124858 56856 124864 56868
rect 124916 56856 124922 56908
rect 113784 56800 120120 56828
rect 113784 56788 113790 56800
rect 123570 56788 123576 56840
rect 123628 56828 123634 56840
rect 123628 56800 125594 56828
rect 123628 56788 123634 56800
rect 109770 56720 109776 56772
rect 109828 56760 109834 56772
rect 110322 56760 110328 56772
rect 109828 56732 110328 56760
rect 109828 56720 109834 56732
rect 110322 56720 110328 56732
rect 110380 56720 110386 56772
rect 110414 56720 110420 56772
rect 110472 56760 110478 56772
rect 111426 56760 111432 56772
rect 110472 56732 111432 56760
rect 110472 56720 110478 56732
rect 111426 56720 111432 56732
rect 111484 56720 111490 56772
rect 112162 56720 112168 56772
rect 112220 56760 112226 56772
rect 112990 56760 112996 56772
rect 112220 56732 112996 56760
rect 112220 56720 112226 56732
rect 112990 56720 112996 56732
rect 113048 56720 113054 56772
rect 114554 56720 114560 56772
rect 114612 56760 114618 56772
rect 115474 56760 115480 56772
rect 114612 56732 115480 56760
rect 114612 56720 114618 56732
rect 115474 56720 115480 56732
rect 115532 56720 115538 56772
rect 116670 56720 116676 56772
rect 116728 56760 116734 56772
rect 117038 56760 117044 56772
rect 116728 56732 117044 56760
rect 116728 56720 116734 56732
rect 117038 56720 117044 56732
rect 117096 56720 117102 56772
rect 120258 56720 120264 56772
rect 120316 56760 120322 56772
rect 121270 56760 121276 56772
rect 120316 56732 121276 56760
rect 120316 56720 120322 56732
rect 121270 56720 121276 56732
rect 121328 56720 121334 56772
rect 109218 56652 109224 56704
rect 109276 56692 109282 56704
rect 109954 56692 109960 56704
rect 109276 56664 109960 56692
rect 109276 56652 109282 56664
rect 109954 56652 109960 56664
rect 110012 56652 110018 56704
rect 110966 56652 110972 56704
rect 111024 56692 111030 56704
rect 111518 56692 111524 56704
rect 111024 56664 111524 56692
rect 111024 56652 111030 56664
rect 111518 56652 111524 56664
rect 111576 56652 111582 56704
rect 112714 56652 112720 56704
rect 112772 56692 112778 56704
rect 113082 56692 113088 56704
rect 112772 56664 113088 56692
rect 112772 56652 112778 56664
rect 113082 56652 113088 56664
rect 113140 56652 113146 56704
rect 113634 56652 113640 56704
rect 113692 56692 113698 56704
rect 114462 56692 114468 56704
rect 113692 56664 114468 56692
rect 113692 56652 113698 56664
rect 114462 56652 114468 56664
rect 114520 56652 114526 56704
rect 114830 56652 114836 56704
rect 114888 56692 114894 56704
rect 115566 56692 115572 56704
rect 114888 56664 115572 56692
rect 114888 56652 114894 56664
rect 115566 56652 115572 56664
rect 115624 56652 115630 56704
rect 116394 56652 116400 56704
rect 116452 56692 116458 56704
rect 116854 56692 116860 56704
rect 116452 56664 116860 56692
rect 116452 56652 116458 56664
rect 116854 56652 116860 56664
rect 116912 56652 116918 56704
rect 125566 56692 125594 56800
rect 127710 56788 127716 56840
rect 127768 56828 127774 56840
rect 128188 56828 128216 56936
rect 144178 56924 144184 56936
rect 144236 56924 144242 56976
rect 128354 56856 128360 56908
rect 128412 56896 128418 56908
rect 129366 56896 129372 56908
rect 128412 56868 129372 56896
rect 128412 56856 128418 56868
rect 129366 56856 129372 56868
rect 129424 56856 129430 56908
rect 131850 56856 131856 56908
rect 131908 56896 131914 56908
rect 135346 56896 135352 56908
rect 131908 56868 135352 56896
rect 131908 56856 131914 56868
rect 135346 56856 135352 56868
rect 135404 56856 135410 56908
rect 139118 56856 139124 56908
rect 139176 56896 139182 56908
rect 146110 56896 146116 56908
rect 139176 56868 146116 56896
rect 139176 56856 139182 56868
rect 146110 56856 146116 56868
rect 146168 56856 146174 56908
rect 147646 56896 147674 57004
rect 152550 56992 152556 57044
rect 152608 57032 152614 57044
rect 159358 57032 159364 57044
rect 152608 57004 159364 57032
rect 152608 56992 152614 57004
rect 159358 56992 159364 57004
rect 159416 56992 159422 57044
rect 149146 56924 149152 56976
rect 149204 56964 149210 56976
rect 150158 56964 150164 56976
rect 149204 56936 150164 56964
rect 149204 56924 149210 56936
rect 150158 56924 150164 56936
rect 150216 56924 150222 56976
rect 155310 56924 155316 56976
rect 155368 56964 155374 56976
rect 162136 56964 162164 57072
rect 216858 57060 216864 57112
rect 216916 57100 216922 57112
rect 225690 57100 225696 57112
rect 216916 57072 225696 57100
rect 216916 57060 216922 57072
rect 225690 57060 225696 57072
rect 225748 57060 225754 57112
rect 155368 56936 162164 56964
rect 162964 57004 217272 57032
rect 155368 56924 155374 56936
rect 158806 56896 158812 56908
rect 147646 56868 158812 56896
rect 158806 56856 158812 56868
rect 158864 56856 158870 56908
rect 158898 56856 158904 56908
rect 158956 56896 158962 56908
rect 162964 56896 162992 57004
rect 170306 56924 170312 56976
rect 170364 56964 170370 56976
rect 170858 56964 170864 56976
rect 170364 56936 170864 56964
rect 170364 56924 170370 56936
rect 170858 56924 170864 56936
rect 170916 56924 170922 56976
rect 217134 56964 217140 56976
rect 171106 56936 217140 56964
rect 158956 56868 162992 56896
rect 158956 56856 158962 56868
rect 163406 56856 163412 56908
rect 163464 56896 163470 56908
rect 171106 56896 171134 56936
rect 217134 56924 217140 56936
rect 217192 56924 217198 56976
rect 217244 56964 217272 57004
rect 217410 56992 217416 57044
rect 217468 57032 217474 57044
rect 218974 57032 218980 57044
rect 217468 57004 218980 57032
rect 217468 56992 217474 57004
rect 218974 56992 218980 57004
rect 219032 56992 219038 57044
rect 218606 56964 218612 56976
rect 217244 56936 218612 56964
rect 218606 56924 218612 56936
rect 218664 56924 218670 56976
rect 218790 56924 218796 56976
rect 218848 56964 218854 56976
rect 258718 56964 258724 56976
rect 218848 56936 258724 56964
rect 218848 56924 218854 56936
rect 258718 56924 258724 56936
rect 258776 56924 258782 56976
rect 163464 56868 171134 56896
rect 163464 56856 163470 56868
rect 174998 56856 175004 56908
rect 175056 56896 175062 56908
rect 180518 56896 180524 56908
rect 175056 56868 180524 56896
rect 175056 56856 175062 56868
rect 180518 56856 180524 56868
rect 180576 56856 180582 56908
rect 180766 56868 200114 56896
rect 127768 56800 128216 56828
rect 127768 56788 127774 56800
rect 133138 56788 133144 56840
rect 133196 56828 133202 56840
rect 133782 56828 133788 56840
rect 133196 56800 133788 56828
rect 133196 56788 133202 56800
rect 133782 56788 133788 56800
rect 133840 56788 133846 56840
rect 134058 56788 134064 56840
rect 134116 56828 134122 56840
rect 135070 56828 135076 56840
rect 134116 56800 135076 56828
rect 134116 56788 134122 56800
rect 135070 56788 135076 56800
rect 135128 56788 135134 56840
rect 138566 56788 138572 56840
rect 138624 56828 138630 56840
rect 143626 56828 143632 56840
rect 138624 56800 143632 56828
rect 138624 56788 138630 56800
rect 143626 56788 143632 56800
rect 143684 56788 143690 56840
rect 145466 56788 145472 56840
rect 145524 56828 145530 56840
rect 145524 56800 150388 56828
rect 145524 56788 145530 56800
rect 125962 56720 125968 56772
rect 126020 56760 126026 56772
rect 126790 56760 126796 56772
rect 126020 56732 126796 56760
rect 126020 56720 126026 56732
rect 126790 56720 126796 56732
rect 126848 56720 126854 56772
rect 141878 56760 141884 56772
rect 129568 56732 141884 56760
rect 129568 56692 129596 56732
rect 141878 56720 141884 56732
rect 141936 56720 141942 56772
rect 145098 56720 145104 56772
rect 145156 56760 145162 56772
rect 147674 56760 147680 56772
rect 145156 56732 147680 56760
rect 145156 56720 145162 56732
rect 147674 56720 147680 56732
rect 147732 56720 147738 56772
rect 149054 56720 149060 56772
rect 149112 56760 149118 56772
rect 150250 56760 150256 56772
rect 149112 56732 150256 56760
rect 149112 56720 149118 56732
rect 150250 56720 150256 56732
rect 150308 56720 150314 56772
rect 150360 56760 150388 56800
rect 150802 56788 150808 56840
rect 150860 56828 150866 56840
rect 151630 56828 151636 56840
rect 150860 56800 151636 56828
rect 150860 56788 150866 56800
rect 151630 56788 151636 56800
rect 151688 56788 151694 56840
rect 177298 56828 177304 56840
rect 151786 56800 177304 56828
rect 151786 56760 151814 56800
rect 177298 56788 177304 56800
rect 177356 56788 177362 56840
rect 180766 56828 180794 56868
rect 179800 56800 180794 56828
rect 150360 56732 151814 56760
rect 154114 56720 154120 56772
rect 154172 56760 154178 56772
rect 157334 56760 157340 56772
rect 154172 56732 157340 56760
rect 154172 56720 154178 56732
rect 157334 56720 157340 56732
rect 157392 56720 157398 56772
rect 157426 56720 157432 56772
rect 157484 56760 157490 56772
rect 157484 56732 158576 56760
rect 157484 56720 157490 56732
rect 158548 56704 158576 56732
rect 171502 56720 171508 56772
rect 171560 56760 171566 56772
rect 179800 56760 179828 56800
rect 180886 56788 180892 56840
rect 180944 56828 180950 56840
rect 181898 56828 181904 56840
rect 180944 56800 181904 56828
rect 180944 56788 180950 56800
rect 181898 56788 181904 56800
rect 181956 56788 181962 56840
rect 184106 56788 184112 56840
rect 184164 56828 184170 56840
rect 184658 56828 184664 56840
rect 184164 56800 184664 56828
rect 184164 56788 184170 56800
rect 184658 56788 184664 56800
rect 184716 56788 184722 56840
rect 184934 56788 184940 56840
rect 184992 56828 184998 56840
rect 186038 56828 186044 56840
rect 184992 56800 186044 56828
rect 184992 56788 184998 56800
rect 186038 56788 186044 56800
rect 186096 56788 186102 56840
rect 189442 56788 189448 56840
rect 189500 56828 189506 56840
rect 190270 56828 190276 56840
rect 189500 56800 190276 56828
rect 189500 56788 189506 56800
rect 190270 56788 190276 56800
rect 190328 56788 190334 56840
rect 191282 56788 191288 56840
rect 191340 56828 191346 56840
rect 191558 56828 191564 56840
rect 191340 56800 191564 56828
rect 191340 56788 191346 56800
rect 191558 56788 191564 56800
rect 191616 56788 191622 56840
rect 192202 56788 192208 56840
rect 192260 56828 192266 56840
rect 192938 56828 192944 56840
rect 192260 56800 192944 56828
rect 192260 56788 192266 56800
rect 192938 56788 192944 56800
rect 192996 56788 193002 56840
rect 193398 56788 193404 56840
rect 193456 56828 193462 56840
rect 194226 56828 194232 56840
rect 193456 56800 194232 56828
rect 193456 56788 193462 56800
rect 194226 56788 194232 56800
rect 194284 56788 194290 56840
rect 196894 56788 196900 56840
rect 196952 56828 196958 56840
rect 197262 56828 197268 56840
rect 196952 56800 197268 56828
rect 196952 56788 196958 56800
rect 197262 56788 197268 56800
rect 197320 56788 197326 56840
rect 197814 56788 197820 56840
rect 197872 56828 197878 56840
rect 198642 56828 198648 56840
rect 197872 56800 198648 56828
rect 197872 56788 197878 56800
rect 198642 56788 198648 56800
rect 198700 56788 198706 56840
rect 199654 56788 199660 56840
rect 199712 56828 199718 56840
rect 199930 56828 199936 56840
rect 199712 56800 199936 56828
rect 199712 56788 199718 56800
rect 199930 56788 199936 56800
rect 199988 56788 199994 56840
rect 200086 56828 200114 56868
rect 200574 56856 200580 56908
rect 200632 56896 200638 56908
rect 201402 56896 201408 56908
rect 200632 56868 201408 56896
rect 200632 56856 200638 56868
rect 201402 56856 201408 56868
rect 201460 56856 201466 56908
rect 202322 56856 202328 56908
rect 202380 56896 202386 56908
rect 202690 56896 202696 56908
rect 202380 56868 202696 56896
rect 202380 56856 202386 56868
rect 202690 56856 202696 56868
rect 202748 56856 202754 56908
rect 203242 56856 203248 56908
rect 203300 56896 203306 56908
rect 203886 56896 203892 56908
rect 203300 56868 203892 56896
rect 203300 56856 203306 56868
rect 203886 56856 203892 56868
rect 203944 56856 203950 56908
rect 204438 56856 204444 56908
rect 204496 56896 204502 56908
rect 205358 56896 205364 56908
rect 204496 56868 205364 56896
rect 204496 56856 204502 56868
rect 205358 56856 205364 56868
rect 205416 56856 205422 56908
rect 205634 56856 205640 56908
rect 205692 56896 205698 56908
rect 206646 56896 206652 56908
rect 205692 56868 206652 56896
rect 205692 56856 205698 56868
rect 206646 56856 206652 56868
rect 206704 56856 206710 56908
rect 207474 56856 207480 56908
rect 207532 56896 207538 56908
rect 208302 56896 208308 56908
rect 207532 56868 208308 56896
rect 207532 56856 207538 56868
rect 208302 56856 208308 56868
rect 208360 56856 208366 56908
rect 210418 56856 210424 56908
rect 210476 56896 210482 56908
rect 229554 56896 229560 56908
rect 210476 56868 229560 56896
rect 210476 56856 210482 56868
rect 229554 56856 229560 56868
rect 229612 56856 229618 56908
rect 200086 56800 202552 56828
rect 171560 56732 179828 56760
rect 171560 56720 171566 56732
rect 179874 56720 179880 56772
rect 179932 56760 179938 56772
rect 180518 56760 180524 56772
rect 179932 56732 180524 56760
rect 179932 56720 179938 56732
rect 180518 56720 180524 56732
rect 180576 56720 180582 56772
rect 180766 56732 200114 56760
rect 125566 56664 129596 56692
rect 129826 56652 129832 56704
rect 129884 56692 129890 56704
rect 130930 56692 130936 56704
rect 129884 56664 130936 56692
rect 129884 56652 129890 56664
rect 130930 56652 130936 56664
rect 130988 56652 130994 56704
rect 131390 56652 131396 56704
rect 131448 56692 131454 56704
rect 132310 56692 132316 56704
rect 131448 56664 132316 56692
rect 131448 56652 131454 56664
rect 132310 56652 132316 56664
rect 132368 56652 132374 56704
rect 132586 56652 132592 56704
rect 132644 56692 132650 56704
rect 133598 56692 133604 56704
rect 132644 56664 133604 56692
rect 132644 56652 132650 56664
rect 133598 56652 133604 56664
rect 133656 56652 133662 56704
rect 134610 56652 134616 56704
rect 134668 56692 134674 56704
rect 135162 56692 135168 56704
rect 134668 56664 135168 56692
rect 134668 56652 134674 56664
rect 135162 56652 135168 56664
rect 135220 56652 135226 56704
rect 135254 56652 135260 56704
rect 135312 56692 135318 56704
rect 136082 56692 136088 56704
rect 135312 56664 136088 56692
rect 135312 56652 135318 56664
rect 136082 56652 136088 56664
rect 136140 56652 136146 56704
rect 136266 56652 136272 56704
rect 136324 56692 136330 56704
rect 141418 56692 141424 56704
rect 136324 56664 137876 56692
rect 136324 56652 136330 56664
rect 109006 56596 115934 56624
rect 115906 56488 115934 56596
rect 120534 56584 120540 56636
rect 120592 56624 120598 56636
rect 121362 56624 121368 56636
rect 120592 56596 121368 56624
rect 120592 56584 120598 56596
rect 121362 56584 121368 56596
rect 121420 56584 121426 56636
rect 121454 56584 121460 56636
rect 121512 56624 121518 56636
rect 122742 56624 122748 56636
rect 121512 56596 122748 56624
rect 121512 56584 121518 56596
rect 122742 56584 122748 56596
rect 122800 56584 122806 56636
rect 122926 56584 122932 56636
rect 122984 56624 122990 56636
rect 123754 56624 123760 56636
rect 122984 56596 123760 56624
rect 122984 56584 122990 56596
rect 123754 56584 123760 56596
rect 123812 56584 123818 56636
rect 124766 56584 124772 56636
rect 124824 56624 124830 56636
rect 125410 56624 125416 56636
rect 124824 56596 125416 56624
rect 124824 56584 124830 56596
rect 125410 56584 125416 56596
rect 125468 56584 125474 56636
rect 125686 56584 125692 56636
rect 125744 56624 125750 56636
rect 126422 56624 126428 56636
rect 125744 56596 126428 56624
rect 125744 56584 125750 56596
rect 126422 56584 126428 56596
rect 126480 56584 126486 56636
rect 127158 56584 127164 56636
rect 127216 56624 127222 56636
rect 127216 56596 127388 56624
rect 127216 56584 127222 56596
rect 117866 56516 117872 56568
rect 117924 56556 117930 56568
rect 127250 56556 127256 56568
rect 117924 56528 127256 56556
rect 117924 56516 117930 56528
rect 127250 56516 127256 56528
rect 127308 56516 127314 56568
rect 122006 56488 122012 56500
rect 115906 56460 122012 56488
rect 122006 56448 122012 56460
rect 122064 56448 122070 56500
rect 127360 56488 127388 56596
rect 127434 56584 127440 56636
rect 127492 56624 127498 56636
rect 127986 56624 127992 56636
rect 127492 56596 127992 56624
rect 127492 56584 127498 56596
rect 127986 56584 127992 56596
rect 128044 56584 128050 56636
rect 128096 56596 128860 56624
rect 127894 56516 127900 56568
rect 127952 56556 127958 56568
rect 128096 56556 128124 56596
rect 127952 56528 128124 56556
rect 128832 56556 128860 56596
rect 128906 56584 128912 56636
rect 128964 56624 128970 56636
rect 129458 56624 129464 56636
rect 128964 56596 129464 56624
rect 128964 56584 128970 56596
rect 129458 56584 129464 56596
rect 129516 56584 129522 56636
rect 130102 56584 130108 56636
rect 130160 56624 130166 56636
rect 130654 56624 130660 56636
rect 130160 56596 130660 56624
rect 130160 56584 130166 56596
rect 130654 56584 130660 56596
rect 130712 56584 130718 56636
rect 131114 56624 131120 56636
rect 130764 56596 131120 56624
rect 130764 56556 130792 56596
rect 131114 56584 131120 56596
rect 131172 56584 131178 56636
rect 131666 56584 131672 56636
rect 131724 56624 131730 56636
rect 132402 56624 132408 56636
rect 131724 56596 132408 56624
rect 131724 56584 131730 56596
rect 132402 56584 132408 56596
rect 132460 56584 132466 56636
rect 132862 56584 132868 56636
rect 132920 56624 132926 56636
rect 133322 56624 133328 56636
rect 132920 56596 133328 56624
rect 132920 56584 132926 56596
rect 133322 56584 133328 56596
rect 133380 56584 133386 56636
rect 134334 56584 134340 56636
rect 134392 56624 134398 56636
rect 134886 56624 134892 56636
rect 134392 56596 134892 56624
rect 134392 56584 134398 56596
rect 134886 56584 134892 56596
rect 134944 56584 134950 56636
rect 135806 56584 135812 56636
rect 135864 56624 135870 56636
rect 136542 56624 136548 56636
rect 135864 56596 136548 56624
rect 135864 56584 135870 56596
rect 136542 56584 136548 56596
rect 136600 56584 136606 56636
rect 137002 56584 137008 56636
rect 137060 56624 137066 56636
rect 137738 56624 137744 56636
rect 137060 56596 137744 56624
rect 137060 56584 137066 56596
rect 137738 56584 137744 56596
rect 137796 56584 137802 56636
rect 137848 56624 137876 56664
rect 137986 56664 141424 56692
rect 137986 56624 138014 56664
rect 141418 56652 141424 56664
rect 141476 56652 141482 56704
rect 146662 56652 146668 56704
rect 146720 56692 146726 56704
rect 147398 56692 147404 56704
rect 146720 56664 147404 56692
rect 146720 56652 146726 56664
rect 147398 56652 147404 56664
rect 147456 56652 147462 56704
rect 149882 56652 149888 56704
rect 149940 56692 149946 56704
rect 150342 56692 150348 56704
rect 149940 56664 150348 56692
rect 149940 56652 149946 56664
rect 150342 56652 150348 56664
rect 150400 56652 150406 56704
rect 150710 56652 150716 56704
rect 150768 56692 150774 56704
rect 151354 56692 151360 56704
rect 150768 56664 151360 56692
rect 150768 56652 150774 56664
rect 151354 56652 151360 56664
rect 151412 56652 151418 56704
rect 157978 56652 157984 56704
rect 158036 56692 158042 56704
rect 158438 56692 158444 56704
rect 158036 56664 158444 56692
rect 158036 56652 158042 56664
rect 158438 56652 158444 56664
rect 158496 56652 158502 56704
rect 158530 56652 158536 56704
rect 158588 56652 158594 56704
rect 160738 56652 160744 56704
rect 160796 56692 160802 56704
rect 161382 56692 161388 56704
rect 160796 56664 161388 56692
rect 160796 56652 160802 56664
rect 161382 56652 161388 56664
rect 161440 56652 161446 56704
rect 164326 56652 164332 56704
rect 164384 56692 164390 56704
rect 165062 56692 165068 56704
rect 164384 56664 165068 56692
rect 164384 56652 164390 56664
rect 165062 56652 165068 56664
rect 165120 56652 165126 56704
rect 165798 56652 165804 56704
rect 165856 56692 165862 56704
rect 166810 56692 166816 56704
rect 165856 56664 166816 56692
rect 165856 56652 165862 56664
rect 166810 56652 166816 56664
rect 166868 56652 166874 56704
rect 137848 56596 138014 56624
rect 138198 56584 138204 56636
rect 138256 56624 138262 56636
rect 139302 56624 139308 56636
rect 138256 56596 139308 56624
rect 138256 56584 138262 56596
rect 139302 56584 139308 56596
rect 139360 56584 139366 56636
rect 139762 56584 139768 56636
rect 139820 56624 139826 56636
rect 140498 56624 140504 56636
rect 139820 56596 140504 56624
rect 139820 56584 139826 56596
rect 140498 56584 140504 56596
rect 140556 56584 140562 56636
rect 141510 56584 141516 56636
rect 141568 56624 141574 56636
rect 142062 56624 142068 56636
rect 141568 56596 142068 56624
rect 141568 56584 141574 56596
rect 142062 56584 142068 56596
rect 142120 56584 142126 56636
rect 142430 56584 142436 56636
rect 142488 56624 142494 56636
rect 143166 56624 143172 56636
rect 142488 56596 143172 56624
rect 142488 56584 142494 56596
rect 143166 56584 143172 56596
rect 143224 56584 143230 56636
rect 144270 56584 144276 56636
rect 144328 56624 144334 56636
rect 144638 56624 144644 56636
rect 144328 56596 144644 56624
rect 144328 56584 144334 56596
rect 144638 56584 144644 56596
rect 144696 56584 144702 56636
rect 145742 56584 145748 56636
rect 145800 56624 145806 56636
rect 146202 56624 146208 56636
rect 145800 56596 146208 56624
rect 145800 56584 145806 56596
rect 146202 56584 146208 56596
rect 146260 56584 146266 56636
rect 147214 56584 147220 56636
rect 147272 56624 147278 56636
rect 147582 56624 147588 56636
rect 147272 56596 147588 56624
rect 147272 56584 147278 56596
rect 147582 56584 147588 56596
rect 147640 56584 147646 56636
rect 149330 56584 149336 56636
rect 149388 56624 149394 56636
rect 150066 56624 150072 56636
rect 149388 56596 150072 56624
rect 149388 56584 149394 56596
rect 150066 56584 150072 56596
rect 150124 56584 150130 56636
rect 151078 56584 151084 56636
rect 151136 56624 151142 56636
rect 151538 56624 151544 56636
rect 151136 56596 151544 56624
rect 151136 56584 151142 56596
rect 151538 56584 151544 56596
rect 151596 56584 151602 56636
rect 157702 56584 157708 56636
rect 157760 56624 157766 56636
rect 158254 56624 158260 56636
rect 157760 56596 158260 56624
rect 157760 56584 157766 56596
rect 158254 56584 158260 56596
rect 158312 56584 158318 56636
rect 158346 56584 158352 56636
rect 158404 56624 158410 56636
rect 158714 56624 158720 56636
rect 158404 56596 158720 56624
rect 158404 56584 158410 56596
rect 158714 56584 158720 56596
rect 158772 56584 158778 56636
rect 159174 56584 159180 56636
rect 159232 56624 159238 56636
rect 159726 56624 159732 56636
rect 159232 56596 159732 56624
rect 159232 56584 159238 56596
rect 159726 56584 159732 56596
rect 159784 56584 159790 56636
rect 160370 56584 160376 56636
rect 160428 56624 160434 56636
rect 160922 56624 160928 56636
rect 160428 56596 160928 56624
rect 160428 56584 160434 56596
rect 160922 56584 160928 56596
rect 160980 56584 160986 56636
rect 161566 56584 161572 56636
rect 161624 56624 161630 56636
rect 162670 56624 162676 56636
rect 161624 56596 162676 56624
rect 161624 56584 161630 56596
rect 162670 56584 162676 56596
rect 162728 56584 162734 56636
rect 163130 56584 163136 56636
rect 163188 56624 163194 56636
rect 163866 56624 163872 56636
rect 163188 56596 163872 56624
rect 163188 56584 163194 56596
rect 163866 56584 163872 56596
rect 163924 56584 163930 56636
rect 164878 56584 164884 56636
rect 164936 56624 164942 56636
rect 165338 56624 165344 56636
rect 164936 56596 165344 56624
rect 164936 56584 164942 56596
rect 165338 56584 165344 56596
rect 165396 56584 165402 56636
rect 166074 56584 166080 56636
rect 166132 56624 166138 56636
rect 166626 56624 166632 56636
rect 166132 56596 166632 56624
rect 166132 56584 166138 56596
rect 166626 56584 166632 56596
rect 166684 56584 166690 56636
rect 173250 56584 173256 56636
rect 173308 56624 173314 56636
rect 180766 56624 180794 56732
rect 181162 56652 181168 56704
rect 181220 56692 181226 56704
rect 182082 56692 182088 56704
rect 181220 56664 182088 56692
rect 181220 56652 181226 56664
rect 182082 56652 182088 56664
rect 182140 56652 182146 56704
rect 182910 56652 182916 56704
rect 182968 56692 182974 56704
rect 183370 56692 183376 56704
rect 182968 56664 183376 56692
rect 182968 56652 182974 56664
rect 183370 56652 183376 56664
rect 183428 56652 183434 56704
rect 183554 56652 183560 56704
rect 183612 56692 183618 56704
rect 190362 56692 190368 56704
rect 183612 56664 190368 56692
rect 183612 56652 183618 56664
rect 190362 56652 190368 56664
rect 190420 56652 190426 56704
rect 196066 56652 196072 56704
rect 196124 56692 196130 56704
rect 197170 56692 197176 56704
rect 196124 56664 197176 56692
rect 196124 56652 196130 56664
rect 197170 56652 197176 56664
rect 197228 56652 197234 56704
rect 198734 56652 198740 56704
rect 198792 56692 198798 56704
rect 199654 56692 199660 56704
rect 198792 56664 199660 56692
rect 198792 56652 198798 56664
rect 199654 56652 199660 56664
rect 199712 56652 199718 56704
rect 173308 56596 180794 56624
rect 173308 56584 173314 56596
rect 180978 56584 180984 56636
rect 181036 56624 181042 56636
rect 187602 56624 187608 56636
rect 181036 56596 187608 56624
rect 181036 56584 181042 56596
rect 187602 56584 187608 56596
rect 187660 56584 187666 56636
rect 200086 56624 200114 56732
rect 201494 56652 201500 56704
rect 201552 56692 201558 56704
rect 202414 56692 202420 56704
rect 201552 56664 202420 56692
rect 201552 56652 201558 56664
rect 202414 56652 202420 56664
rect 202472 56652 202478 56704
rect 202524 56692 202552 56800
rect 203150 56788 203156 56840
rect 203208 56828 203214 56840
rect 203794 56828 203800 56840
rect 203208 56800 203800 56828
rect 203208 56788 203214 56800
rect 203794 56788 203800 56800
rect 203852 56788 203858 56840
rect 205910 56788 205916 56840
rect 205968 56828 205974 56840
rect 206922 56828 206928 56840
rect 205968 56800 206928 56828
rect 205968 56788 205974 56800
rect 206922 56788 206928 56800
rect 206980 56788 206986 56840
rect 208118 56788 208124 56840
rect 208176 56828 208182 56840
rect 233878 56828 233884 56840
rect 208176 56800 233884 56828
rect 208176 56788 208182 56800
rect 233878 56788 233884 56800
rect 233936 56788 233942 56840
rect 271138 56760 271144 56772
rect 209746 56732 271144 56760
rect 209038 56692 209044 56704
rect 202524 56664 209044 56692
rect 209038 56652 209044 56664
rect 209096 56652 209102 56704
rect 209746 56624 209774 56732
rect 271138 56720 271144 56732
rect 271196 56720 271202 56772
rect 214006 56652 214012 56704
rect 214064 56692 214070 56704
rect 228266 56692 228272 56704
rect 214064 56664 228272 56692
rect 214064 56652 214070 56664
rect 228266 56652 228272 56664
rect 228324 56652 228330 56704
rect 200086 56596 209774 56624
rect 213454 56584 213460 56636
rect 213512 56624 213518 56636
rect 225782 56624 225788 56636
rect 213512 56596 225788 56624
rect 213512 56584 213518 56596
rect 225782 56584 225788 56596
rect 225840 56584 225846 56636
rect 128832 56528 130792 56556
rect 127952 56516 127958 56528
rect 163682 56516 163688 56568
rect 163740 56556 163746 56568
rect 407758 56556 407764 56568
rect 163740 56528 407764 56556
rect 163740 56516 163746 56528
rect 407758 56516 407764 56528
rect 407816 56516 407822 56568
rect 128170 56488 128176 56500
rect 127360 56460 128176 56488
rect 128170 56448 128176 56460
rect 128228 56448 128234 56500
rect 167270 56448 167276 56500
rect 167328 56488 167334 56500
rect 421558 56488 421564 56500
rect 167328 56460 421564 56488
rect 167328 56448 167334 56460
rect 421558 56448 421564 56460
rect 421616 56448 421622 56500
rect 183462 56380 183468 56432
rect 183520 56420 183526 56432
rect 443638 56420 443644 56432
rect 183520 56392 443644 56420
rect 183520 56380 183526 56392
rect 443638 56380 443644 56392
rect 443696 56380 443702 56432
rect 185302 56312 185308 56364
rect 185360 56352 185366 56364
rect 450538 56352 450544 56364
rect 185360 56324 450544 56352
rect 185360 56312 185366 56324
rect 450538 56312 450544 56324
rect 450596 56312 450602 56364
rect 184382 56244 184388 56296
rect 184440 56284 184446 56296
rect 447778 56284 447784 56296
rect 184440 56256 447784 56284
rect 184440 56244 184446 56256
rect 447778 56244 447784 56256
rect 447836 56244 447842 56296
rect 186222 56176 186228 56228
rect 186280 56216 186286 56228
rect 454678 56216 454684 56228
rect 186280 56188 454684 56216
rect 186280 56176 186286 56188
rect 454678 56176 454684 56188
rect 454736 56176 454742 56228
rect 187970 56108 187976 56160
rect 188028 56148 188034 56160
rect 461578 56148 461584 56160
rect 188028 56120 461584 56148
rect 188028 56108 188034 56120
rect 461578 56108 461584 56120
rect 461636 56108 461642 56160
rect 189166 56040 189172 56092
rect 189224 56080 189230 56092
rect 472618 56080 472624 56092
rect 189224 56052 472624 56080
rect 189224 56040 189230 56052
rect 472618 56040 472624 56052
rect 472676 56040 472682 56092
rect 187050 55972 187056 56024
rect 187108 56012 187114 56024
rect 500954 56012 500960 56024
rect 187108 55984 500960 56012
rect 187108 55972 187114 55984
rect 500954 55972 500960 55984
rect 501012 55972 501018 56024
rect 188982 55904 188988 55956
rect 189040 55944 189046 55956
rect 507854 55944 507860 55956
rect 189040 55916 507860 55944
rect 189040 55904 189046 55916
rect 507854 55904 507860 55916
rect 507912 55904 507918 55956
rect 202966 55836 202972 55888
rect 203024 55876 203030 55888
rect 564434 55876 564440 55888
rect 203024 55848 564440 55876
rect 203024 55836 203030 55848
rect 564434 55836 564440 55848
rect 564492 55836 564498 55888
rect 139394 55768 139400 55820
rect 139452 55808 139458 55820
rect 313274 55808 313280 55820
rect 139452 55780 313280 55808
rect 139452 55768 139458 55780
rect 313274 55768 313280 55780
rect 313332 55768 313338 55820
rect 118786 55700 118792 55752
rect 118844 55740 118850 55752
rect 231854 55740 231860 55752
rect 118844 55712 231860 55740
rect 118844 55700 118850 55712
rect 231854 55700 231860 55712
rect 231912 55700 231918 55752
rect 116026 55632 116032 55684
rect 116084 55672 116090 55684
rect 220814 55672 220820 55684
rect 116084 55644 220820 55672
rect 116084 55632 116090 55644
rect 220814 55632 220820 55644
rect 220872 55632 220878 55684
rect 115198 55564 115204 55616
rect 115256 55604 115262 55616
rect 218054 55604 218060 55616
rect 115256 55576 218060 55604
rect 115256 55564 115262 55576
rect 218054 55564 218060 55576
rect 218112 55564 218118 55616
rect 218606 55564 218612 55616
rect 218664 55604 218670 55616
rect 219066 55604 219072 55616
rect 218664 55576 219072 55604
rect 218664 55564 218670 55576
rect 219066 55564 219072 55576
rect 219124 55564 219130 55616
rect 112438 55496 112444 55548
rect 112496 55536 112502 55548
rect 113082 55536 113088 55548
rect 112496 55508 113088 55536
rect 112496 55496 112502 55508
rect 113082 55496 113088 55508
rect 113140 55496 113146 55548
rect 127250 55496 127256 55548
rect 127308 55536 127314 55548
rect 227714 55536 227720 55548
rect 127308 55508 227720 55536
rect 127308 55496 127314 55508
rect 227714 55496 227720 55508
rect 227772 55496 227778 55548
rect 103790 55428 103796 55480
rect 103848 55468 103854 55480
rect 104710 55468 104716 55480
rect 103848 55440 104716 55468
rect 103848 55428 103854 55440
rect 104710 55428 104716 55440
rect 104768 55428 104774 55480
rect 119338 55428 119344 55480
rect 119396 55468 119402 55480
rect 119890 55468 119896 55480
rect 119396 55440 119896 55468
rect 119396 55428 119402 55440
rect 119890 55428 119896 55440
rect 119948 55428 119954 55480
rect 130746 55428 130752 55480
rect 130804 55468 130810 55480
rect 131022 55468 131028 55480
rect 130804 55440 131028 55468
rect 130804 55428 130810 55440
rect 131022 55428 131028 55440
rect 131080 55428 131086 55480
rect 146386 55428 146392 55480
rect 146444 55468 146450 55480
rect 213914 55468 213920 55480
rect 146444 55440 213920 55468
rect 146444 55428 146450 55440
rect 213914 55428 213920 55440
rect 213972 55428 213978 55480
rect 143534 55360 143540 55412
rect 143592 55400 143598 55412
rect 209774 55400 209780 55412
rect 143592 55372 209780 55400
rect 143592 55360 143598 55372
rect 209774 55360 209780 55372
rect 209832 55360 209838 55412
rect 100754 55292 100760 55344
rect 100812 55332 100818 55344
rect 102042 55332 102048 55344
rect 100812 55304 102048 55332
rect 100812 55292 100818 55304
rect 102042 55292 102048 55304
rect 102100 55292 102106 55344
rect 130470 55292 130476 55344
rect 130528 55332 130534 55344
rect 131022 55332 131028 55344
rect 130528 55304 131028 55332
rect 130528 55292 130534 55304
rect 131022 55292 131028 55304
rect 131080 55292 131086 55344
rect 142154 55156 142160 55208
rect 142212 55196 142218 55208
rect 324314 55196 324320 55208
rect 142212 55168 324320 55196
rect 142212 55156 142218 55168
rect 324314 55156 324320 55168
rect 324372 55156 324378 55208
rect 143074 55088 143080 55140
rect 143132 55128 143138 55140
rect 327074 55128 327080 55140
rect 143132 55100 327080 55128
rect 143132 55088 143138 55100
rect 327074 55088 327080 55100
rect 327132 55088 327138 55140
rect 143902 55020 143908 55072
rect 143960 55060 143966 55072
rect 331214 55060 331220 55072
rect 143960 55032 331220 55060
rect 143960 55020 143966 55032
rect 331214 55020 331220 55032
rect 331272 55020 331278 55072
rect 162762 54952 162768 55004
rect 162820 54992 162826 55004
rect 405734 54992 405740 55004
rect 162820 54964 405740 54992
rect 162820 54952 162826 54964
rect 405734 54952 405740 54964
rect 405792 54952 405798 55004
rect 164602 54884 164608 54936
rect 164660 54924 164666 54936
rect 412634 54924 412640 54936
rect 164660 54896 412640 54924
rect 164660 54884 164666 54896
rect 412634 54884 412640 54896
rect 412692 54884 412698 54936
rect 53650 54816 53656 54868
rect 53708 54856 53714 54868
rect 73246 54856 73252 54868
rect 53708 54828 73252 54856
rect 53708 54816 53714 54828
rect 73246 54816 73252 54828
rect 73304 54816 73310 54868
rect 165522 54816 165528 54868
rect 165580 54856 165586 54868
rect 414658 54856 414664 54868
rect 165580 54828 414664 54856
rect 165580 54816 165586 54828
rect 414658 54816 414664 54828
rect 414716 54816 414722 54868
rect 49602 54748 49608 54800
rect 49660 54788 49666 54800
rect 72326 54788 72332 54800
rect 49660 54760 72332 54788
rect 49660 54748 49666 54760
rect 72326 54748 72332 54760
rect 72384 54748 72390 54800
rect 166442 54748 166448 54800
rect 166500 54788 166506 54800
rect 417418 54788 417424 54800
rect 166500 54760 417424 54788
rect 166500 54748 166506 54760
rect 417418 54748 417424 54760
rect 417476 54748 417482 54800
rect 45462 54680 45468 54732
rect 45520 54720 45526 54732
rect 71406 54720 71412 54732
rect 45520 54692 71412 54720
rect 45520 54680 45526 54692
rect 71406 54680 71412 54692
rect 71464 54680 71470 54732
rect 167178 54680 167184 54732
rect 167236 54720 167242 54732
rect 425790 54720 425796 54732
rect 167236 54692 425796 54720
rect 167236 54680 167242 54692
rect 425790 54680 425796 54692
rect 425848 54680 425854 54732
rect 45370 54612 45376 54664
rect 45428 54652 45434 54664
rect 71130 54652 71136 54664
rect 45428 54624 71136 54652
rect 45428 54612 45434 54624
rect 71130 54612 71136 54624
rect 71188 54612 71194 54664
rect 161014 54612 161020 54664
rect 161072 54652 161078 54664
rect 161290 54652 161296 54664
rect 161072 54624 161296 54652
rect 161072 54612 161078 54624
rect 161290 54612 161296 54624
rect 161348 54612 161354 54664
rect 172054 54612 172060 54664
rect 172112 54652 172118 54664
rect 439498 54652 439504 54664
rect 172112 54624 439504 54652
rect 172112 54612 172118 54624
rect 439498 54612 439504 54624
rect 439556 54612 439562 54664
rect 44082 54544 44088 54596
rect 44140 54584 44146 54596
rect 70854 54584 70860 54596
rect 44140 54556 70860 54584
rect 44140 54544 44146 54556
rect 70854 54544 70860 54556
rect 70912 54544 70918 54596
rect 189074 54544 189080 54596
rect 189132 54584 189138 54596
rect 475378 54584 475384 54596
rect 189132 54556 475384 54584
rect 189132 54544 189138 54556
rect 475378 54544 475384 54556
rect 475436 54544 475442 54596
rect 37182 54476 37188 54528
rect 37240 54516 37246 54528
rect 69290 54516 69296 54528
rect 37240 54488 69296 54516
rect 37240 54476 37246 54488
rect 69290 54476 69296 54488
rect 69348 54476 69354 54528
rect 136082 54476 136088 54528
rect 136140 54516 136146 54528
rect 136450 54516 136456 54528
rect 136140 54488 136456 54516
rect 136140 54476 136146 54488
rect 136450 54476 136456 54488
rect 136508 54476 136514 54528
rect 160094 54476 160100 54528
rect 160152 54516 160158 54528
rect 161290 54516 161296 54528
rect 160152 54488 161296 54516
rect 160152 54476 160158 54488
rect 161290 54476 161296 54488
rect 161348 54476 161354 54528
rect 203150 54476 203156 54528
rect 203208 54516 203214 54528
rect 544378 54516 544384 54528
rect 203208 54488 544384 54516
rect 203208 54476 203214 54488
rect 544378 54476 544384 54488
rect 544436 54476 544442 54528
rect 141234 54408 141240 54460
rect 141292 54448 141298 54460
rect 320174 54448 320180 54460
rect 141292 54420 320180 54448
rect 141292 54408 141298 54420
rect 320174 54408 320180 54420
rect 320232 54408 320238 54460
rect 140314 54340 140320 54392
rect 140372 54380 140378 54392
rect 316034 54380 316040 54392
rect 140372 54352 316040 54380
rect 140372 54340 140378 54352
rect 316034 54340 316040 54352
rect 316092 54340 316098 54392
rect 143626 54272 143632 54324
rect 143684 54312 143690 54324
rect 309134 54312 309140 54324
rect 143684 54284 309140 54312
rect 143684 54272 143690 54284
rect 309134 54272 309140 54284
rect 309192 54272 309198 54324
rect 136726 54204 136732 54256
rect 136784 54244 136790 54256
rect 302234 54244 302240 54256
rect 136784 54216 302240 54244
rect 136784 54204 136790 54216
rect 302234 54204 302240 54216
rect 302292 54204 302298 54256
rect 153194 53728 153200 53780
rect 153252 53768 153258 53780
rect 367094 53768 367100 53780
rect 153252 53740 367100 53768
rect 153252 53728 153258 53740
rect 367094 53728 367100 53740
rect 367152 53728 367158 53780
rect 169110 53660 169116 53712
rect 169168 53700 169174 53712
rect 430574 53700 430580 53712
rect 169168 53672 430580 53700
rect 169168 53660 169174 53672
rect 430574 53660 430580 53672
rect 430632 53660 430638 53712
rect 170030 53592 170036 53644
rect 170088 53632 170094 53644
rect 432598 53632 432604 53644
rect 170088 53604 432604 53632
rect 170088 53592 170094 53604
rect 432598 53592 432604 53604
rect 432656 53592 432662 53644
rect 136174 53524 136180 53576
rect 136232 53564 136238 53576
rect 136358 53564 136364 53576
rect 136232 53536 136364 53564
rect 136232 53524 136238 53536
rect 136358 53524 136364 53536
rect 136416 53524 136422 53576
rect 188246 53524 188252 53576
rect 188304 53564 188310 53576
rect 468478 53564 468484 53576
rect 188304 53536 468484 53564
rect 188304 53524 188310 53536
rect 468478 53524 468484 53536
rect 468536 53524 468542 53576
rect 175642 53456 175648 53508
rect 175700 53496 175706 53508
rect 456794 53496 456800 53508
rect 175700 53468 456800 53496
rect 175700 53456 175706 53468
rect 456794 53456 456800 53468
rect 456852 53456 456858 53508
rect 128630 53388 128636 53440
rect 128688 53428 128694 53440
rect 129550 53428 129556 53440
rect 128688 53400 129556 53428
rect 128688 53388 128694 53400
rect 129550 53388 129556 53400
rect 129608 53388 129614 53440
rect 191006 53388 191012 53440
rect 191064 53428 191070 53440
rect 479518 53428 479524 53440
rect 191064 53400 479524 53428
rect 191064 53388 191070 53400
rect 479518 53388 479524 53400
rect 479576 53388 479582 53440
rect 192018 53320 192024 53372
rect 192076 53360 192082 53372
rect 483658 53360 483664 53372
rect 192076 53332 483664 53360
rect 192076 53320 192082 53332
rect 483658 53320 483664 53332
rect 483716 53320 483722 53372
rect 193674 53252 193680 53304
rect 193732 53292 193738 53304
rect 512638 53292 512644 53304
rect 193732 53264 512644 53292
rect 193732 53252 193738 53264
rect 512638 53252 512644 53264
rect 512696 53252 512702 53304
rect 194594 53184 194600 53236
rect 194652 53224 194658 53236
rect 519538 53224 519544 53236
rect 194652 53196 519544 53224
rect 194652 53184 194658 53196
rect 519538 53184 519544 53196
rect 519596 53184 519602 53236
rect 191834 53116 191840 53168
rect 191892 53156 191898 53168
rect 520274 53156 520280 53168
rect 191892 53128 520280 53156
rect 191892 53116 191898 53128
rect 520274 53116 520280 53128
rect 520332 53116 520338 53168
rect 195422 53048 195428 53100
rect 195480 53088 195486 53100
rect 526438 53088 526444 53100
rect 195480 53060 526444 53088
rect 195480 53048 195486 53060
rect 526438 53048 526444 53060
rect 526496 53048 526502 53100
rect 125318 52980 125324 53032
rect 125376 53020 125382 53032
rect 258074 53020 258080 53032
rect 125376 52992 258080 53020
rect 125376 52980 125382 52992
rect 258074 52980 258080 52992
rect 258132 52980 258138 53032
rect 124490 52912 124496 52964
rect 124548 52952 124554 52964
rect 253934 52952 253940 52964
rect 124548 52924 253940 52952
rect 124548 52912 124554 52924
rect 253934 52912 253940 52924
rect 253992 52912 253998 52964
rect 119062 52844 119068 52896
rect 119120 52884 119126 52896
rect 233234 52884 233240 52896
rect 119120 52856 233240 52884
rect 119120 52844 119126 52856
rect 233234 52844 233240 52856
rect 233292 52844 233298 52896
rect 141878 52776 141884 52828
rect 141936 52816 141942 52828
rect 251174 52816 251180 52828
rect 141936 52788 251180 52816
rect 141936 52776 141942 52788
rect 251174 52776 251180 52788
rect 251232 52776 251238 52828
rect 136634 52708 136640 52760
rect 136692 52748 136698 52760
rect 240134 52748 240140 52760
rect 136692 52720 240140 52748
rect 136692 52708 136698 52720
rect 240134 52708 240140 52720
rect 240192 52708 240198 52760
rect 147674 52368 147680 52420
rect 147732 52408 147738 52420
rect 335354 52408 335360 52420
rect 147732 52380 335360 52408
rect 147732 52368 147738 52380
rect 335354 52368 335360 52380
rect 335412 52368 335418 52420
rect 146018 52300 146024 52352
rect 146076 52340 146082 52352
rect 339494 52340 339500 52352
rect 146076 52312 339500 52340
rect 146076 52300 146082 52312
rect 339494 52300 339500 52312
rect 339552 52300 339558 52352
rect 146938 52232 146944 52284
rect 146996 52272 147002 52284
rect 342254 52272 342260 52284
rect 146996 52244 342260 52272
rect 146996 52232 147002 52244
rect 342254 52232 342260 52244
rect 342312 52232 342318 52284
rect 147858 52164 147864 52216
rect 147916 52204 147922 52216
rect 346394 52204 346400 52216
rect 147916 52176 346400 52204
rect 147916 52164 147922 52176
rect 346394 52164 346400 52176
rect 346452 52164 346458 52216
rect 150434 52096 150440 52148
rect 150492 52136 150498 52148
rect 357434 52136 357440 52148
rect 150492 52108 357440 52136
rect 150492 52096 150498 52108
rect 357434 52096 357440 52108
rect 357492 52096 357498 52148
rect 150526 52028 150532 52080
rect 150584 52068 150590 52080
rect 360194 52068 360200 52080
rect 150584 52040 360200 52068
rect 150584 52028 150590 52040
rect 360194 52028 360200 52040
rect 360252 52028 360258 52080
rect 152274 51960 152280 52012
rect 152332 52000 152338 52012
rect 364334 52000 364340 52012
rect 152332 51972 364340 52000
rect 152332 51960 152338 51972
rect 364334 51960 364340 51972
rect 364392 51960 364398 52012
rect 172974 51892 172980 51944
rect 173032 51932 173038 51944
rect 445754 51932 445760 51944
rect 173032 51904 445760 51932
rect 173032 51892 173038 51904
rect 445754 51892 445760 51904
rect 445812 51892 445818 51944
rect 108022 51824 108028 51876
rect 108080 51864 108086 51876
rect 108850 51864 108856 51876
rect 108080 51836 108856 51864
rect 108080 51824 108086 51836
rect 108850 51824 108856 51836
rect 108908 51824 108914 51876
rect 173894 51824 173900 51876
rect 173952 51864 173958 51876
rect 448514 51864 448520 51876
rect 173952 51836 448520 51864
rect 173952 51824 173958 51836
rect 448514 51824 448520 51836
rect 448572 51824 448578 51876
rect 175550 51756 175556 51808
rect 175608 51796 175614 51808
rect 459554 51796 459560 51808
rect 175608 51768 459560 51796
rect 175608 51756 175614 51768
rect 459554 51756 459560 51768
rect 459612 51756 459618 51808
rect 199378 51688 199384 51740
rect 199436 51728 199442 51740
rect 530578 51728 530584 51740
rect 199436 51700 530584 51728
rect 199436 51688 199442 51700
rect 530578 51688 530584 51700
rect 530636 51688 530642 51740
rect 146110 51008 146116 51060
rect 146168 51048 146174 51060
rect 311894 51048 311900 51060
rect 146168 51020 311900 51048
rect 146168 51008 146174 51020
rect 311894 51008 311900 51020
rect 311952 51008 311958 51060
rect 174814 50940 174820 50992
rect 174872 50980 174878 50992
rect 452654 50980 452660 50992
rect 174872 50952 452660 50980
rect 174872 50940 174878 50952
rect 452654 50940 452660 50952
rect 452712 50940 452718 50992
rect 177482 50872 177488 50924
rect 177540 50912 177546 50924
rect 463694 50912 463700 50924
rect 177540 50884 463700 50912
rect 177540 50872 177546 50884
rect 463694 50872 463700 50884
rect 463752 50872 463758 50924
rect 178402 50804 178408 50856
rect 178460 50844 178466 50856
rect 466454 50844 466460 50856
rect 178460 50816 466460 50844
rect 178460 50804 178466 50816
rect 466454 50804 466460 50816
rect 466512 50804 466518 50856
rect 178034 50736 178040 50788
rect 178092 50776 178098 50788
rect 470594 50776 470600 50788
rect 178092 50748 470600 50776
rect 178092 50736 178098 50748
rect 470594 50736 470600 50748
rect 470652 50736 470658 50788
rect 200206 50668 200212 50720
rect 200264 50708 200270 50720
rect 533338 50708 533344 50720
rect 200264 50680 533344 50708
rect 200264 50668 200270 50680
rect 533338 50668 533344 50680
rect 533396 50668 533402 50720
rect 201126 50600 201132 50652
rect 201184 50640 201190 50652
rect 537478 50640 537484 50652
rect 201184 50612 537484 50640
rect 201184 50600 201190 50612
rect 537478 50600 537484 50612
rect 537536 50600 537542 50652
rect 197538 50532 197544 50584
rect 197596 50572 197602 50584
rect 542354 50572 542360 50584
rect 197596 50544 542360 50572
rect 197596 50532 197602 50544
rect 542354 50532 542360 50544
rect 542412 50532 542418 50584
rect 204714 50464 204720 50516
rect 204772 50504 204778 50516
rect 551278 50504 551284 50516
rect 204772 50476 551284 50504
rect 204772 50464 204778 50476
rect 551278 50464 551284 50476
rect 551336 50464 551342 50516
rect 197630 50396 197636 50448
rect 197688 50436 197694 50448
rect 546494 50436 546500 50448
rect 197688 50408 546500 50436
rect 197688 50396 197694 50408
rect 546494 50396 546500 50408
rect 546552 50396 546558 50448
rect 123294 50328 123300 50380
rect 123352 50368 123358 50380
rect 124122 50368 124128 50380
rect 123352 50340 124128 50368
rect 123352 50328 123358 50340
rect 124122 50328 124128 50340
rect 124180 50328 124186 50380
rect 202046 50328 202052 50380
rect 202104 50368 202110 50380
rect 560294 50368 560300 50380
rect 202104 50340 560300 50368
rect 202104 50328 202110 50340
rect 560294 50328 560300 50340
rect 560352 50328 560358 50380
rect 139486 50260 139492 50312
rect 139544 50300 139550 50312
rect 291194 50300 291200 50312
rect 139544 50272 291200 50300
rect 139544 50260 139550 50272
rect 291194 50260 291200 50272
rect 291252 50260 291258 50312
rect 158714 49104 158720 49156
rect 158772 49144 158778 49156
rect 316126 49144 316132 49156
rect 158772 49116 316132 49144
rect 158772 49104 158778 49116
rect 316126 49104 316132 49116
rect 316184 49104 316190 49156
rect 165706 49036 165712 49088
rect 165764 49076 165770 49088
rect 329834 49076 329840 49088
rect 165764 49048 329840 49076
rect 165764 49036 165770 49048
rect 329834 49036 329840 49048
rect 329892 49036 329898 49088
rect 155126 48968 155132 49020
rect 155184 49008 155190 49020
rect 340874 49008 340880 49020
rect 155184 48980 340880 49008
rect 155184 48968 155190 48980
rect 340874 48968 340880 48980
rect 340932 48968 340938 49020
rect 55766 46180 55772 46232
rect 55824 46220 55830 46232
rect 580350 46220 580356 46232
rect 55824 46192 580356 46220
rect 55824 46180 55830 46192
rect 580350 46180 580356 46192
rect 580408 46180 580414 46232
rect 3326 45500 3332 45552
rect 3384 45540 3390 45552
rect 21358 45540 21364 45552
rect 3384 45512 21364 45540
rect 3384 45500 3390 45512
rect 21358 45500 21364 45512
rect 21416 45500 21422 45552
rect 238110 33056 238116 33108
rect 238168 33096 238174 33108
rect 580166 33096 580172 33108
rect 238168 33068 580172 33096
rect 238168 33056 238174 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 2774 32852 2780 32904
rect 2832 32892 2838 32904
rect 4798 32892 4804 32904
rect 2832 32864 4804 32892
rect 2832 32852 2838 32864
rect 4798 32852 4804 32864
rect 4856 32852 4862 32904
rect 234062 20612 234068 20664
rect 234120 20652 234126 20664
rect 580074 20652 580080 20664
rect 234120 20624 580080 20652
rect 234120 20612 234126 20624
rect 580074 20612 580080 20624
rect 580132 20612 580138 20664
rect 159358 19932 159364 19984
rect 159416 19972 159422 19984
rect 347774 19972 347780 19984
rect 159416 19944 347780 19972
rect 159416 19932 159422 19944
rect 347774 19932 347780 19944
rect 347832 19932 347838 19984
rect 119798 18640 119804 18692
rect 119856 18680 119862 18692
rect 235994 18680 236000 18692
rect 119856 18652 236000 18680
rect 119856 18640 119862 18652
rect 235994 18640 236000 18652
rect 236052 18640 236058 18692
rect 209038 18572 209044 18624
rect 209096 18612 209102 18624
rect 440234 18612 440240 18624
rect 209096 18584 440240 18612
rect 209096 18572 209102 18584
rect 440234 18572 440240 18584
rect 440292 18572 440298 18624
rect 146938 17892 146944 17944
rect 146996 17932 147002 17944
rect 260834 17932 260840 17944
rect 146996 17904 260840 17932
rect 146996 17892 147002 17904
rect 260834 17892 260840 17904
rect 260892 17892 260898 17944
rect 129366 17824 129372 17876
rect 129424 17864 129430 17876
rect 269114 17864 269120 17876
rect 129424 17836 269120 17864
rect 129424 17824 129430 17836
rect 269114 17824 269120 17836
rect 269172 17824 269178 17876
rect 129274 17756 129280 17808
rect 129332 17796 129338 17808
rect 273254 17796 273260 17808
rect 129332 17768 273260 17796
rect 129332 17756 129338 17768
rect 273254 17756 273260 17768
rect 273312 17756 273318 17808
rect 130654 17688 130660 17740
rect 130712 17728 130718 17740
rect 276014 17728 276020 17740
rect 130712 17700 276020 17728
rect 130712 17688 130718 17700
rect 276014 17688 276020 17700
rect 276072 17688 276078 17740
rect 130746 17620 130752 17672
rect 130804 17660 130810 17672
rect 280154 17660 280160 17672
rect 130804 17632 280160 17660
rect 130804 17620 130810 17632
rect 280154 17620 280160 17632
rect 280212 17620 280218 17672
rect 132126 17552 132132 17604
rect 132184 17592 132190 17604
rect 284294 17592 284300 17604
rect 132184 17564 284300 17592
rect 132184 17552 132190 17564
rect 284294 17552 284300 17564
rect 284352 17552 284358 17604
rect 133506 17484 133512 17536
rect 133564 17524 133570 17536
rect 287054 17524 287060 17536
rect 133564 17496 287060 17524
rect 133564 17484 133570 17496
rect 287054 17484 287060 17496
rect 287112 17484 287118 17536
rect 177298 17416 177304 17468
rect 177356 17456 177362 17468
rect 336734 17456 336740 17468
rect 177356 17428 336740 17456
rect 177356 17416 177362 17428
rect 336734 17416 336740 17428
rect 336792 17416 336798 17468
rect 162118 17348 162124 17400
rect 162176 17388 162182 17400
rect 325694 17388 325700 17400
rect 162176 17360 325700 17388
rect 162176 17348 162182 17360
rect 325694 17348 325700 17360
rect 325752 17348 325758 17400
rect 136266 17280 136272 17332
rect 136324 17320 136330 17332
rect 300854 17320 300860 17332
rect 136324 17292 300860 17320
rect 136324 17280 136330 17292
rect 300854 17280 300860 17292
rect 300912 17280 300918 17332
rect 148318 17212 148324 17264
rect 148376 17252 148382 17264
rect 318794 17252 318800 17264
rect 148376 17224 318800 17252
rect 148376 17212 148382 17224
rect 318794 17212 318800 17224
rect 318852 17212 318858 17264
rect 137278 17144 137284 17196
rect 137336 17184 137342 17196
rect 247034 17184 247040 17196
rect 137336 17156 247040 17184
rect 137336 17144 137342 17156
rect 247034 17144 247040 17156
rect 247092 17144 247098 17196
rect 116946 17076 116952 17128
rect 117004 17116 117010 17128
rect 224954 17116 224960 17128
rect 117004 17088 224960 17116
rect 117004 17076 117010 17088
rect 224954 17076 224960 17088
rect 225012 17076 225018 17128
rect 144178 17008 144184 17060
rect 144236 17048 144242 17060
rect 242894 17048 242900 17060
rect 144236 17020 242900 17048
rect 144236 17008 144242 17020
rect 242894 17008 242900 17020
rect 242952 17008 242958 17060
rect 121270 16532 121276 16584
rect 121328 16572 121334 16584
rect 238110 16572 238116 16584
rect 121328 16544 238116 16572
rect 121328 16532 121334 16544
rect 238110 16532 238116 16544
rect 238168 16532 238174 16584
rect 121178 16464 121184 16516
rect 121236 16504 121242 16516
rect 241698 16504 241704 16516
rect 121236 16476 241704 16504
rect 121236 16464 121242 16476
rect 241698 16464 241704 16476
rect 241756 16464 241762 16516
rect 122558 16396 122564 16448
rect 122616 16436 122622 16448
rect 245194 16436 245200 16448
rect 122616 16408 245200 16436
rect 122616 16396 122622 16408
rect 245194 16396 245200 16408
rect 245252 16396 245258 16448
rect 123846 16328 123852 16380
rect 123904 16368 123910 16380
rect 248782 16368 248788 16380
rect 123904 16340 248788 16368
rect 123904 16328 123910 16340
rect 248782 16328 248788 16340
rect 248840 16328 248846 16380
rect 123938 16260 123944 16312
rect 123996 16300 124002 16312
rect 252370 16300 252376 16312
rect 123996 16272 252376 16300
rect 123996 16260 124002 16272
rect 252370 16260 252376 16272
rect 252428 16260 252434 16312
rect 125410 16192 125416 16244
rect 125468 16232 125474 16244
rect 255866 16232 255872 16244
rect 125468 16204 255872 16232
rect 125468 16192 125474 16204
rect 255866 16192 255872 16204
rect 255924 16192 255930 16244
rect 126606 16124 126612 16176
rect 126664 16164 126670 16176
rect 259454 16164 259460 16176
rect 126664 16136 259460 16164
rect 126664 16124 126670 16136
rect 259454 16124 259460 16136
rect 259512 16124 259518 16176
rect 126698 16056 126704 16108
rect 126756 16096 126762 16108
rect 262950 16096 262956 16108
rect 126756 16068 262956 16096
rect 126756 16056 126762 16068
rect 262950 16056 262956 16068
rect 263008 16056 263014 16108
rect 127986 15988 127992 16040
rect 128044 16028 128050 16040
rect 266538 16028 266544 16040
rect 128044 16000 266544 16028
rect 128044 15988 128050 16000
rect 266538 15988 266544 16000
rect 266596 15988 266602 16040
rect 206646 15920 206652 15972
rect 206704 15960 206710 15972
rect 575106 15960 575112 15972
rect 206704 15932 575112 15960
rect 206704 15920 206710 15932
rect 575106 15920 575112 15932
rect 575164 15920 575170 15972
rect 206738 15852 206744 15904
rect 206796 15892 206802 15904
rect 578602 15892 578608 15904
rect 206796 15864 578608 15892
rect 206796 15852 206802 15864
rect 578602 15852 578608 15864
rect 578660 15852 578666 15904
rect 119890 15784 119896 15836
rect 119948 15824 119954 15836
rect 234614 15824 234620 15836
rect 119948 15796 234620 15824
rect 119948 15784 119954 15796
rect 234614 15784 234620 15796
rect 234672 15784 234678 15836
rect 118418 15716 118424 15768
rect 118476 15756 118482 15768
rect 231026 15756 231032 15768
rect 118476 15728 231032 15756
rect 118476 15716 118482 15728
rect 231026 15716 231032 15728
rect 231084 15716 231090 15768
rect 118510 15648 118516 15700
rect 118568 15688 118574 15700
rect 227530 15688 227536 15700
rect 118568 15660 227536 15688
rect 118568 15648 118574 15660
rect 227530 15648 227536 15660
rect 227588 15648 227594 15700
rect 117038 15580 117044 15632
rect 117096 15620 117102 15632
rect 223942 15620 223948 15632
rect 117096 15592 223948 15620
rect 117096 15580 117102 15592
rect 223942 15580 223948 15592
rect 224000 15580 224006 15632
rect 115658 15512 115664 15564
rect 115716 15552 115722 15564
rect 220446 15552 220452 15564
rect 115716 15524 220452 15552
rect 115716 15512 115722 15524
rect 220446 15512 220452 15524
rect 220504 15512 220510 15564
rect 115566 15444 115572 15496
rect 115624 15484 115630 15496
rect 216858 15484 216864 15496
rect 115624 15456 216864 15484
rect 115624 15444 115630 15456
rect 216858 15444 216864 15456
rect 216916 15444 216922 15496
rect 114370 15376 114376 15428
rect 114428 15416 114434 15428
rect 213362 15416 213368 15428
rect 114428 15388 213368 15416
rect 114428 15376 114434 15388
rect 213362 15376 213368 15388
rect 213420 15376 213426 15428
rect 112714 15308 112720 15360
rect 112772 15348 112778 15360
rect 209866 15348 209872 15360
rect 112772 15320 209872 15348
rect 112772 15308 112778 15320
rect 209866 15308 209872 15320
rect 209924 15308 209930 15360
rect 188890 15104 188896 15156
rect 188948 15144 188954 15156
rect 504174 15144 504180 15156
rect 188948 15116 504180 15144
rect 188948 15104 188954 15116
rect 504174 15104 504180 15116
rect 504232 15104 504238 15156
rect 188706 15036 188712 15088
rect 188764 15076 188770 15088
rect 507670 15076 507676 15088
rect 188764 15048 507676 15076
rect 188764 15036 188770 15048
rect 507670 15036 507676 15048
rect 507728 15036 507734 15088
rect 190270 14968 190276 15020
rect 190328 15008 190334 15020
rect 511258 15008 511264 15020
rect 190328 14980 511264 15008
rect 190328 14968 190334 14980
rect 511258 14968 511264 14980
rect 511316 14968 511322 15020
rect 190178 14900 190184 14952
rect 190236 14940 190242 14952
rect 514754 14940 514760 14952
rect 190236 14912 514760 14940
rect 190236 14900 190242 14912
rect 514754 14900 514760 14912
rect 514812 14900 514818 14952
rect 191558 14832 191564 14884
rect 191616 14872 191622 14884
rect 518342 14872 518348 14884
rect 191616 14844 518348 14872
rect 191616 14832 191622 14844
rect 518342 14832 518348 14844
rect 518400 14832 518406 14884
rect 192938 14764 192944 14816
rect 192996 14804 193002 14816
rect 521838 14804 521844 14816
rect 192996 14776 521844 14804
rect 192996 14764 193002 14776
rect 521838 14764 521844 14776
rect 521896 14764 521902 14816
rect 193030 14696 193036 14748
rect 193088 14736 193094 14748
rect 525426 14736 525432 14748
rect 193088 14708 525432 14736
rect 193088 14696 193094 14708
rect 525426 14696 525432 14708
rect 525484 14696 525490 14748
rect 194318 14628 194324 14680
rect 194376 14668 194382 14680
rect 529014 14668 529020 14680
rect 194376 14640 529020 14668
rect 194376 14628 194382 14640
rect 529014 14628 529020 14640
rect 529072 14628 529078 14680
rect 195698 14560 195704 14612
rect 195756 14600 195762 14612
rect 532510 14600 532516 14612
rect 195756 14572 532516 14600
rect 195756 14560 195762 14572
rect 532510 14560 532516 14572
rect 532568 14560 532574 14612
rect 195790 14492 195796 14544
rect 195848 14532 195854 14544
rect 536098 14532 536104 14544
rect 195848 14504 536104 14532
rect 195848 14492 195854 14504
rect 536098 14492 536104 14504
rect 536156 14492 536162 14544
rect 141510 14424 141516 14476
rect 141568 14464 141574 14476
rect 182542 14464 182548 14476
rect 141568 14436 182548 14464
rect 141568 14424 141574 14436
rect 182542 14424 182548 14436
rect 182600 14424 182606 14476
rect 196894 14424 196900 14476
rect 196952 14464 196958 14476
rect 539594 14464 539600 14476
rect 196952 14436 539600 14464
rect 196952 14424 196958 14436
rect 539594 14424 539600 14436
rect 539652 14424 539658 14476
rect 187418 14356 187424 14408
rect 187476 14396 187482 14408
rect 500586 14396 500592 14408
rect 187476 14368 500592 14396
rect 187476 14356 187482 14368
rect 500586 14356 500592 14368
rect 500644 14356 500650 14408
rect 186130 14288 186136 14340
rect 186188 14328 186194 14340
rect 497090 14328 497096 14340
rect 186188 14300 497096 14328
rect 186188 14288 186194 14300
rect 497090 14288 497096 14300
rect 497148 14288 497154 14340
rect 186038 14220 186044 14272
rect 186096 14260 186102 14272
rect 493502 14260 493508 14272
rect 186096 14232 493508 14260
rect 186096 14220 186102 14232
rect 493502 14220 493508 14232
rect 493560 14220 493566 14272
rect 184658 14152 184664 14204
rect 184716 14192 184722 14204
rect 489914 14192 489920 14204
rect 184716 14164 489920 14192
rect 184716 14152 184722 14164
rect 489914 14152 489920 14164
rect 489972 14152 489978 14204
rect 183186 14084 183192 14136
rect 183244 14124 183250 14136
rect 486418 14124 486424 14136
rect 183244 14096 486424 14124
rect 183244 14084 183250 14096
rect 486418 14084 486424 14096
rect 486476 14084 486482 14136
rect 183278 14016 183284 14068
rect 183336 14056 183342 14068
rect 481634 14056 481640 14068
rect 183336 14028 481640 14056
rect 183336 14016 183342 14028
rect 481634 14016 481640 14028
rect 481692 14016 481698 14068
rect 181714 13948 181720 14000
rect 181772 13988 181778 14000
rect 478138 13988 478144 14000
rect 181772 13960 478144 13988
rect 181772 13948 181778 13960
rect 478138 13948 478144 13960
rect 478196 13948 478202 14000
rect 180518 13880 180524 13932
rect 180576 13920 180582 13932
rect 473354 13920 473360 13932
rect 180576 13892 473360 13920
rect 180576 13880 180582 13892
rect 473354 13880 473360 13892
rect 473412 13880 473418 13932
rect 162486 13744 162492 13796
rect 162544 13784 162550 13796
rect 403618 13784 403624 13796
rect 162544 13756 403624 13784
rect 162544 13744 162550 13756
rect 403618 13744 403624 13756
rect 403676 13744 403682 13796
rect 163958 13676 163964 13728
rect 164016 13716 164022 13728
rect 407206 13716 407212 13728
rect 164016 13688 407212 13716
rect 164016 13676 164022 13688
rect 407206 13676 407212 13688
rect 407264 13676 407270 13728
rect 164050 13608 164056 13660
rect 164108 13648 164114 13660
rect 410794 13648 410800 13660
rect 164108 13620 410800 13648
rect 164108 13608 164114 13620
rect 410794 13608 410800 13620
rect 410852 13608 410858 13660
rect 165338 13540 165344 13592
rect 165396 13580 165402 13592
rect 414290 13580 414296 13592
rect 165396 13552 414296 13580
rect 165396 13540 165402 13552
rect 414290 13540 414296 13552
rect 414348 13540 414354 13592
rect 166810 13472 166816 13524
rect 166868 13512 166874 13524
rect 417418 13512 417424 13524
rect 166868 13484 417424 13512
rect 166868 13472 166874 13484
rect 417418 13472 417424 13484
rect 417476 13472 417482 13524
rect 166718 13404 166724 13456
rect 166776 13444 166782 13456
rect 421374 13444 421380 13456
rect 166776 13416 421380 13444
rect 166776 13404 166782 13416
rect 421374 13404 421380 13416
rect 421432 13404 421438 13456
rect 168098 13336 168104 13388
rect 168156 13376 168162 13388
rect 423766 13376 423772 13388
rect 168156 13348 423772 13376
rect 168156 13336 168162 13348
rect 423766 13336 423772 13348
rect 423824 13336 423830 13388
rect 169478 13268 169484 13320
rect 169536 13308 169542 13320
rect 428458 13308 428464 13320
rect 169536 13280 428464 13308
rect 169536 13268 169542 13280
rect 428458 13268 428464 13280
rect 428516 13268 428522 13320
rect 169386 13200 169392 13252
rect 169444 13240 169450 13252
rect 432046 13240 432052 13252
rect 169444 13212 432052 13240
rect 169444 13200 169450 13212
rect 432046 13200 432052 13212
rect 432104 13200 432110 13252
rect 170858 13132 170864 13184
rect 170916 13172 170922 13184
rect 435542 13172 435548 13184
rect 170916 13144 435548 13172
rect 170916 13132 170922 13144
rect 435542 13132 435548 13144
rect 435600 13132 435606 13184
rect 172238 13064 172244 13116
rect 172296 13104 172302 13116
rect 439130 13104 439136 13116
rect 172296 13076 439136 13104
rect 172296 13064 172302 13076
rect 439130 13064 439136 13076
rect 439188 13064 439194 13116
rect 161014 12996 161020 13048
rect 161072 13036 161078 13048
rect 398834 13036 398840 13048
rect 161072 13008 398840 13036
rect 161072 12996 161078 13008
rect 398834 12996 398840 13008
rect 398892 12996 398898 13048
rect 161106 12928 161112 12980
rect 161164 12968 161170 12980
rect 396534 12968 396540 12980
rect 161164 12940 396540 12968
rect 161164 12928 161170 12940
rect 396534 12928 396540 12940
rect 396592 12928 396598 12980
rect 159818 12860 159824 12912
rect 159876 12900 159882 12912
rect 393038 12900 393044 12912
rect 159876 12872 393044 12900
rect 159876 12860 159882 12872
rect 393038 12860 393044 12872
rect 393096 12860 393102 12912
rect 158346 12792 158352 12844
rect 158404 12832 158410 12844
rect 389450 12832 389456 12844
rect 158404 12804 389456 12832
rect 158404 12792 158410 12804
rect 389450 12792 389456 12804
rect 389508 12792 389514 12844
rect 158254 12724 158260 12776
rect 158312 12764 158318 12776
rect 385954 12764 385960 12776
rect 158312 12736 385960 12764
rect 158312 12724 158318 12736
rect 385954 12724 385960 12736
rect 386012 12724 386018 12776
rect 156966 12656 156972 12708
rect 157024 12696 157030 12708
rect 382366 12696 382372 12708
rect 157024 12668 382372 12696
rect 157024 12656 157030 12668
rect 382366 12656 382372 12668
rect 382424 12656 382430 12708
rect 156874 12588 156880 12640
rect 156932 12628 156938 12640
rect 378870 12628 378876 12640
rect 156932 12600 378876 12628
rect 156932 12588 156938 12600
rect 378870 12588 378876 12600
rect 378928 12588 378934 12640
rect 155678 12520 155684 12572
rect 155736 12560 155742 12572
rect 373994 12560 374000 12572
rect 155736 12532 374000 12560
rect 155736 12520 155742 12532
rect 373994 12520 374000 12532
rect 374052 12520 374058 12572
rect 137738 12384 137744 12436
rect 137796 12424 137802 12436
rect 304350 12424 304356 12436
rect 137796 12396 304356 12424
rect 137796 12384 137802 12396
rect 304350 12384 304356 12396
rect 304408 12384 304414 12436
rect 137830 12316 137836 12368
rect 137888 12356 137894 12368
rect 307938 12356 307944 12368
rect 137888 12328 307944 12356
rect 137888 12316 137894 12328
rect 307938 12316 307944 12328
rect 307996 12316 308002 12368
rect 139210 12248 139216 12300
rect 139268 12288 139274 12300
rect 311434 12288 311440 12300
rect 139268 12260 311440 12288
rect 139268 12248 139274 12260
rect 311434 12248 311440 12260
rect 311492 12248 311498 12300
rect 140498 12180 140504 12232
rect 140556 12220 140562 12232
rect 315022 12220 315028 12232
rect 140556 12192 315028 12220
rect 140556 12180 140562 12192
rect 315022 12180 315028 12192
rect 315080 12180 315086 12232
rect 140590 12112 140596 12164
rect 140648 12152 140654 12164
rect 318518 12152 318524 12164
rect 140648 12124 318524 12152
rect 140648 12112 140654 12124
rect 318518 12112 318524 12124
rect 318576 12112 318582 12164
rect 142062 12044 142068 12096
rect 142120 12084 142126 12096
rect 322106 12084 322112 12096
rect 142120 12056 322112 12084
rect 142120 12044 142126 12056
rect 322106 12044 322112 12056
rect 322164 12044 322170 12096
rect 143166 11976 143172 12028
rect 143224 12016 143230 12028
rect 325602 12016 325608 12028
rect 143224 11988 325608 12016
rect 143224 11976 143230 11988
rect 325602 11976 325608 11988
rect 325660 11976 325666 12028
rect 143350 11908 143356 11960
rect 143408 11948 143414 11960
rect 329190 11948 329196 11960
rect 143408 11920 329196 11948
rect 143408 11908 143414 11920
rect 329190 11908 329196 11920
rect 329248 11908 329254 11960
rect 144638 11840 144644 11892
rect 144696 11880 144702 11892
rect 332686 11880 332692 11892
rect 144696 11852 332692 11880
rect 144696 11840 144702 11852
rect 332686 11840 332692 11852
rect 332744 11840 332750 11892
rect 175090 11772 175096 11824
rect 175148 11812 175154 11824
rect 450446 11812 450452 11824
rect 175148 11784 450452 11812
rect 175148 11772 175154 11784
rect 450446 11772 450452 11784
rect 450504 11772 450510 11824
rect 177850 11704 177856 11756
rect 177908 11744 177914 11756
rect 465166 11744 465172 11756
rect 177908 11716 465172 11744
rect 177908 11704 177914 11716
rect 465166 11704 465172 11716
rect 465224 11704 465230 11756
rect 136358 11636 136364 11688
rect 136416 11676 136422 11688
rect 299474 11676 299480 11688
rect 136416 11648 299480 11676
rect 136416 11636 136422 11648
rect 299474 11636 299480 11648
rect 299532 11636 299538 11688
rect 136450 11568 136456 11620
rect 136508 11608 136514 11620
rect 297266 11608 297272 11620
rect 136508 11580 297272 11608
rect 136508 11568 136514 11580
rect 297266 11568 297272 11580
rect 297324 11568 297330 11620
rect 134886 11500 134892 11552
rect 134944 11540 134950 11552
rect 293678 11540 293684 11552
rect 134944 11512 293684 11540
rect 134944 11500 134950 11512
rect 293678 11500 293684 11512
rect 293736 11500 293742 11552
rect 133690 11432 133696 11484
rect 133748 11472 133754 11484
rect 290182 11472 290188 11484
rect 133748 11444 290188 11472
rect 133748 11432 133754 11444
rect 290182 11432 290188 11444
rect 290240 11432 290246 11484
rect 133598 11364 133604 11416
rect 133656 11404 133662 11416
rect 286594 11404 286600 11416
rect 133656 11376 286600 11404
rect 133656 11364 133662 11376
rect 286594 11364 286600 11376
rect 286652 11364 286658 11416
rect 130838 11296 130844 11348
rect 130896 11336 130902 11348
rect 279510 11336 279516 11348
rect 130896 11308 279516 11336
rect 130896 11296 130902 11308
rect 279510 11296 279516 11308
rect 279568 11296 279574 11348
rect 130930 11228 130936 11280
rect 130988 11268 130994 11280
rect 276106 11268 276112 11280
rect 130988 11240 276112 11268
rect 130988 11228 130994 11240
rect 276106 11228 276112 11240
rect 276164 11228 276170 11280
rect 128078 11160 128084 11212
rect 128136 11200 128142 11212
rect 268838 11200 268844 11212
rect 128136 11172 268844 11200
rect 128136 11160 128142 11172
rect 268838 11160 268844 11172
rect 268896 11160 268902 11212
rect 128170 11092 128176 11144
rect 128228 11132 128234 11144
rect 265342 11132 265348 11144
rect 128228 11104 265348 11132
rect 128228 11092 128234 11104
rect 265342 11092 265348 11104
rect 265400 11092 265406 11144
rect 209774 11024 209780 11076
rect 209832 11064 209838 11076
rect 210970 11064 210976 11076
rect 209832 11036 210976 11064
rect 209832 11024 209838 11036
rect 210970 11024 210976 11036
rect 211028 11024 211034 11076
rect 197078 10956 197084 11008
rect 197136 10996 197142 11008
rect 541986 10996 541992 11008
rect 197136 10968 541992 10996
rect 197136 10956 197142 10968
rect 541986 10956 541992 10968
rect 542044 10956 542050 11008
rect 108666 10888 108672 10940
rect 108724 10928 108730 10940
rect 188522 10928 188528 10940
rect 108724 10900 188528 10928
rect 108724 10888 108730 10900
rect 188522 10888 188528 10900
rect 188580 10888 188586 10940
rect 198550 10888 198556 10940
rect 198608 10928 198614 10940
rect 545482 10928 545488 10940
rect 198608 10900 545488 10928
rect 198608 10888 198614 10900
rect 545482 10888 545488 10900
rect 545540 10888 545546 10940
rect 108574 10820 108580 10872
rect 108632 10860 108638 10872
rect 190822 10860 190828 10872
rect 108632 10832 190828 10860
rect 108632 10820 108638 10832
rect 190822 10820 190828 10832
rect 190880 10820 190886 10872
rect 199746 10820 199752 10872
rect 199804 10860 199810 10872
rect 547874 10860 547880 10872
rect 199804 10832 547880 10860
rect 199804 10820 199810 10832
rect 547874 10820 547880 10832
rect 547932 10820 547938 10872
rect 108758 10752 108764 10804
rect 108816 10792 108822 10804
rect 192018 10792 192024 10804
rect 108816 10764 192024 10792
rect 108816 10752 108822 10764
rect 192018 10752 192024 10764
rect 192076 10752 192082 10804
rect 199838 10752 199844 10804
rect 199896 10792 199902 10804
rect 552658 10792 552664 10804
rect 199896 10764 552664 10792
rect 199896 10752 199902 10764
rect 552658 10752 552664 10764
rect 552716 10752 552722 10804
rect 110046 10684 110052 10736
rect 110104 10724 110110 10736
rect 193214 10724 193220 10736
rect 110104 10696 193220 10724
rect 110104 10684 110110 10696
rect 193214 10684 193220 10696
rect 193272 10684 193278 10736
rect 201310 10684 201316 10736
rect 201368 10724 201374 10736
rect 556154 10724 556160 10736
rect 201368 10696 556160 10724
rect 201368 10684 201374 10696
rect 556154 10684 556160 10696
rect 556212 10684 556218 10736
rect 110230 10616 110236 10668
rect 110288 10656 110294 10668
rect 195422 10656 195428 10668
rect 110288 10628 195428 10656
rect 110288 10616 110294 10628
rect 195422 10616 195428 10628
rect 195480 10616 195486 10668
rect 202506 10616 202512 10668
rect 202564 10656 202570 10668
rect 559742 10656 559748 10668
rect 202564 10628 559748 10656
rect 202564 10616 202570 10628
rect 559742 10616 559748 10628
rect 559800 10616 559806 10668
rect 110138 10548 110144 10600
rect 110196 10588 110202 10600
rect 197906 10588 197912 10600
rect 110196 10560 197912 10588
rect 110196 10548 110202 10560
rect 197906 10548 197912 10560
rect 197964 10548 197970 10600
rect 202598 10548 202604 10600
rect 202656 10588 202662 10600
rect 563238 10588 563244 10600
rect 202656 10560 563244 10588
rect 202656 10548 202662 10560
rect 563238 10548 563244 10560
rect 563296 10548 563302 10600
rect 111426 10480 111432 10532
rect 111484 10520 111490 10532
rect 199102 10520 199108 10532
rect 111484 10492 199108 10520
rect 111484 10480 111490 10492
rect 199102 10480 199108 10492
rect 199160 10480 199166 10532
rect 203978 10480 203984 10532
rect 204036 10520 204042 10532
rect 566826 10520 566832 10532
rect 204036 10492 566832 10520
rect 204036 10480 204042 10492
rect 566826 10480 566832 10492
rect 566884 10480 566890 10532
rect 111518 10412 111524 10464
rect 111576 10452 111582 10464
rect 201586 10452 201592 10464
rect 111576 10424 201592 10452
rect 111576 10412 111582 10424
rect 201586 10412 201592 10424
rect 201644 10412 201650 10464
rect 205358 10412 205364 10464
rect 205416 10452 205422 10464
rect 570322 10452 570328 10464
rect 205416 10424 570328 10452
rect 205416 10412 205422 10424
rect 570322 10412 570328 10424
rect 570380 10412 570386 10464
rect 111334 10344 111340 10396
rect 111392 10384 111398 10396
rect 201494 10384 201500 10396
rect 111392 10356 201500 10384
rect 111392 10344 111398 10356
rect 201494 10344 201500 10356
rect 201552 10344 201558 10396
rect 205450 10344 205456 10396
rect 205508 10384 205514 10396
rect 572714 10384 572720 10396
rect 205508 10356 572720 10384
rect 205508 10344 205514 10356
rect 572714 10344 572720 10356
rect 572772 10344 572778 10396
rect 112898 10276 112904 10328
rect 112956 10316 112962 10328
rect 205082 10316 205088 10328
rect 112956 10288 205088 10316
rect 112956 10276 112962 10288
rect 205082 10276 205088 10288
rect 205140 10276 205146 10328
rect 206830 10276 206836 10328
rect 206888 10316 206894 10328
rect 577406 10316 577412 10328
rect 206888 10288 577412 10316
rect 206888 10276 206894 10288
rect 577406 10276 577412 10288
rect 577464 10276 577470 10328
rect 196986 10208 196992 10260
rect 197044 10248 197050 10260
rect 538398 10248 538404 10260
rect 197044 10220 538404 10248
rect 197044 10208 197050 10220
rect 538398 10208 538404 10220
rect 538456 10208 538462 10260
rect 118602 10140 118608 10192
rect 118660 10180 118666 10192
rect 229830 10180 229836 10192
rect 118660 10152 229836 10180
rect 118660 10140 118666 10152
rect 229830 10140 229836 10152
rect 229888 10140 229894 10192
rect 117130 10072 117136 10124
rect 117188 10112 117194 10124
rect 226426 10112 226432 10124
rect 117188 10084 226432 10112
rect 117188 10072 117194 10084
rect 226426 10072 226432 10084
rect 226484 10072 226490 10124
rect 116854 10004 116860 10056
rect 116912 10044 116918 10056
rect 222746 10044 222752 10056
rect 116912 10016 222752 10044
rect 116912 10004 116918 10016
rect 222746 10004 222752 10016
rect 222804 10004 222810 10056
rect 115750 9936 115756 9988
rect 115808 9976 115814 9988
rect 218606 9976 218612 9988
rect 115808 9948 218612 9976
rect 115808 9936 115814 9948
rect 218606 9936 218612 9948
rect 218664 9936 218670 9988
rect 115474 9868 115480 9920
rect 115532 9908 115538 9920
rect 215662 9908 215668 9920
rect 115532 9880 215668 9908
rect 115532 9868 115538 9880
rect 215662 9868 215668 9880
rect 215720 9868 215726 9920
rect 114462 9800 114468 9852
rect 114520 9840 114526 9852
rect 212166 9840 212172 9852
rect 114520 9812 212172 9840
rect 114520 9800 114526 9812
rect 212166 9800 212172 9812
rect 212224 9800 212230 9852
rect 112806 9732 112812 9784
rect 112864 9772 112870 9784
rect 208578 9772 208584 9784
rect 112864 9744 208584 9772
rect 112864 9732 112870 9744
rect 208578 9732 208584 9744
rect 208636 9732 208642 9784
rect 173710 9596 173716 9648
rect 173768 9636 173774 9648
rect 448606 9636 448612 9648
rect 173768 9608 448612 9636
rect 173768 9596 173774 9608
rect 448606 9596 448612 9608
rect 448664 9596 448670 9648
rect 175182 9528 175188 9580
rect 175240 9568 175246 9580
rect 452102 9568 452108 9580
rect 175240 9540 452108 9568
rect 175240 9528 175246 9540
rect 452102 9528 452108 9540
rect 452160 9528 452166 9580
rect 176470 9460 176476 9512
rect 176528 9500 176534 9512
rect 455690 9500 455696 9512
rect 176528 9472 455696 9500
rect 176528 9460 176534 9472
rect 455690 9460 455696 9472
rect 455748 9460 455754 9512
rect 101674 9392 101680 9444
rect 101732 9432 101738 9444
rect 163682 9432 163688 9444
rect 101732 9404 163688 9432
rect 101732 9392 101738 9404
rect 163682 9392 163688 9404
rect 163740 9392 163746 9444
rect 176378 9392 176384 9444
rect 176436 9432 176442 9444
rect 459186 9432 459192 9444
rect 176436 9404 459192 9432
rect 176436 9392 176442 9404
rect 459186 9392 459192 9404
rect 459244 9392 459250 9444
rect 103238 9324 103244 9376
rect 103296 9364 103302 9376
rect 167178 9364 167184 9376
rect 103296 9336 167184 9364
rect 103296 9324 103302 9336
rect 167178 9324 167184 9336
rect 167236 9324 167242 9376
rect 177942 9324 177948 9376
rect 178000 9364 178006 9376
rect 462774 9364 462780 9376
rect 178000 9336 462780 9364
rect 178000 9324 178006 9336
rect 462774 9324 462780 9336
rect 462832 9324 462838 9376
rect 103330 9256 103336 9308
rect 103388 9296 103394 9308
rect 170674 9296 170680 9308
rect 103388 9268 170680 9296
rect 103388 9256 103394 9268
rect 170674 9256 170680 9268
rect 170732 9256 170738 9308
rect 179230 9256 179236 9308
rect 179288 9296 179294 9308
rect 466270 9296 466276 9308
rect 179288 9268 466276 9296
rect 179288 9256 179294 9268
rect 466270 9256 466276 9268
rect 466328 9256 466334 9308
rect 104526 9188 104532 9240
rect 104584 9228 104590 9240
rect 174262 9228 174268 9240
rect 104584 9200 174268 9228
rect 104584 9188 104590 9200
rect 174262 9188 174268 9200
rect 174320 9188 174326 9240
rect 179322 9188 179328 9240
rect 179380 9228 179386 9240
rect 469858 9228 469864 9240
rect 179380 9200 469864 9228
rect 179380 9188 179386 9200
rect 469858 9188 469864 9200
rect 469916 9188 469922 9240
rect 105906 9120 105912 9172
rect 105964 9160 105970 9172
rect 177850 9160 177856 9172
rect 105964 9132 177856 9160
rect 105964 9120 105970 9132
rect 177850 9120 177856 9132
rect 177908 9120 177914 9172
rect 180610 9120 180616 9172
rect 180668 9160 180674 9172
rect 473446 9160 473452 9172
rect 180668 9132 473452 9160
rect 180668 9120 180674 9132
rect 473446 9120 473452 9132
rect 473504 9120 473510 9172
rect 105998 9052 106004 9104
rect 106056 9092 106062 9104
rect 181438 9092 181444 9104
rect 106056 9064 181444 9092
rect 106056 9052 106062 9064
rect 181438 9052 181444 9064
rect 181496 9052 181502 9104
rect 181898 9052 181904 9104
rect 181956 9092 181962 9104
rect 476942 9092 476948 9104
rect 181956 9064 476948 9092
rect 181956 9052 181962 9064
rect 476942 9052 476948 9064
rect 477000 9052 477006 9104
rect 107470 8984 107476 9036
rect 107528 9024 107534 9036
rect 184934 9024 184940 9036
rect 107528 8996 184940 9024
rect 107528 8984 107534 8996
rect 184934 8984 184940 8996
rect 184992 8984 184998 9036
rect 185946 8984 185952 9036
rect 186004 9024 186010 9036
rect 495894 9024 495900 9036
rect 186004 8996 495900 9024
rect 186004 8984 186010 8996
rect 495894 8984 495900 8996
rect 495952 8984 495958 9036
rect 107378 8916 107384 8968
rect 107436 8956 107442 8968
rect 187326 8956 187332 8968
rect 107436 8928 187332 8956
rect 107436 8916 107442 8928
rect 187326 8916 187332 8928
rect 187384 8916 187390 8968
rect 187510 8916 187516 8968
rect 187568 8956 187574 8968
rect 499390 8956 499396 8968
rect 187568 8928 499396 8956
rect 187568 8916 187574 8928
rect 499390 8916 499396 8928
rect 499448 8916 499454 8968
rect 172330 8848 172336 8900
rect 172388 8888 172394 8900
rect 443822 8888 443828 8900
rect 172388 8860 443828 8888
rect 172388 8848 172394 8860
rect 443822 8848 443828 8860
rect 443880 8848 443886 8900
rect 173802 8780 173808 8832
rect 173860 8820 173866 8832
rect 445018 8820 445024 8832
rect 173860 8792 445024 8820
rect 173860 8780 173866 8792
rect 445018 8780 445024 8792
rect 445076 8780 445082 8832
rect 172146 8712 172152 8764
rect 172204 8752 172210 8764
rect 441522 8752 441528 8764
rect 172204 8724 441528 8752
rect 172204 8712 172210 8724
rect 441522 8712 441528 8724
rect 441580 8712 441586 8764
rect 170950 8644 170956 8696
rect 171008 8684 171014 8696
rect 437934 8684 437940 8696
rect 171008 8656 437940 8684
rect 171008 8644 171014 8656
rect 437934 8644 437940 8656
rect 437992 8644 437998 8696
rect 168190 8576 168196 8628
rect 168248 8616 168254 8628
rect 422570 8616 422576 8628
rect 168248 8588 422576 8616
rect 168248 8576 168254 8588
rect 422570 8576 422576 8588
rect 422628 8576 422634 8628
rect 166626 8508 166632 8560
rect 166684 8548 166690 8560
rect 418982 8548 418988 8560
rect 166684 8520 418988 8548
rect 166684 8508 166690 8520
rect 418982 8508 418988 8520
rect 419040 8508 419046 8560
rect 97258 8440 97264 8492
rect 97316 8480 97322 8492
rect 103698 8480 103704 8492
rect 97316 8452 103704 8480
rect 97316 8440 97322 8452
rect 103698 8440 103704 8452
rect 103756 8440 103762 8492
rect 162578 8440 162584 8492
rect 162636 8480 162642 8492
rect 404814 8480 404820 8492
rect 162636 8452 404820 8480
rect 162636 8440 162642 8452
rect 404814 8440 404820 8452
rect 404872 8440 404878 8492
rect 162670 8372 162676 8424
rect 162728 8412 162734 8424
rect 401318 8412 401324 8424
rect 162728 8384 401324 8412
rect 162728 8372 162734 8384
rect 401318 8372 401324 8384
rect 401376 8372 401382 8424
rect 158438 8304 158444 8356
rect 158496 8344 158502 8356
rect 387150 8344 387156 8356
rect 158496 8316 387156 8344
rect 158496 8304 158502 8316
rect 387150 8304 387156 8316
rect 387208 8304 387214 8356
rect 152918 8236 152924 8288
rect 152976 8276 152982 8288
rect 367002 8276 367008 8288
rect 152976 8248 367008 8276
rect 152976 8236 152982 8248
rect 367002 8236 367008 8248
rect 367060 8236 367066 8288
rect 154298 8168 154304 8220
rect 154356 8208 154362 8220
rect 370590 8208 370596 8220
rect 154356 8180 370596 8208
rect 154356 8168 154362 8180
rect 370590 8168 370596 8180
rect 370648 8168 370654 8220
rect 155862 8100 155868 8152
rect 155920 8140 155926 8152
rect 374086 8140 374092 8152
rect 155920 8112 374092 8140
rect 155920 8100 155926 8112
rect 374086 8100 374092 8112
rect 374144 8100 374150 8152
rect 155770 8032 155776 8084
rect 155828 8072 155834 8084
rect 377674 8072 377680 8084
rect 155828 8044 377680 8072
rect 155828 8032 155834 8044
rect 377674 8032 377680 8044
rect 377732 8032 377738 8084
rect 157058 7964 157064 8016
rect 157116 8004 157122 8016
rect 381170 8004 381176 8016
rect 157116 7976 381176 8004
rect 157116 7964 157122 7976
rect 381170 7964 381176 7976
rect 381228 7964 381234 8016
rect 94958 7896 94964 7948
rect 95016 7936 95022 7948
rect 137646 7936 137652 7948
rect 95016 7908 137652 7936
rect 95016 7896 95022 7908
rect 137646 7896 137652 7908
rect 137704 7896 137710 7948
rect 158530 7896 158536 7948
rect 158588 7936 158594 7948
rect 384758 7936 384764 7948
rect 158588 7908 384764 7936
rect 158588 7896 158594 7908
rect 384758 7896 384764 7908
rect 384816 7896 384822 7948
rect 96338 7828 96344 7880
rect 96396 7868 96402 7880
rect 141234 7868 141240 7880
rect 96396 7840 141240 7868
rect 96396 7828 96402 7840
rect 141234 7828 141240 7840
rect 141292 7828 141298 7880
rect 158622 7828 158628 7880
rect 158680 7868 158686 7880
rect 388254 7868 388260 7880
rect 158680 7840 388260 7868
rect 158680 7828 158686 7840
rect 388254 7828 388260 7840
rect 388312 7828 388318 7880
rect 97626 7760 97632 7812
rect 97684 7800 97690 7812
rect 144730 7800 144736 7812
rect 97684 7772 144736 7800
rect 97684 7760 97690 7772
rect 144730 7760 144736 7772
rect 144788 7760 144794 7812
rect 159910 7760 159916 7812
rect 159968 7800 159974 7812
rect 391842 7800 391848 7812
rect 159968 7772 391848 7800
rect 159968 7760 159974 7772
rect 391842 7760 391848 7772
rect 391900 7760 391906 7812
rect 99006 7692 99012 7744
rect 99064 7732 99070 7744
rect 151814 7732 151820 7744
rect 99064 7704 151820 7732
rect 99064 7692 99070 7704
rect 151814 7692 151820 7704
rect 151872 7692 151878 7744
rect 161290 7692 161296 7744
rect 161348 7732 161354 7744
rect 395338 7732 395344 7744
rect 161348 7704 395344 7732
rect 161348 7692 161354 7704
rect 395338 7692 395344 7704
rect 395396 7692 395402 7744
rect 86310 7624 86316 7676
rect 86368 7664 86374 7676
rect 97442 7664 97448 7676
rect 86368 7636 97448 7664
rect 86368 7624 86374 7636
rect 97442 7624 97448 7636
rect 97500 7624 97506 7676
rect 98914 7624 98920 7676
rect 98972 7664 98978 7676
rect 155402 7664 155408 7676
rect 98972 7636 155408 7664
rect 98972 7624 98978 7636
rect 155402 7624 155408 7636
rect 155460 7624 155466 7676
rect 161198 7624 161204 7676
rect 161256 7664 161262 7676
rect 398926 7664 398932 7676
rect 161256 7636 398932 7664
rect 161256 7624 161262 7636
rect 398926 7624 398932 7636
rect 398984 7624 398990 7676
rect 85482 7556 85488 7608
rect 85540 7596 85546 7608
rect 98822 7596 98828 7608
rect 85540 7568 98828 7596
rect 85540 7556 85546 7568
rect 98822 7556 98828 7568
rect 98880 7556 98886 7608
rect 100386 7556 100392 7608
rect 100444 7596 100450 7608
rect 158898 7596 158904 7608
rect 100444 7568 158904 7596
rect 100444 7556 100450 7568
rect 158898 7556 158904 7568
rect 158956 7556 158962 7608
rect 162394 7556 162400 7608
rect 162452 7596 162458 7608
rect 402514 7596 402520 7608
rect 162452 7568 402520 7596
rect 162452 7556 162458 7568
rect 402514 7556 402520 7568
rect 402572 7556 402578 7608
rect 153010 7488 153016 7540
rect 153068 7528 153074 7540
rect 363506 7528 363512 7540
rect 153068 7500 363512 7528
rect 153068 7488 153074 7500
rect 363506 7488 363512 7500
rect 363564 7488 363570 7540
rect 151538 7420 151544 7472
rect 151596 7460 151602 7472
rect 359918 7460 359924 7472
rect 151596 7432 359924 7460
rect 151596 7420 151602 7432
rect 359918 7420 359924 7432
rect 359976 7420 359982 7472
rect 150066 7352 150072 7404
rect 150124 7392 150130 7404
rect 356330 7392 356336 7404
rect 150124 7364 356336 7392
rect 150124 7352 150130 7364
rect 356330 7352 356336 7364
rect 356388 7352 356394 7404
rect 150158 7284 150164 7336
rect 150216 7324 150222 7336
rect 352834 7324 352840 7336
rect 150216 7296 352840 7324
rect 150216 7284 150222 7296
rect 352834 7284 352840 7296
rect 352892 7284 352898 7336
rect 147490 7216 147496 7268
rect 147548 7256 147554 7268
rect 345750 7256 345756 7268
rect 147548 7228 345756 7256
rect 147548 7216 147554 7228
rect 345750 7216 345756 7228
rect 345808 7216 345814 7268
rect 147398 7148 147404 7200
rect 147456 7188 147462 7200
rect 342162 7188 342168 7200
rect 147456 7160 342168 7188
rect 147456 7148 147462 7160
rect 342162 7148 342168 7160
rect 342220 7148 342226 7200
rect 146202 7080 146208 7132
rect 146260 7120 146266 7132
rect 338666 7120 338672 7132
rect 146260 7092 338672 7120
rect 146260 7080 146266 7092
rect 338666 7080 338672 7092
rect 338724 7080 338730 7132
rect 144822 7012 144828 7064
rect 144880 7052 144886 7064
rect 335078 7052 335084 7064
rect 144880 7024 335084 7052
rect 144880 7012 144886 7024
rect 335078 7012 335084 7024
rect 335136 7012 335142 7064
rect 128262 6808 128268 6860
rect 128320 6848 128326 6860
rect 267734 6848 267740 6860
rect 128320 6820 267740 6848
rect 128320 6808 128326 6820
rect 267734 6808 267740 6820
rect 267792 6808 267798 6860
rect 129458 6740 129464 6792
rect 129516 6780 129522 6792
rect 270402 6780 270408 6792
rect 129516 6752 270408 6780
rect 129516 6740 129522 6752
rect 270402 6740 270408 6752
rect 270460 6740 270466 6792
rect 129642 6672 129648 6724
rect 129700 6712 129706 6724
rect 274818 6712 274824 6724
rect 129700 6684 274824 6712
rect 129700 6672 129706 6684
rect 274818 6672 274824 6684
rect 274876 6672 274882 6724
rect 131022 6604 131028 6656
rect 131080 6644 131086 6656
rect 278314 6644 278320 6656
rect 131080 6616 278320 6644
rect 131080 6604 131086 6616
rect 278314 6604 278320 6616
rect 278372 6604 278378 6656
rect 132310 6536 132316 6588
rect 132368 6576 132374 6588
rect 281902 6576 281908 6588
rect 132368 6548 281908 6576
rect 132368 6536 132374 6548
rect 281902 6536 281908 6548
rect 281960 6536 281966 6588
rect 132218 6468 132224 6520
rect 132276 6508 132282 6520
rect 285398 6508 285404 6520
rect 132276 6480 285404 6508
rect 132276 6468 132282 6480
rect 285398 6468 285404 6480
rect 285456 6468 285462 6520
rect 133782 6400 133788 6452
rect 133840 6440 133846 6452
rect 288986 6440 288992 6452
rect 133840 6412 288992 6440
rect 133840 6400 133846 6412
rect 288986 6400 288992 6412
rect 289044 6400 289050 6452
rect 135070 6332 135076 6384
rect 135128 6372 135134 6384
rect 292574 6372 292580 6384
rect 135128 6344 292580 6372
rect 135128 6332 135134 6344
rect 292574 6332 292580 6344
rect 292632 6332 292638 6384
rect 93670 6264 93676 6316
rect 93728 6304 93734 6316
rect 130562 6304 130568 6316
rect 93728 6276 130568 6304
rect 93728 6264 93734 6276
rect 130562 6264 130568 6276
rect 130620 6264 130626 6316
rect 134978 6264 134984 6316
rect 135036 6304 135042 6316
rect 296070 6304 296076 6316
rect 135036 6276 296076 6304
rect 135036 6264 135042 6276
rect 296070 6264 296076 6276
rect 296128 6264 296134 6316
rect 95050 6196 95056 6248
rect 95108 6236 95114 6248
rect 134150 6236 134156 6248
rect 95108 6208 134156 6236
rect 95108 6196 95114 6208
rect 134150 6196 134156 6208
rect 134208 6196 134214 6248
rect 136542 6196 136548 6248
rect 136600 6236 136606 6248
rect 299658 6236 299664 6248
rect 136600 6208 299664 6236
rect 136600 6196 136606 6208
rect 299658 6196 299664 6208
rect 299716 6196 299722 6248
rect 83826 6128 83832 6180
rect 83884 6168 83890 6180
rect 93946 6168 93952 6180
rect 83884 6140 93952 6168
rect 83884 6128 83890 6140
rect 93946 6128 93952 6140
rect 94004 6128 94010 6180
rect 129550 6128 129556 6180
rect 129608 6168 129614 6180
rect 271230 6168 271236 6180
rect 129608 6140 271236 6168
rect 129608 6128 129614 6140
rect 271230 6128 271236 6140
rect 271288 6128 271294 6180
rect 447410 6168 447416 6180
rect 277366 6140 447416 6168
rect 126882 6060 126888 6112
rect 126940 6100 126946 6112
rect 264146 6100 264152 6112
rect 126940 6072 264152 6100
rect 126940 6060 126946 6072
rect 264146 6060 264152 6072
rect 264204 6060 264210 6112
rect 271138 6060 271144 6112
rect 271196 6100 271202 6112
rect 277366 6100 277394 6140
rect 447410 6128 447416 6140
rect 447468 6128 447474 6180
rect 271196 6072 277394 6100
rect 271196 6060 271202 6072
rect 126790 5992 126796 6044
rect 126848 6032 126854 6044
rect 260650 6032 260656 6044
rect 126848 6004 260656 6032
rect 126848 5992 126854 6004
rect 260650 5992 260656 6004
rect 260708 5992 260714 6044
rect 125226 5924 125232 5976
rect 125284 5964 125290 5976
rect 257062 5964 257068 5976
rect 125284 5936 257068 5964
rect 125284 5924 125290 5936
rect 257062 5924 257068 5936
rect 257120 5924 257126 5976
rect 124030 5856 124036 5908
rect 124088 5896 124094 5908
rect 253474 5896 253480 5908
rect 124088 5868 253480 5896
rect 124088 5856 124094 5868
rect 253474 5856 253480 5868
rect 253532 5856 253538 5908
rect 124122 5788 124128 5840
rect 124180 5828 124186 5840
rect 249978 5828 249984 5840
rect 124180 5800 249984 5828
rect 124180 5788 124186 5800
rect 249978 5788 249984 5800
rect 250036 5788 250042 5840
rect 122650 5720 122656 5772
rect 122708 5760 122714 5772
rect 246390 5760 246396 5772
rect 122708 5732 246396 5760
rect 122708 5720 122714 5732
rect 246390 5720 246396 5732
rect 246448 5720 246454 5772
rect 122742 5652 122748 5704
rect 122800 5692 122806 5704
rect 242986 5692 242992 5704
rect 122800 5664 242992 5692
rect 122800 5652 122806 5664
rect 242986 5652 242992 5664
rect 243044 5652 243050 5704
rect 121362 5584 121368 5636
rect 121420 5624 121426 5636
rect 239306 5624 239312 5636
rect 121420 5596 239312 5624
rect 121420 5584 121426 5596
rect 239306 5584 239312 5596
rect 239364 5584 239370 5636
rect 119706 5516 119712 5568
rect 119764 5556 119770 5568
rect 235810 5556 235816 5568
rect 119764 5528 235816 5556
rect 119764 5516 119770 5528
rect 235810 5516 235816 5528
rect 235868 5516 235874 5568
rect 101766 5448 101772 5500
rect 101824 5488 101830 5500
rect 166074 5488 166080 5500
rect 101824 5460 166080 5488
rect 101824 5448 101830 5460
rect 166074 5448 166080 5460
rect 166132 5448 166138 5500
rect 197262 5448 197268 5500
rect 197320 5488 197326 5500
rect 540790 5488 540796 5500
rect 197320 5460 540796 5488
rect 197320 5448 197326 5460
rect 540790 5448 540796 5460
rect 540848 5448 540854 5500
rect 103422 5380 103428 5432
rect 103480 5420 103486 5432
rect 169570 5420 169576 5432
rect 103480 5392 169576 5420
rect 103480 5380 103486 5392
rect 169570 5380 169576 5392
rect 169628 5380 169634 5432
rect 198642 5380 198648 5432
rect 198700 5420 198706 5432
rect 544286 5420 544292 5432
rect 198700 5392 544292 5420
rect 198700 5380 198706 5392
rect 544286 5380 544292 5392
rect 544344 5380 544350 5432
rect 104710 5312 104716 5364
rect 104768 5352 104774 5364
rect 173158 5352 173164 5364
rect 104768 5324 173164 5352
rect 104768 5312 104774 5324
rect 173158 5312 173164 5324
rect 173216 5312 173222 5364
rect 199654 5312 199660 5364
rect 199712 5352 199718 5364
rect 547966 5352 547972 5364
rect 199712 5324 547972 5352
rect 199712 5312 199718 5324
rect 547966 5312 547972 5324
rect 548024 5312 548030 5364
rect 102778 5244 102784 5296
rect 102836 5284 102842 5296
rect 103422 5284 103428 5296
rect 102836 5256 103428 5284
rect 102836 5244 102842 5256
rect 103422 5244 103428 5256
rect 103480 5244 103486 5296
rect 104618 5244 104624 5296
rect 104676 5284 104682 5296
rect 176654 5284 176660 5296
rect 104676 5256 176660 5284
rect 104676 5244 104682 5256
rect 176654 5244 176660 5256
rect 176712 5244 176718 5296
rect 199930 5244 199936 5296
rect 199988 5284 199994 5296
rect 551462 5284 551468 5296
rect 199988 5256 551468 5284
rect 199988 5244 199994 5256
rect 551462 5244 551468 5256
rect 551520 5244 551526 5296
rect 106090 5176 106096 5228
rect 106148 5216 106154 5228
rect 180242 5216 180248 5228
rect 106148 5188 180248 5216
rect 106148 5176 106154 5188
rect 180242 5176 180248 5188
rect 180300 5176 180306 5228
rect 202414 5176 202420 5228
rect 202472 5216 202478 5228
rect 202472 5188 205772 5216
rect 202472 5176 202478 5188
rect 107562 5108 107568 5160
rect 107620 5148 107626 5160
rect 183738 5148 183744 5160
rect 107620 5120 183744 5148
rect 107620 5108 107626 5120
rect 183738 5108 183744 5120
rect 183796 5108 183802 5160
rect 202690 5108 202696 5160
rect 202748 5148 202754 5160
rect 205744 5148 205772 5188
rect 205818 5176 205824 5228
rect 205876 5216 205882 5228
rect 554958 5216 554964 5228
rect 205876 5188 554964 5216
rect 205876 5176 205882 5188
rect 554958 5176 554964 5188
rect 555016 5176 555022 5228
rect 558546 5148 558552 5160
rect 202748 5120 205680 5148
rect 205744 5120 558552 5148
rect 202748 5108 202754 5120
rect 108850 5040 108856 5092
rect 108908 5080 108914 5092
rect 189718 5080 189724 5092
rect 108908 5052 189724 5080
rect 108908 5040 108914 5052
rect 189718 5040 189724 5052
rect 189776 5040 189782 5092
rect 203886 5040 203892 5092
rect 203944 5080 203950 5092
rect 205652 5080 205680 5120
rect 558546 5108 558552 5120
rect 558604 5108 558610 5160
rect 562042 5080 562048 5092
rect 203944 5052 205220 5080
rect 205652 5052 562048 5080
rect 203944 5040 203950 5052
rect 108942 4972 108948 5024
rect 109000 5012 109006 5024
rect 193306 5012 193312 5024
rect 109000 4984 193312 5012
rect 109000 4972 109006 4984
rect 193306 4972 193312 4984
rect 193364 4972 193370 5024
rect 194226 4972 194232 5024
rect 194284 5012 194290 5024
rect 204990 5012 204996 5024
rect 194284 4984 204996 5012
rect 194284 4972 194290 4984
rect 204990 4972 204996 4984
rect 205048 4972 205054 5024
rect 205192 5012 205220 5052
rect 562042 5040 562048 5052
rect 562100 5040 562106 5092
rect 565630 5012 565636 5024
rect 205192 4984 565636 5012
rect 565630 4972 565636 4984
rect 565688 4972 565694 5024
rect 110322 4904 110328 4956
rect 110380 4944 110386 4956
rect 196802 4944 196808 4956
rect 110380 4916 196808 4944
rect 110380 4904 110386 4916
rect 196802 4904 196808 4916
rect 196860 4904 196866 4956
rect 204070 4904 204076 4956
rect 204128 4944 204134 4956
rect 569126 4944 569132 4956
rect 204128 4916 569132 4944
rect 204128 4904 204134 4916
rect 569126 4904 569132 4916
rect 569184 4904 569190 4956
rect 111702 4836 111708 4888
rect 111760 4876 111766 4888
rect 200298 4876 200304 4888
rect 111760 4848 200304 4876
rect 111760 4836 111766 4848
rect 200298 4836 200304 4848
rect 200356 4836 200362 4888
rect 201402 4836 201408 4888
rect 201460 4876 201466 4888
rect 201460 4848 204024 4876
rect 201460 4836 201466 4848
rect 111610 4768 111616 4820
rect 111668 4808 111674 4820
rect 203886 4808 203892 4820
rect 111668 4780 203892 4808
rect 111668 4768 111674 4780
rect 203886 4768 203892 4780
rect 203944 4768 203950 4820
rect 203996 4808 204024 4848
rect 205542 4836 205548 4888
rect 205600 4876 205606 4888
rect 572806 4876 572812 4888
rect 205600 4848 572812 4876
rect 205600 4836 205606 4848
rect 572806 4836 572812 4848
rect 572864 4836 572870 4888
rect 205818 4808 205824 4820
rect 203996 4780 205824 4808
rect 205818 4768 205824 4780
rect 205876 4768 205882 4820
rect 206922 4768 206928 4820
rect 206980 4808 206986 4820
rect 576302 4808 576308 4820
rect 206980 4780 576308 4808
rect 206980 4768 206986 4780
rect 576302 4768 576308 4780
rect 576360 4768 576366 4820
rect 101858 4700 101864 4752
rect 101916 4740 101922 4752
rect 162486 4740 162492 4752
rect 101916 4712 162492 4740
rect 101916 4700 101922 4712
rect 162486 4700 162492 4712
rect 162544 4700 162550 4752
rect 197170 4700 197176 4752
rect 197228 4740 197234 4752
rect 537202 4740 537208 4752
rect 197228 4712 537208 4740
rect 197228 4700 197234 4712
rect 537202 4700 537208 4712
rect 537260 4700 537266 4752
rect 100478 4632 100484 4684
rect 100536 4672 100542 4684
rect 157794 4672 157800 4684
rect 100536 4644 157800 4672
rect 100536 4632 100542 4644
rect 157794 4632 157800 4644
rect 157852 4632 157858 4684
rect 533706 4672 533712 4684
rect 200086 4644 533712 4672
rect 99098 4564 99104 4616
rect 99156 4604 99162 4616
rect 154206 4604 154212 4616
rect 99156 4576 154212 4604
rect 99156 4564 99162 4576
rect 154206 4564 154212 4576
rect 154264 4564 154270 4616
rect 195514 4564 195520 4616
rect 195572 4604 195578 4616
rect 200086 4604 200114 4644
rect 533706 4632 533712 4644
rect 533764 4632 533770 4684
rect 530118 4604 530124 4616
rect 195572 4576 200114 4604
rect 204916 4576 530124 4604
rect 195572 4564 195578 4576
rect 97718 4496 97724 4548
rect 97776 4536 97782 4548
rect 147122 4536 147128 4548
rect 97776 4508 147128 4536
rect 97776 4496 97782 4508
rect 147122 4496 147128 4508
rect 147180 4496 147186 4548
rect 194502 4496 194508 4548
rect 194560 4536 194566 4548
rect 204916 4536 204944 4576
rect 530118 4564 530124 4576
rect 530176 4564 530182 4616
rect 194560 4508 204944 4536
rect 194560 4496 194566 4508
rect 204990 4496 204996 4548
rect 205048 4536 205054 4548
rect 526622 4536 526628 4548
rect 205048 4508 526628 4536
rect 205048 4496 205054 4508
rect 526622 4496 526628 4508
rect 526680 4496 526686 4548
rect 96430 4428 96436 4480
rect 96488 4468 96494 4480
rect 143534 4468 143540 4480
rect 96488 4440 143540 4468
rect 96488 4428 96494 4440
rect 143534 4428 143540 4440
rect 143592 4428 143598 4480
rect 192754 4428 192760 4480
rect 192812 4468 192818 4480
rect 523034 4468 523040 4480
rect 192812 4440 523040 4468
rect 192812 4428 192818 4440
rect 523034 4428 523040 4440
rect 523092 4428 523098 4480
rect 95142 4360 95148 4412
rect 95200 4400 95206 4412
rect 136450 4400 136456 4412
rect 95200 4372 136456 4400
rect 95200 4360 95206 4372
rect 136450 4360 136456 4372
rect 136508 4360 136514 4412
rect 141418 4360 141424 4412
rect 141476 4400 141482 4412
rect 186130 4400 186136 4412
rect 141476 4372 186136 4400
rect 141476 4360 141482 4372
rect 186130 4360 186136 4372
rect 186188 4360 186194 4412
rect 191466 4360 191472 4412
rect 191524 4400 191530 4412
rect 519538 4400 519544 4412
rect 191524 4372 519544 4400
rect 191524 4360 191530 4372
rect 519538 4360 519544 4372
rect 519596 4360 519602 4412
rect 93762 4292 93768 4344
rect 93820 4332 93826 4344
rect 132954 4332 132960 4344
rect 93820 4304 132960 4332
rect 93820 4292 93826 4304
rect 132954 4292 132960 4304
rect 133012 4292 133018 4344
rect 191650 4292 191656 4344
rect 191708 4332 191714 4344
rect 515950 4332 515956 4344
rect 191708 4304 515956 4332
rect 191708 4292 191714 4304
rect 515950 4292 515956 4304
rect 516008 4292 516014 4344
rect 92290 4224 92296 4276
rect 92348 4264 92354 4276
rect 126974 4264 126980 4276
rect 92348 4236 126980 4264
rect 92348 4224 92354 4236
rect 126974 4224 126980 4236
rect 127032 4224 127038 4276
rect 190086 4224 190092 4276
rect 190144 4264 190150 4276
rect 512454 4264 512460 4276
rect 190144 4236 512460 4264
rect 190144 4224 190150 4236
rect 512454 4224 512460 4236
rect 512512 4224 512518 4276
rect 276014 4156 276020 4208
rect 276072 4196 276078 4208
rect 277118 4196 277124 4208
rect 276072 4168 277124 4196
rect 276072 4156 276078 4168
rect 277118 4156 277124 4168
rect 277176 4156 277182 4208
rect 28902 4088 28908 4140
rect 28960 4128 28966 4140
rect 52454 4128 52460 4140
rect 28960 4100 52460 4128
rect 28960 4088 28966 4100
rect 52454 4088 52460 4100
rect 52512 4088 52518 4140
rect 52546 4088 52552 4140
rect 52604 4128 52610 4140
rect 53650 4128 53656 4140
rect 52604 4100 53656 4128
rect 52604 4088 52610 4100
rect 53650 4088 53656 4100
rect 53708 4088 53714 4140
rect 56042 4088 56048 4140
rect 56100 4128 56106 4140
rect 57238 4128 57244 4140
rect 56100 4100 57244 4128
rect 56100 4088 56106 4100
rect 57238 4088 57244 4100
rect 57296 4088 57302 4140
rect 58434 4088 58440 4140
rect 58492 4128 58498 4140
rect 59262 4128 59268 4140
rect 58492 4100 59268 4128
rect 58492 4088 58498 4100
rect 59262 4088 59268 4100
rect 59320 4088 59326 4140
rect 59630 4088 59636 4140
rect 59688 4128 59694 4140
rect 60642 4128 60648 4140
rect 59688 4100 60648 4128
rect 59688 4088 59694 4100
rect 60642 4088 60648 4100
rect 60700 4088 60706 4140
rect 82446 4088 82452 4140
rect 82504 4128 82510 4140
rect 85666 4128 85672 4140
rect 82504 4100 85672 4128
rect 82504 4088 82510 4100
rect 85666 4088 85672 4100
rect 85724 4088 85730 4140
rect 91002 4088 91008 4140
rect 91060 4128 91066 4140
rect 117590 4128 117596 4140
rect 91060 4100 117596 4128
rect 91060 4088 91066 4100
rect 117590 4088 117596 4100
rect 117648 4088 117654 4140
rect 139302 4088 139308 4140
rect 139360 4128 139366 4140
rect 309042 4128 309048 4140
rect 139360 4100 309048 4128
rect 139360 4088 139366 4100
rect 309042 4088 309048 4100
rect 309100 4088 309106 4140
rect 421558 4088 421564 4140
rect 421616 4128 421622 4140
rect 423674 4128 423680 4140
rect 421616 4100 423680 4128
rect 421616 4088 421622 4100
rect 423674 4088 423680 4100
rect 423732 4088 423738 4140
rect 439498 4088 439504 4140
rect 439556 4128 439562 4140
rect 442626 4128 442632 4140
rect 439556 4100 442632 4128
rect 439556 4088 439562 4100
rect 442626 4088 442632 4100
rect 442684 4088 442690 4140
rect 472618 4088 472624 4140
rect 472676 4128 472682 4140
rect 510062 4128 510068 4140
rect 472676 4100 510068 4128
rect 472676 4088 472682 4100
rect 510062 4088 510068 4100
rect 510120 4088 510126 4140
rect 23014 4020 23020 4072
rect 23072 4060 23078 4072
rect 65702 4060 65708 4072
rect 23072 4032 65708 4060
rect 23072 4020 23078 4032
rect 65702 4020 65708 4032
rect 65760 4020 65766 4072
rect 71498 4020 71504 4072
rect 71556 4060 71562 4072
rect 76558 4060 76564 4072
rect 71556 4032 76564 4060
rect 71556 4020 71562 4032
rect 76558 4020 76564 4032
rect 76616 4020 76622 4072
rect 90726 4020 90732 4072
rect 90784 4060 90790 4072
rect 118786 4060 118792 4072
rect 90784 4032 118792 4060
rect 90784 4020 90790 4032
rect 118786 4020 118792 4032
rect 118844 4020 118850 4072
rect 144546 4020 144552 4072
rect 144604 4060 144610 4072
rect 333882 4060 333888 4072
rect 144604 4032 333888 4060
rect 144604 4020 144610 4032
rect 333882 4020 333888 4032
rect 333940 4020 333946 4072
rect 479518 4020 479524 4072
rect 479576 4060 479582 4072
rect 517146 4060 517152 4072
rect 479576 4032 517152 4060
rect 479576 4020 479582 4032
rect 517146 4020 517152 4032
rect 517204 4020 517210 4072
rect 19426 3952 19432 4004
rect 19484 3992 19490 4004
rect 27614 3992 27620 4004
rect 19484 3964 27620 3992
rect 19484 3952 19490 3964
rect 27614 3952 27620 3964
rect 27672 3952 27678 4004
rect 65150 3992 65156 4004
rect 27724 3964 65156 3992
rect 20622 3884 20628 3936
rect 20680 3924 20686 3936
rect 27724 3924 27752 3964
rect 65150 3952 65156 3964
rect 65208 3952 65214 4004
rect 88058 3952 88064 4004
rect 88116 3992 88122 4004
rect 111610 3992 111616 4004
rect 88116 3964 111616 3992
rect 88116 3952 88122 3964
rect 111610 3952 111616 3964
rect 111668 3952 111674 4004
rect 113082 3952 113088 4004
rect 113140 3992 113146 4004
rect 201402 3992 201408 4004
rect 113140 3964 201408 3992
rect 113140 3952 113146 3964
rect 201402 3952 201408 3964
rect 201460 3952 201466 4004
rect 201494 3952 201500 4004
rect 201552 3992 201558 4004
rect 202690 3992 202696 4004
rect 201552 3964 202696 3992
rect 201552 3952 201558 3964
rect 202690 3952 202696 3964
rect 202748 3952 202754 4004
rect 218974 3952 218980 4004
rect 219032 3992 219038 4004
rect 408402 3992 408408 4004
rect 219032 3964 408408 3992
rect 219032 3952 219038 3964
rect 408402 3952 408408 3964
rect 408460 3952 408466 4004
rect 468478 3952 468484 4004
rect 468536 3992 468542 4004
rect 506474 3992 506480 4004
rect 468536 3964 506480 3992
rect 468536 3952 468542 3964
rect 506474 3952 506480 3964
rect 506532 3952 506538 4004
rect 20680 3896 27752 3924
rect 20680 3884 20686 3896
rect 27798 3884 27804 3936
rect 27856 3924 27862 3936
rect 64966 3924 64972 3936
rect 27856 3896 64972 3924
rect 27856 3884 27862 3896
rect 64966 3884 64972 3896
rect 65024 3884 65030 3936
rect 89622 3884 89628 3936
rect 89680 3924 89686 3936
rect 116394 3924 116400 3936
rect 89680 3896 116400 3924
rect 89680 3884 89686 3896
rect 116394 3884 116400 3896
rect 116452 3884 116458 3936
rect 147582 3884 147588 3936
rect 147640 3924 147646 3936
rect 344554 3924 344560 3936
rect 147640 3896 344560 3924
rect 147640 3884 147646 3896
rect 344554 3884 344560 3896
rect 344612 3884 344618 3936
rect 447778 3884 447784 3936
rect 447836 3924 447842 3936
rect 491110 3924 491116 3936
rect 447836 3896 491116 3924
rect 447836 3884 447842 3896
rect 491110 3884 491116 3896
rect 491168 3884 491174 3936
rect 18230 3816 18236 3868
rect 18288 3856 18294 3868
rect 52362 3856 52368 3868
rect 18288 3828 52368 3856
rect 18288 3816 18294 3828
rect 52362 3816 52368 3828
rect 52420 3816 52426 3868
rect 52454 3816 52460 3868
rect 52512 3856 52518 3868
rect 52512 3828 56088 3856
rect 52512 3816 52518 3828
rect 15930 3748 15936 3800
rect 15988 3788 15994 3800
rect 56060 3788 56088 3828
rect 56134 3816 56140 3868
rect 56192 3856 56198 3868
rect 61838 3856 61844 3868
rect 56192 3828 61844 3856
rect 56192 3816 56198 3828
rect 61838 3816 61844 3828
rect 61896 3816 61902 3868
rect 90634 3816 90640 3868
rect 90692 3856 90698 3868
rect 119890 3856 119896 3868
rect 90692 3828 119896 3856
rect 90692 3816 90698 3828
rect 119890 3816 119896 3828
rect 119948 3816 119954 3868
rect 150250 3816 150256 3868
rect 150308 3856 150314 3868
rect 351638 3856 351644 3868
rect 150308 3828 351644 3856
rect 150308 3816 150314 3828
rect 351638 3816 351644 3828
rect 351696 3816 351702 3868
rect 425698 3816 425704 3868
rect 425756 3856 425762 3868
rect 468662 3856 468668 3868
rect 425756 3828 468668 3856
rect 425756 3816 425762 3828
rect 468662 3816 468668 3828
rect 468720 3816 468726 3868
rect 475378 3816 475384 3868
rect 475436 3856 475442 3868
rect 513558 3856 513564 3868
rect 475436 3828 513564 3856
rect 475436 3816 475442 3828
rect 513558 3816 513564 3828
rect 513616 3816 513622 3868
rect 67266 3788 67272 3800
rect 15988 3760 55904 3788
rect 56060 3760 67272 3788
rect 15988 3748 15994 3760
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 55490 3720 55496 3732
rect 12308 3692 55496 3720
rect 12308 3680 12314 3692
rect 55490 3680 55496 3692
rect 55548 3680 55554 3732
rect 55876 3720 55904 3760
rect 67266 3748 67272 3760
rect 67324 3748 67330 3800
rect 82630 3748 82636 3800
rect 82688 3788 82694 3800
rect 87966 3788 87972 3800
rect 82688 3760 87972 3788
rect 82688 3748 82694 3760
rect 87966 3748 87972 3760
rect 88024 3748 88030 3800
rect 90910 3748 90916 3800
rect 90968 3788 90974 3800
rect 121086 3788 121092 3800
rect 90968 3760 121092 3788
rect 90968 3748 90974 3760
rect 121086 3748 121092 3760
rect 121144 3748 121150 3800
rect 122098 3748 122104 3800
rect 122156 3788 122162 3800
rect 128170 3788 128176 3800
rect 122156 3760 128176 3788
rect 122156 3748 122162 3760
rect 128170 3748 128176 3760
rect 128228 3748 128234 3800
rect 150342 3748 150348 3800
rect 150400 3788 150406 3800
rect 355226 3788 355232 3800
rect 150400 3760 355232 3788
rect 150400 3748 150406 3760
rect 355226 3748 355232 3760
rect 355284 3748 355290 3800
rect 418798 3748 418804 3800
rect 418856 3788 418862 3800
rect 461578 3788 461584 3800
rect 418856 3760 461584 3788
rect 418856 3748 418862 3760
rect 461578 3748 461584 3760
rect 461636 3748 461642 3800
rect 461670 3748 461676 3800
rect 461728 3788 461734 3800
rect 505370 3788 505376 3800
rect 461728 3760 505376 3788
rect 461728 3748 461734 3760
rect 505370 3748 505376 3760
rect 505428 3748 505434 3800
rect 63954 3720 63960 3732
rect 55876 3692 63960 3720
rect 63954 3680 63960 3692
rect 64012 3680 64018 3732
rect 84010 3680 84016 3732
rect 84068 3720 84074 3732
rect 90358 3720 90364 3732
rect 84068 3692 90364 3720
rect 84068 3680 84074 3692
rect 90358 3680 90364 3692
rect 90416 3680 90422 3732
rect 90818 3680 90824 3732
rect 90876 3720 90882 3732
rect 122282 3720 122288 3732
rect 90876 3692 122288 3720
rect 90876 3680 90882 3692
rect 122282 3680 122288 3692
rect 122340 3680 122346 3732
rect 160002 3680 160008 3732
rect 160060 3720 160066 3732
rect 394234 3720 394240 3732
rect 160060 3692 394240 3720
rect 160060 3680 160066 3692
rect 394234 3680 394240 3692
rect 394292 3680 394298 3732
rect 411990 3680 411996 3732
rect 412048 3720 412054 3732
rect 454494 3720 454500 3732
rect 412048 3692 454500 3720
rect 412048 3680 412054 3692
rect 454494 3680 454500 3692
rect 454552 3680 454558 3732
rect 454678 3680 454684 3732
rect 454736 3720 454742 3732
rect 498194 3720 498200 3732
rect 454736 3692 498200 3720
rect 454736 3680 454742 3692
rect 498194 3680 498200 3692
rect 498252 3680 498258 3732
rect 537478 3680 537484 3732
rect 537536 3720 537542 3732
rect 557350 3720 557356 3732
rect 537536 3692 557356 3720
rect 537536 3680 537542 3692
rect 557350 3680 557356 3692
rect 557408 3680 557414 3732
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 56134 3652 56140 3664
rect 7708 3624 56140 3652
rect 7708 3612 7714 3624
rect 56134 3612 56140 3624
rect 56192 3612 56198 3664
rect 61286 3652 61292 3664
rect 60706 3624 61292 3652
rect 1670 3544 1676 3596
rect 1728 3584 1734 3596
rect 1728 3556 4200 3584
rect 1728 3544 1734 3556
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 3970 3516 3976 3528
rect 2924 3488 3976 3516
rect 2924 3476 2930 3488
rect 3970 3476 3976 3488
rect 4028 3476 4034 3528
rect 4172 3516 4200 3556
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 60706 3584 60734 3624
rect 61286 3612 61292 3624
rect 61344 3612 61350 3664
rect 82538 3612 82544 3664
rect 82596 3652 82602 3664
rect 89162 3652 89168 3664
rect 82596 3624 89168 3652
rect 82596 3612 82602 3624
rect 89162 3612 89168 3624
rect 89220 3612 89226 3664
rect 92382 3612 92388 3664
rect 92440 3652 92446 3664
rect 124674 3652 124680 3664
rect 92440 3624 124680 3652
rect 92440 3612 92446 3624
rect 124674 3612 124680 3624
rect 124732 3612 124738 3664
rect 138658 3612 138664 3664
rect 138716 3652 138722 3664
rect 140038 3652 140044 3664
rect 138716 3624 140044 3652
rect 138716 3612 138722 3624
rect 140038 3612 140044 3624
rect 140096 3612 140102 3664
rect 161382 3612 161388 3664
rect 161440 3652 161446 3664
rect 397730 3652 397736 3664
rect 161440 3624 397736 3652
rect 161440 3612 161446 3624
rect 397730 3612 397736 3624
rect 397788 3612 397794 3664
rect 443638 3612 443644 3664
rect 443696 3652 443702 3664
rect 443696 3624 449940 3652
rect 443696 3612 443702 3624
rect 5316 3556 60734 3584
rect 5316 3544 5322 3556
rect 64322 3544 64328 3596
rect 64380 3584 64386 3596
rect 64782 3584 64788 3596
rect 64380 3556 64788 3584
rect 64380 3544 64386 3556
rect 64782 3544 64788 3556
rect 64840 3544 64846 3596
rect 72418 3584 72424 3596
rect 65444 3556 72424 3584
rect 55214 3516 55220 3528
rect 4172 3488 55220 3516
rect 55214 3476 55220 3488
rect 55272 3476 55278 3528
rect 55490 3476 55496 3528
rect 55548 3516 55554 3528
rect 59998 3516 60004 3528
rect 55548 3488 60004 3516
rect 55548 3476 55554 3488
rect 59998 3476 60004 3488
rect 60056 3476 60062 3528
rect 63218 3476 63224 3528
rect 63276 3516 63282 3528
rect 65444 3516 65472 3556
rect 72418 3544 72424 3556
rect 72476 3544 72482 3596
rect 74994 3544 75000 3596
rect 75052 3584 75058 3596
rect 75822 3584 75828 3596
rect 75052 3556 75828 3584
rect 75052 3544 75058 3556
rect 75822 3544 75828 3556
rect 75880 3544 75886 3596
rect 81342 3544 81348 3596
rect 81400 3584 81406 3596
rect 81400 3556 82400 3584
rect 81400 3544 81406 3556
rect 63276 3488 65472 3516
rect 63276 3476 63282 3488
rect 65518 3476 65524 3528
rect 65576 3516 65582 3528
rect 66162 3516 66168 3528
rect 65576 3488 66168 3516
rect 65576 3476 65582 3488
rect 66162 3476 66168 3488
rect 66220 3476 66226 3528
rect 66714 3476 66720 3528
rect 66772 3516 66778 3528
rect 67542 3516 67548 3528
rect 66772 3488 67548 3516
rect 66772 3476 66778 3488
rect 67542 3476 67548 3488
rect 67600 3476 67606 3528
rect 67910 3476 67916 3528
rect 67968 3516 67974 3528
rect 68922 3516 68928 3528
rect 67968 3488 68928 3516
rect 67968 3476 67974 3488
rect 68922 3476 68928 3488
rect 68980 3476 68986 3528
rect 69106 3476 69112 3528
rect 69164 3516 69170 3528
rect 70210 3516 70216 3528
rect 69164 3488 70216 3516
rect 69164 3476 69170 3488
rect 70210 3476 70216 3488
rect 70268 3476 70274 3528
rect 72602 3476 72608 3528
rect 72660 3516 72666 3528
rect 73062 3516 73068 3528
rect 72660 3488 73068 3516
rect 72660 3476 72666 3488
rect 73062 3476 73068 3488
rect 73120 3476 73126 3528
rect 75362 3516 75368 3528
rect 73172 3488 75368 3516
rect 566 3408 572 3460
rect 624 3448 630 3460
rect 59354 3448 59360 3460
rect 624 3420 59360 3448
rect 624 3408 630 3420
rect 59354 3408 59360 3420
rect 59412 3408 59418 3460
rect 60826 3408 60832 3460
rect 60884 3448 60890 3460
rect 73172 3448 73200 3488
rect 75362 3476 75368 3488
rect 75420 3476 75426 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 79686 3476 79692 3528
rect 79744 3516 79750 3528
rect 80330 3516 80336 3528
rect 79744 3488 80336 3516
rect 79744 3476 79750 3488
rect 80330 3476 80336 3488
rect 80388 3476 80394 3528
rect 80422 3476 80428 3528
rect 80480 3516 80486 3528
rect 80882 3516 80888 3528
rect 80480 3488 80888 3516
rect 80480 3476 80486 3488
rect 80882 3476 80888 3488
rect 80940 3476 80946 3528
rect 81250 3476 81256 3528
rect 81308 3516 81314 3528
rect 82078 3516 82084 3528
rect 81308 3488 82084 3516
rect 81308 3476 81314 3488
rect 82078 3476 82084 3488
rect 82136 3476 82142 3528
rect 82372 3516 82400 3556
rect 84102 3544 84108 3596
rect 84160 3584 84166 3596
rect 91554 3584 91560 3596
rect 84160 3556 91560 3584
rect 84160 3544 84166 3556
rect 91554 3544 91560 3556
rect 91612 3544 91618 3596
rect 97810 3544 97816 3596
rect 97868 3584 97874 3596
rect 97868 3556 100616 3584
rect 97868 3544 97874 3556
rect 84470 3516 84476 3528
rect 82372 3488 84476 3516
rect 84470 3476 84476 3488
rect 84528 3476 84534 3528
rect 95142 3516 95148 3528
rect 88996 3488 95148 3516
rect 60884 3420 73200 3448
rect 60884 3408 60890 3420
rect 73798 3408 73804 3460
rect 73856 3448 73862 3460
rect 75178 3448 75184 3460
rect 73856 3420 75184 3448
rect 73856 3408 73862 3420
rect 75178 3408 75184 3420
rect 75236 3408 75242 3460
rect 83918 3408 83924 3460
rect 83976 3448 83982 3460
rect 88996 3448 89024 3488
rect 95142 3476 95148 3488
rect 95200 3476 95206 3528
rect 96522 3476 96528 3528
rect 96580 3516 96586 3528
rect 98454 3516 98460 3528
rect 96580 3488 98460 3516
rect 96580 3476 96586 3488
rect 98454 3476 98460 3488
rect 98512 3476 98518 3528
rect 98822 3476 98828 3528
rect 98880 3516 98886 3528
rect 100588 3516 100616 3556
rect 100662 3544 100668 3596
rect 100720 3584 100726 3596
rect 100720 3556 101352 3584
rect 100720 3544 100726 3556
rect 101214 3516 101220 3528
rect 98880 3488 100248 3516
rect 100588 3488 101220 3516
rect 98880 3476 98886 3488
rect 99190 3448 99196 3460
rect 83976 3420 89024 3448
rect 89088 3420 99196 3448
rect 83976 3408 83982 3420
rect 8754 3340 8760 3392
rect 8812 3380 8818 3392
rect 9582 3380 9588 3392
rect 8812 3352 9588 3380
rect 8812 3340 8818 3352
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 9950 3340 9956 3392
rect 10008 3380 10014 3392
rect 10962 3380 10968 3392
rect 10008 3352 10968 3380
rect 10008 3340 10014 3352
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 12342 3380 12348 3392
rect 11204 3352 12348 3380
rect 11204 3340 11210 3352
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 17034 3340 17040 3392
rect 17092 3380 17098 3392
rect 17862 3380 17868 3392
rect 17092 3352 17868 3380
rect 17092 3340 17098 3352
rect 17862 3340 17868 3352
rect 17920 3340 17926 3392
rect 25314 3340 25320 3392
rect 25372 3380 25378 3392
rect 26142 3380 26148 3392
rect 25372 3352 26148 3380
rect 25372 3340 25378 3352
rect 26142 3340 26148 3352
rect 26200 3340 26206 3392
rect 27706 3340 27712 3392
rect 27764 3380 27770 3392
rect 28810 3380 28816 3392
rect 27764 3352 28816 3380
rect 27764 3340 27770 3352
rect 28810 3340 28816 3352
rect 28868 3340 28874 3392
rect 32398 3340 32404 3392
rect 32456 3380 32462 3392
rect 33042 3380 33048 3392
rect 32456 3352 33048 3380
rect 32456 3340 32462 3352
rect 33042 3340 33048 3352
rect 33100 3340 33106 3392
rect 33594 3340 33600 3392
rect 33652 3380 33658 3392
rect 34422 3380 34428 3392
rect 33652 3352 34428 3380
rect 33652 3340 33658 3352
rect 34422 3340 34428 3352
rect 34480 3340 34486 3392
rect 34790 3340 34796 3392
rect 34848 3380 34854 3392
rect 35802 3380 35808 3392
rect 34848 3352 35808 3380
rect 34848 3340 34854 3352
rect 35802 3340 35808 3352
rect 35860 3340 35866 3392
rect 40678 3340 40684 3392
rect 40736 3380 40742 3392
rect 41322 3380 41328 3392
rect 40736 3352 41328 3380
rect 40736 3340 40742 3352
rect 41322 3340 41328 3352
rect 41380 3340 41386 3392
rect 43070 3340 43076 3392
rect 43128 3380 43134 3392
rect 44082 3380 44088 3392
rect 43128 3352 44088 3380
rect 43128 3340 43134 3352
rect 44082 3340 44088 3352
rect 44140 3340 44146 3392
rect 67818 3380 67824 3392
rect 45388 3352 67824 3380
rect 31294 3272 31300 3324
rect 31352 3312 31358 3324
rect 45388 3312 45416 3352
rect 67818 3340 67824 3352
rect 67876 3340 67882 3392
rect 78582 3340 78588 3392
rect 78640 3380 78646 3392
rect 79778 3380 79784 3392
rect 78640 3352 79784 3380
rect 78640 3340 78646 3352
rect 79778 3340 79784 3352
rect 79836 3340 79842 3392
rect 86218 3340 86224 3392
rect 86276 3380 86282 3392
rect 89088 3380 89116 3420
rect 99190 3408 99196 3420
rect 99248 3408 99254 3460
rect 99558 3408 99564 3460
rect 99616 3448 99622 3460
rect 100110 3448 100116 3460
rect 99616 3420 100116 3448
rect 99616 3408 99622 3420
rect 100110 3408 100116 3420
rect 100168 3408 100174 3460
rect 86276 3352 89116 3380
rect 86276 3340 86282 3352
rect 89438 3340 89444 3392
rect 89496 3380 89502 3392
rect 100220 3380 100248 3488
rect 101214 3476 101220 3488
rect 101272 3476 101278 3528
rect 100294 3408 100300 3460
rect 100352 3448 100358 3460
rect 101324 3448 101352 3556
rect 101398 3544 101404 3596
rect 101456 3584 101462 3596
rect 103330 3584 103336 3596
rect 101456 3556 103336 3584
rect 101456 3544 101462 3556
rect 103330 3544 103336 3556
rect 103388 3544 103394 3596
rect 103422 3544 103428 3596
rect 103480 3584 103486 3596
rect 106826 3584 106832 3596
rect 103480 3556 106832 3584
rect 103480 3544 103486 3556
rect 106826 3544 106832 3556
rect 106884 3544 106890 3596
rect 107212 3556 107424 3584
rect 101490 3476 101496 3528
rect 101548 3516 101554 3528
rect 107212 3516 107240 3556
rect 101548 3488 107240 3516
rect 107396 3516 107424 3556
rect 107470 3544 107476 3596
rect 107528 3584 107534 3596
rect 142430 3584 142436 3596
rect 107528 3556 142436 3584
rect 107528 3544 107534 3556
rect 142430 3544 142436 3556
rect 142488 3544 142494 3596
rect 165246 3544 165252 3596
rect 165304 3584 165310 3596
rect 415486 3584 415492 3596
rect 165304 3556 415492 3584
rect 165304 3544 165310 3556
rect 415486 3544 415492 3556
rect 415544 3544 415550 3596
rect 429838 3544 429844 3596
rect 429896 3584 429902 3596
rect 429896 3556 431954 3584
rect 429896 3544 429902 3556
rect 145926 3516 145932 3528
rect 107396 3488 145932 3516
rect 101548 3476 101554 3488
rect 145926 3476 145932 3488
rect 145984 3476 145990 3528
rect 168006 3476 168012 3528
rect 168064 3516 168070 3528
rect 168064 3488 423720 3516
rect 168064 3476 168070 3488
rect 102318 3448 102324 3460
rect 100352 3420 101168 3448
rect 101324 3420 102324 3448
rect 100352 3408 100358 3420
rect 101030 3380 101036 3392
rect 89496 3352 98776 3380
rect 100220 3352 101036 3380
rect 89496 3340 89502 3352
rect 31352 3284 45416 3312
rect 31352 3272 31358 3284
rect 48958 3272 48964 3324
rect 49016 3312 49022 3324
rect 49602 3312 49608 3324
rect 49016 3284 49608 3312
rect 49016 3272 49022 3284
rect 49602 3272 49608 3284
rect 49660 3272 49666 3324
rect 69198 3312 69204 3324
rect 55876 3284 69204 3312
rect 41874 3204 41880 3256
rect 41932 3244 41938 3256
rect 43438 3244 43444 3256
rect 41932 3216 43444 3244
rect 41932 3204 41938 3216
rect 43438 3204 43444 3216
rect 43496 3204 43502 3256
rect 43548 3216 45554 3244
rect 38378 3136 38384 3188
rect 38436 3176 38442 3188
rect 43548 3176 43576 3216
rect 38436 3148 43576 3176
rect 38436 3136 38442 3148
rect 44266 3136 44272 3188
rect 44324 3176 44330 3188
rect 45370 3176 45376 3188
rect 44324 3148 45376 3176
rect 44324 3136 44330 3148
rect 45370 3136 45376 3148
rect 45428 3136 45434 3188
rect 45526 3176 45554 3216
rect 55766 3176 55772 3188
rect 45526 3148 55772 3176
rect 55766 3136 55772 3148
rect 55824 3136 55830 3188
rect 35986 3068 35992 3120
rect 36044 3108 36050 3120
rect 55876 3108 55904 3284
rect 69198 3272 69204 3284
rect 69256 3272 69262 3324
rect 88978 3272 88984 3324
rect 89036 3312 89042 3324
rect 96246 3312 96252 3324
rect 89036 3284 96252 3312
rect 89036 3272 89042 3284
rect 96246 3272 96252 3284
rect 96304 3272 96310 3324
rect 98748 3312 98776 3352
rect 101030 3340 101036 3352
rect 101088 3340 101094 3392
rect 101140 3380 101168 3420
rect 102318 3408 102324 3420
rect 102376 3408 102382 3460
rect 102870 3408 102876 3460
rect 102928 3448 102934 3460
rect 106918 3448 106924 3460
rect 102928 3420 106924 3448
rect 102928 3408 102934 3420
rect 106918 3408 106924 3420
rect 106976 3408 106982 3460
rect 110138 3408 110144 3460
rect 110196 3448 110202 3460
rect 156598 3448 156604 3460
rect 110196 3420 156604 3448
rect 110196 3408 110202 3420
rect 156598 3408 156604 3420
rect 156656 3408 156662 3460
rect 169662 3408 169668 3460
rect 169720 3448 169726 3460
rect 169720 3420 412634 3448
rect 169720 3408 169726 3420
rect 107010 3380 107016 3392
rect 101140 3352 107016 3380
rect 107010 3340 107016 3352
rect 107068 3340 107074 3392
rect 107102 3340 107108 3392
rect 107160 3380 107166 3392
rect 110506 3380 110512 3392
rect 107160 3352 110512 3380
rect 107160 3340 107166 3352
rect 110506 3340 110512 3352
rect 110564 3340 110570 3392
rect 110598 3340 110604 3392
rect 110656 3380 110662 3392
rect 123478 3380 123484 3392
rect 110656 3352 123484 3380
rect 110656 3340 110662 3352
rect 123478 3340 123484 3352
rect 123536 3340 123542 3392
rect 124858 3340 124864 3392
rect 124916 3380 124922 3392
rect 125870 3380 125876 3392
rect 124916 3352 125876 3380
rect 124916 3340 124922 3352
rect 125870 3340 125876 3352
rect 125928 3340 125934 3392
rect 137738 3340 137744 3392
rect 137796 3380 137802 3392
rect 306742 3380 306748 3392
rect 137796 3352 306748 3380
rect 137796 3340 137802 3352
rect 306742 3340 306748 3352
rect 306800 3340 306806 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 347038 3340 347044 3392
rect 347096 3380 347102 3392
rect 349246 3380 349252 3392
rect 347096 3352 349252 3380
rect 347096 3340 347102 3352
rect 349246 3340 349252 3352
rect 349304 3340 349310 3392
rect 373994 3340 374000 3392
rect 374052 3380 374058 3392
rect 375282 3380 375288 3392
rect 374052 3352 375288 3380
rect 374052 3340 374058 3352
rect 375282 3340 375288 3352
rect 375340 3340 375346 3392
rect 398834 3340 398840 3392
rect 398892 3380 398898 3392
rect 400122 3380 400128 3392
rect 398892 3352 400128 3380
rect 398892 3340 398898 3352
rect 400122 3340 400128 3352
rect 400180 3340 400186 3392
rect 407758 3340 407764 3392
rect 407816 3380 407822 3392
rect 409598 3380 409604 3392
rect 407816 3352 409604 3380
rect 407816 3340 407822 3352
rect 409598 3340 409604 3352
rect 409656 3340 409662 3392
rect 412606 3380 412634 3420
rect 414658 3408 414664 3460
rect 414716 3448 414722 3460
rect 416682 3448 416688 3460
rect 414716 3420 416688 3448
rect 414716 3408 414722 3420
rect 416682 3408 416688 3420
rect 416740 3408 416746 3460
rect 423692 3448 423720 3488
rect 423766 3476 423772 3528
rect 423824 3516 423830 3528
rect 424962 3516 424968 3528
rect 423824 3488 424968 3516
rect 423824 3476 423830 3488
rect 424962 3476 424968 3488
rect 425020 3476 425026 3528
rect 425790 3476 425796 3528
rect 425848 3516 425854 3528
rect 427262 3516 427268 3528
rect 425848 3488 427268 3516
rect 425848 3476 425854 3488
rect 427262 3476 427268 3488
rect 427320 3476 427326 3528
rect 431926 3516 431954 3556
rect 448514 3544 448520 3596
rect 448572 3584 448578 3596
rect 449802 3584 449808 3596
rect 448572 3556 449808 3584
rect 448572 3544 448578 3556
rect 449802 3544 449808 3556
rect 449860 3544 449866 3596
rect 449912 3584 449940 3624
rect 450538 3612 450544 3664
rect 450596 3652 450602 3664
rect 494698 3652 494704 3664
rect 450596 3624 494704 3652
rect 450596 3612 450602 3624
rect 494698 3612 494704 3624
rect 494756 3612 494762 3664
rect 519630 3612 519636 3664
rect 519688 3652 519694 3664
rect 531314 3652 531320 3664
rect 519688 3624 531320 3652
rect 519688 3612 519694 3624
rect 531314 3612 531320 3624
rect 531372 3612 531378 3664
rect 533338 3612 533344 3664
rect 533396 3652 533402 3664
rect 553762 3652 553768 3664
rect 533396 3624 553768 3652
rect 533396 3612 533402 3624
rect 553762 3612 553768 3624
rect 553820 3612 553826 3664
rect 487614 3584 487620 3596
rect 449912 3556 487620 3584
rect 487614 3544 487620 3556
rect 487672 3544 487678 3596
rect 512638 3544 512644 3596
rect 512696 3584 512702 3596
rect 527818 3584 527824 3596
rect 512696 3556 527824 3584
rect 512696 3544 512702 3556
rect 527818 3544 527824 3556
rect 527876 3544 527882 3596
rect 530578 3544 530584 3596
rect 530636 3584 530642 3596
rect 550266 3584 550272 3596
rect 530636 3556 550272 3584
rect 530636 3544 530642 3556
rect 550266 3544 550272 3556
rect 550324 3544 550330 3596
rect 551278 3544 551284 3596
rect 551336 3584 551342 3596
rect 571518 3584 571524 3596
rect 551336 3556 571524 3584
rect 551336 3544 551342 3556
rect 571518 3544 571524 3556
rect 571576 3544 571582 3596
rect 431926 3488 473216 3516
rect 426158 3448 426164 3460
rect 423692 3420 426164 3448
rect 426158 3408 426164 3420
rect 426216 3408 426222 3460
rect 432598 3408 432604 3460
rect 432656 3448 432662 3460
rect 434438 3448 434444 3460
rect 432656 3420 434444 3448
rect 432656 3408 432662 3420
rect 434438 3408 434444 3420
rect 434496 3408 434502 3460
rect 436830 3408 436836 3460
rect 436888 3448 436894 3460
rect 436888 3420 470594 3448
rect 436888 3408 436894 3420
rect 429654 3380 429660 3392
rect 412606 3352 429660 3380
rect 429654 3340 429660 3352
rect 429712 3340 429718 3392
rect 115198 3312 115204 3324
rect 98748 3284 115204 3312
rect 115198 3272 115204 3284
rect 115256 3272 115262 3324
rect 135162 3272 135168 3324
rect 135220 3312 135226 3324
rect 294874 3312 294880 3324
rect 135220 3284 294880 3312
rect 135220 3272 135226 3284
rect 294874 3272 294880 3284
rect 294932 3272 294938 3324
rect 299474 3272 299480 3324
rect 299532 3312 299538 3324
rect 300762 3312 300768 3324
rect 299532 3284 300768 3312
rect 299532 3272 299538 3284
rect 300762 3272 300768 3284
rect 300820 3272 300826 3324
rect 347130 3272 347136 3324
rect 347188 3312 347194 3324
rect 350442 3312 350448 3324
rect 347188 3284 350448 3312
rect 347188 3272 347194 3284
rect 350442 3272 350448 3284
rect 350500 3272 350506 3324
rect 470566 3312 470594 3420
rect 473188 3380 473216 3488
rect 473354 3476 473360 3528
rect 473412 3516 473418 3528
rect 474550 3516 474556 3528
rect 473412 3488 474556 3516
rect 473412 3476 473418 3488
rect 474550 3476 474556 3488
rect 474608 3476 474614 3528
rect 481634 3476 481640 3528
rect 481692 3516 481698 3528
rect 482830 3516 482836 3528
rect 481692 3488 482836 3516
rect 481692 3476 481698 3488
rect 482830 3476 482836 3488
rect 482888 3476 482894 3528
rect 483658 3476 483664 3528
rect 483716 3516 483722 3528
rect 524230 3516 524236 3528
rect 483716 3488 524236 3516
rect 483716 3476 483722 3488
rect 524230 3476 524236 3488
rect 524288 3476 524294 3528
rect 526438 3476 526444 3528
rect 526496 3516 526502 3528
rect 534902 3516 534908 3528
rect 526496 3488 534908 3516
rect 526496 3476 526502 3488
rect 534902 3476 534908 3488
rect 534960 3476 534966 3528
rect 544378 3476 544384 3528
rect 544436 3516 544442 3528
rect 568022 3516 568028 3528
rect 544436 3488 568028 3516
rect 544436 3476 544442 3488
rect 568022 3476 568028 3488
rect 568080 3476 568086 3528
rect 572714 3476 572720 3528
rect 572772 3516 572778 3528
rect 573910 3516 573916 3528
rect 572772 3488 573916 3516
rect 572772 3476 572778 3488
rect 573910 3476 573916 3488
rect 573968 3476 573974 3528
rect 580994 3448 581000 3460
rect 480226 3420 581000 3448
rect 475746 3380 475752 3392
rect 473188 3352 475752 3380
rect 475746 3340 475752 3352
rect 475804 3340 475810 3392
rect 480226 3312 480254 3420
rect 580994 3408 581000 3420
rect 581052 3408 581058 3460
rect 547874 3340 547880 3392
rect 547932 3380 547938 3392
rect 549070 3380 549076 3392
rect 547932 3352 549076 3380
rect 547932 3340 547938 3352
rect 549070 3340 549076 3352
rect 549128 3340 549134 3392
rect 470566 3284 480254 3312
rect 55950 3204 55956 3256
rect 56008 3244 56014 3256
rect 69658 3244 69664 3256
rect 56008 3216 69664 3244
rect 56008 3204 56014 3216
rect 69658 3204 69664 3216
rect 69716 3204 69722 3256
rect 89530 3204 89536 3256
rect 89588 3244 89594 3256
rect 112806 3244 112812 3256
rect 89588 3216 112812 3244
rect 89588 3204 89594 3216
rect 112806 3204 112812 3216
rect 112864 3204 112870 3256
rect 112990 3204 112996 3256
rect 113048 3244 113054 3256
rect 206186 3244 206192 3256
rect 113048 3216 206192 3244
rect 113048 3204 113054 3216
rect 206186 3204 206192 3216
rect 206244 3204 206250 3256
rect 218698 3204 218704 3256
rect 218756 3244 218762 3256
rect 376478 3244 376484 3256
rect 218756 3216 376484 3244
rect 218756 3204 218762 3216
rect 376478 3204 376484 3216
rect 376536 3204 376542 3256
rect 72510 3176 72516 3188
rect 55968 3148 72516 3176
rect 55968 3120 55996 3148
rect 72510 3136 72516 3148
rect 72568 3136 72574 3188
rect 77386 3136 77392 3188
rect 77444 3176 77450 3188
rect 79502 3176 79508 3188
rect 77444 3148 79508 3176
rect 77444 3136 77450 3148
rect 79502 3136 79508 3148
rect 79560 3136 79566 3188
rect 88242 3136 88248 3188
rect 88300 3176 88306 3188
rect 109310 3176 109316 3188
rect 88300 3148 109316 3176
rect 88300 3136 88306 3148
rect 109310 3136 109316 3148
rect 109368 3136 109374 3188
rect 109420 3148 113174 3176
rect 36044 3080 55904 3108
rect 36044 3068 36050 3080
rect 55950 3068 55956 3120
rect 56008 3068 56014 3120
rect 56134 3068 56140 3120
rect 56192 3108 56198 3120
rect 72970 3108 72976 3120
rect 56192 3080 72976 3108
rect 56192 3068 56198 3080
rect 72970 3068 72976 3080
rect 73028 3068 73034 3120
rect 86678 3068 86684 3120
rect 86736 3108 86742 3120
rect 105722 3108 105728 3120
rect 86736 3080 105728 3108
rect 86736 3068 86742 3080
rect 105722 3068 105728 3080
rect 105780 3068 105786 3120
rect 106182 3068 106188 3120
rect 106240 3108 106246 3120
rect 109420 3108 109448 3148
rect 106240 3080 109448 3108
rect 113146 3108 113174 3148
rect 126330 3136 126336 3188
rect 126388 3176 126394 3188
rect 129366 3176 129372 3188
rect 126388 3148 129372 3176
rect 126388 3136 126394 3148
rect 129366 3136 129372 3148
rect 129424 3136 129430 3188
rect 132402 3136 132408 3188
rect 132460 3176 132466 3188
rect 283098 3176 283104 3188
rect 132460 3148 283104 3176
rect 132460 3136 132466 3148
rect 283098 3136 283104 3148
rect 283156 3136 283162 3188
rect 179046 3108 179052 3120
rect 113146 3080 179052 3108
rect 106240 3068 106246 3080
rect 179046 3068 179052 3080
rect 179104 3068 179110 3120
rect 193214 3068 193220 3120
rect 193272 3108 193278 3120
rect 194410 3108 194416 3120
rect 193272 3080 194416 3108
rect 193272 3068 193278 3080
rect 194410 3068 194416 3080
rect 194468 3068 194474 3120
rect 201402 3068 201408 3120
rect 201460 3108 201466 3120
rect 207382 3108 207388 3120
rect 201460 3080 207388 3108
rect 201460 3068 201466 3080
rect 207382 3068 207388 3080
rect 207440 3068 207446 3120
rect 221642 3068 221648 3120
rect 221700 3108 221706 3120
rect 371694 3108 371700 3120
rect 221700 3080 371700 3108
rect 221700 3068 221706 3080
rect 371694 3068 371700 3080
rect 371752 3068 371758 3120
rect 24210 3000 24216 3052
rect 24268 3040 24274 3052
rect 24762 3040 24768 3052
rect 24268 3012 24768 3040
rect 24268 3000 24274 3012
rect 24762 3000 24768 3012
rect 24820 3000 24826 3052
rect 57238 3000 57244 3052
rect 57296 3040 57302 3052
rect 74442 3040 74448 3052
rect 57296 3012 74448 3040
rect 57296 3000 57302 3012
rect 74442 3000 74448 3012
rect 74500 3000 74506 3052
rect 88150 3000 88156 3052
rect 88208 3040 88214 3052
rect 108114 3040 108120 3052
rect 88208 3012 108120 3040
rect 88208 3000 88214 3012
rect 108114 3000 108120 3012
rect 108172 3000 108178 3052
rect 109006 3012 113174 3040
rect 26510 2932 26516 2984
rect 26568 2972 26574 2984
rect 27522 2972 27528 2984
rect 26568 2944 27528 2972
rect 26568 2932 26574 2944
rect 27522 2932 27528 2944
rect 27580 2932 27586 2984
rect 50154 2932 50160 2984
rect 50212 2972 50218 2984
rect 55858 2972 55864 2984
rect 50212 2944 55864 2972
rect 50212 2932 50218 2944
rect 55858 2932 55864 2944
rect 55916 2932 55922 2984
rect 64506 2972 64512 2984
rect 60706 2944 64512 2972
rect 52362 2864 52368 2916
rect 52420 2904 52426 2916
rect 60706 2904 60734 2944
rect 64506 2932 64512 2944
rect 64564 2932 64570 2984
rect 86862 2932 86868 2984
rect 86920 2972 86926 2984
rect 104526 2972 104532 2984
rect 86920 2944 104532 2972
rect 86920 2932 86926 2944
rect 104526 2932 104532 2944
rect 104584 2932 104590 2984
rect 104618 2932 104624 2984
rect 104676 2972 104682 2984
rect 109006 2972 109034 3012
rect 104676 2944 109034 2972
rect 113146 2972 113174 3012
rect 219342 3000 219348 3052
rect 219400 3040 219406 3052
rect 323302 3040 323308 3052
rect 219400 3012 323308 3040
rect 219400 3000 219406 3012
rect 323302 3000 323308 3012
rect 323360 3000 323366 3052
rect 417510 3000 417516 3052
rect 417568 3040 417574 3052
rect 420178 3040 420184 3052
rect 417568 3012 420184 3040
rect 417568 3000 417574 3012
rect 420178 3000 420184 3012
rect 420236 3000 420242 3052
rect 114002 2972 114008 2984
rect 113146 2944 114008 2972
rect 104676 2932 104682 2944
rect 114002 2932 114008 2944
rect 114060 2932 114066 2984
rect 221458 2932 221464 2984
rect 221516 2972 221522 2984
rect 305546 2972 305552 2984
rect 221516 2944 305552 2972
rect 221516 2932 221522 2944
rect 305546 2932 305552 2944
rect 305604 2932 305610 2984
rect 52420 2876 60734 2904
rect 52420 2864 52426 2876
rect 86770 2864 86776 2916
rect 86828 2904 86834 2916
rect 102226 2904 102232 2916
rect 86828 2876 102232 2904
rect 86828 2864 86834 2876
rect 102226 2864 102232 2876
rect 102284 2864 102290 2916
rect 102318 2864 102324 2916
rect 102376 2904 102382 2916
rect 103606 2904 103612 2916
rect 102376 2876 103612 2904
rect 102376 2864 102382 2876
rect 103606 2864 103612 2876
rect 103664 2864 103670 2916
rect 103698 2864 103704 2916
rect 103756 2904 103762 2916
rect 110598 2904 110604 2916
rect 103756 2876 110604 2904
rect 103756 2864 103762 2876
rect 110598 2864 110604 2876
rect 110656 2864 110662 2916
rect 221550 2864 221556 2916
rect 221608 2904 221614 2916
rect 298462 2904 298468 2916
rect 221608 2876 298468 2904
rect 221608 2864 221614 2876
rect 298462 2864 298468 2876
rect 298520 2864 298526 2916
rect 55214 2796 55220 2848
rect 55272 2836 55278 2848
rect 59446 2836 59452 2848
rect 55272 2808 59452 2836
rect 55272 2796 55278 2808
rect 59446 2796 59452 2808
rect 59504 2796 59510 2848
rect 82722 2796 82728 2848
rect 82780 2836 82786 2848
rect 86862 2836 86868 2848
rect 82780 2808 86868 2836
rect 82780 2796 82786 2808
rect 86862 2796 86868 2808
rect 86920 2796 86926 2848
rect 87598 2796 87604 2848
rect 87656 2836 87662 2848
rect 98638 2836 98644 2848
rect 87656 2808 98644 2836
rect 87656 2796 87662 2808
rect 98638 2796 98644 2808
rect 98696 2796 98702 2848
rect 99374 2836 99380 2848
rect 98748 2808 99380 2836
rect 98454 2728 98460 2780
rect 98512 2768 98518 2780
rect 98748 2768 98776 2808
rect 99374 2796 99380 2808
rect 99432 2796 99438 2848
rect 103882 2796 103888 2848
rect 103940 2836 103946 2848
rect 110138 2836 110144 2848
rect 103940 2808 110144 2836
rect 103940 2796 103946 2808
rect 110138 2796 110144 2808
rect 110196 2796 110202 2848
rect 242894 2796 242900 2848
rect 242952 2836 242958 2848
rect 244090 2836 244096 2848
rect 242952 2808 244096 2836
rect 242952 2796 242958 2808
rect 244090 2796 244096 2808
rect 244148 2796 244154 2848
rect 270402 2796 270408 2848
rect 270460 2836 270466 2848
rect 272426 2836 272432 2848
rect 270460 2808 272432 2836
rect 270460 2796 270466 2808
rect 272426 2796 272432 2808
rect 272484 2796 272490 2848
rect 98512 2740 98776 2768
rect 98512 2728 98518 2740
rect 154298 2116 154304 2168
rect 154356 2156 154362 2168
rect 369394 2156 369400 2168
rect 154356 2128 369400 2156
rect 154356 2116 154362 2128
rect 369394 2116 369400 2128
rect 369452 2116 369458 2168
rect 154390 2048 154396 2100
rect 154448 2088 154454 2100
rect 372890 2088 372896 2100
rect 154448 2060 372896 2088
rect 154448 2048 154454 2060
rect 372890 2048 372896 2060
rect 372948 2048 372954 2100
rect 99190 960 99196 1012
rect 99248 1000 99254 1012
rect 99834 1000 99840 1012
rect 99248 972 99840 1000
rect 99248 960 99254 972
rect 99834 960 99840 972
rect 99892 960 99898 1012
rect 51350 688 51356 740
rect 51408 728 51414 740
rect 56134 728 56140 740
rect 51408 700 56140 728
rect 51408 688 51414 700
rect 56134 688 56140 700
rect 56192 688 56198 740
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 215944 700680 215996 700732
rect 235172 700680 235224 700732
rect 209044 700612 209096 700664
rect 267648 700612 267700 700664
rect 206376 700544 206428 700596
rect 283840 700544 283892 700596
rect 385684 700544 385736 700596
rect 397460 700544 397512 700596
rect 399484 700544 399536 700596
rect 478512 700544 478564 700596
rect 206284 700476 206336 700528
rect 300124 700476 300176 700528
rect 382924 700476 382976 700528
rect 462320 700476 462372 700528
rect 204904 700408 204956 700460
rect 332508 700408 332560 700460
rect 370504 700408 370556 700460
rect 494796 700408 494848 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 170312 700340 170364 700392
rect 196532 700340 196584 700392
rect 213184 700340 213236 700392
rect 348792 700340 348844 700392
rect 381544 700340 381596 700392
rect 527180 700340 527232 700392
rect 24308 700272 24360 700324
rect 33784 700272 33836 700324
rect 58900 700272 58952 700324
rect 72976 700272 73028 700324
rect 154120 700272 154172 700324
rect 196624 700272 196676 700324
rect 198004 700272 198056 700324
rect 364984 700272 365036 700324
rect 367744 700272 367796 700324
rect 559656 700272 559708 700324
rect 88340 699660 88392 699712
rect 89168 699660 89220 699712
rect 104900 699660 104952 699712
rect 105452 699660 105504 699712
rect 210424 699660 210476 699712
rect 218980 699660 219032 699712
rect 134156 698572 134208 698624
rect 137836 698572 137888 698624
rect 128912 696872 128964 696924
rect 134156 696940 134208 696992
rect 378784 696940 378836 696992
rect 580172 696940 580224 696992
rect 126520 693744 126572 693796
rect 128912 693744 128964 693796
rect 124588 690140 124640 690192
rect 126520 690140 126572 690192
rect 121460 688644 121512 688696
rect 124588 688644 124640 688696
rect 114560 684360 114612 684412
rect 121460 684360 121512 684412
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 396724 683136 396776 683188
rect 580172 683136 580224 683188
rect 106280 681640 106332 681692
rect 114560 681708 114612 681760
rect 104256 674704 104308 674756
rect 106188 674704 106240 674756
rect 3516 670692 3568 670744
rect 35164 670692 35216 670744
rect 363604 670692 363656 670744
rect 580172 670692 580224 670744
rect 102784 667360 102836 667412
rect 104256 667360 104308 667412
rect 100760 662396 100812 662448
rect 102784 662396 102836 662448
rect 96528 659608 96580 659660
rect 100760 659676 100812 659728
rect 94504 657976 94556 658028
rect 96528 657976 96580 658028
rect 3424 656888 3476 656940
rect 21364 656888 21416 656940
rect 92480 650088 92532 650140
rect 94504 650088 94556 650140
rect 77208 647844 77260 647896
rect 92480 647844 92532 647896
rect 74540 645872 74592 645924
rect 77208 645872 77260 645924
rect 377404 643084 377456 643136
rect 580172 643084 580224 643136
rect 74540 638936 74592 638988
rect 71780 638868 71832 638920
rect 69020 636148 69072 636200
rect 71780 636216 71832 636268
rect 3424 632068 3476 632120
rect 11704 632068 11756 632120
rect 65524 632000 65576 632052
rect 69020 632068 69072 632120
rect 395344 630640 395396 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 36544 618264 36596 618316
rect 360844 616836 360896 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 22744 605820 22796 605872
rect 64144 604460 64196 604512
rect 65524 604460 65576 604512
rect 558184 590656 558236 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 14464 579640 14516 579692
rect 393964 576852 394016 576904
rect 580172 576852 580224 576904
rect 62764 572704 62816 572756
rect 64144 572704 64196 572756
rect 3424 565836 3476 565888
rect 39304 565836 39356 565888
rect 358084 563048 358136 563100
rect 579804 563048 579856 563100
rect 61384 561008 61436 561060
rect 62764 561008 62816 561060
rect 3424 553392 3476 553444
rect 25504 553392 25556 553444
rect 60004 553392 60056 553444
rect 61384 553392 61436 553444
rect 376024 536800 376076 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 15844 527144 15896 527196
rect 392584 524424 392636 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 43444 514768 43496 514820
rect 213368 510620 213420 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 29644 500964 29696 501016
rect 374644 484372 374696 484424
rect 580172 484372 580224 484424
rect 3424 474716 3476 474768
rect 17224 474716 17276 474768
rect 389824 470568 389876 470620
rect 579988 470568 580040 470620
rect 3240 462340 3292 462392
rect 47584 462340 47636 462392
rect 425704 456764 425756 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 32404 448536 32456 448588
rect 209228 430584 209280 430636
rect 216680 430584 216732 430636
rect 388444 430584 388496 430636
rect 580172 430584 580224 430636
rect 3424 422288 3476 422340
rect 18604 422288 18656 422340
rect 214564 408348 214616 408400
rect 216680 408348 216732 408400
rect 371884 404336 371936 404388
rect 580172 404336 580224 404388
rect 218612 400052 218664 400104
rect 218152 399984 218204 400036
rect 226340 399984 226392 400036
rect 226708 399984 226760 400036
rect 218244 399916 218296 399968
rect 226524 399916 226576 399968
rect 217600 399848 217652 399900
rect 231860 399848 231912 399900
rect 58900 399780 58952 399832
rect 121460 399780 121512 399832
rect 177948 399780 178000 399832
rect 209228 399780 209280 399832
rect 217692 399780 217744 399832
rect 232136 399780 232188 399832
rect 111708 399712 111760 399764
rect 204904 399712 204956 399764
rect 217416 399712 217468 399764
rect 233240 399712 233292 399764
rect 57060 399644 57112 399696
rect 230756 399644 230808 399696
rect 57244 399576 57296 399628
rect 232044 399576 232096 399628
rect 57152 399508 57204 399560
rect 231952 399508 232004 399560
rect 244924 399508 244976 399560
rect 359004 399508 359056 399560
rect 57336 399440 57388 399492
rect 232228 399440 232280 399492
rect 242256 399440 242308 399492
rect 359096 399440 359148 399492
rect 218428 399372 218480 399424
rect 226432 399372 226484 399424
rect 60004 398828 60056 398880
rect 62028 398828 62080 398880
rect 59360 398760 59412 398812
rect 214564 398760 214616 398812
rect 219532 398692 219584 398744
rect 224960 398692 225012 398744
rect 219624 398556 219676 398608
rect 225236 398556 225288 398608
rect 219900 398488 219952 398540
rect 226616 398488 226668 398540
rect 121368 398216 121420 398268
rect 196624 398216 196676 398268
rect 115848 398148 115900 398200
rect 206376 398148 206428 398200
rect 218060 398148 218112 398200
rect 225144 398216 225196 398268
rect 219716 398148 219768 398200
rect 225052 398148 225104 398200
rect 57888 398080 57940 398132
rect 165620 398080 165672 398132
rect 217508 398080 217560 398132
rect 232320 398080 232372 398132
rect 3516 397468 3568 397520
rect 140780 397468 140832 397520
rect 216588 397332 216640 397384
rect 275284 397332 275336 397384
rect 85488 397264 85540 397316
rect 230572 397264 230624 397316
rect 304264 397264 304316 397316
rect 308588 397264 308640 397316
rect 62948 397196 63000 397248
rect 239220 397196 239272 397248
rect 79600 397128 79652 397180
rect 230664 397128 230716 397180
rect 253296 397128 253348 397180
rect 259460 397128 259512 397180
rect 89352 397060 89404 397112
rect 94504 397060 94556 397112
rect 183468 397060 183520 397112
rect 229284 397060 229336 397112
rect 62764 396992 62816 397044
rect 113824 396992 113876 397044
rect 206928 396992 206980 397044
rect 268660 396992 268712 397044
rect 61476 396924 61528 396976
rect 109132 396924 109184 396976
rect 188344 396924 188396 396976
rect 250076 396924 250128 396976
rect 82360 396856 82412 396908
rect 162124 396856 162176 396908
rect 173164 396856 173216 396908
rect 236184 396856 236236 396908
rect 78312 396788 78364 396840
rect 168380 396788 168432 396840
rect 186964 396788 187016 396840
rect 252744 396788 252796 396840
rect 113364 396720 113416 396772
rect 230848 396720 230900 396772
rect 250444 396720 250496 396772
rect 256884 396720 256936 396772
rect 262864 396720 262916 396772
rect 265164 396720 265216 396772
rect 268476 396720 268528 396772
rect 269396 396720 269448 396772
rect 282184 396720 282236 396772
rect 283748 396720 283800 396772
rect 291844 396720 291896 396772
rect 292672 396720 292724 396772
rect 112352 396652 112404 396704
rect 230940 396652 230992 396704
rect 242164 396652 242216 396704
rect 244556 396652 244608 396704
rect 249064 396652 249116 396704
rect 251364 396652 251416 396704
rect 251916 396652 251968 396704
rect 254124 396652 254176 396704
rect 268384 396652 268436 396704
rect 273628 396652 273680 396704
rect 284944 396652 284996 396704
rect 285956 396652 286008 396704
rect 58624 396584 58676 396636
rect 95884 396584 95936 396636
rect 106924 396584 106976 396636
rect 230480 396584 230532 396636
rect 61384 396516 61436 396568
rect 98092 396516 98144 396568
rect 104808 396516 104860 396568
rect 229376 396516 229428 396568
rect 95056 396448 95108 396500
rect 229100 396448 229152 396500
rect 246304 396448 246356 396500
rect 263600 396448 263652 396500
rect 90088 396380 90140 396432
rect 227720 396380 227772 396432
rect 260104 396380 260156 396432
rect 325884 396380 325936 396432
rect 60004 396312 60056 396364
rect 76196 396312 76248 396364
rect 91468 396312 91520 396364
rect 229192 396312 229244 396364
rect 235264 396312 235316 396364
rect 272340 396312 272392 396364
rect 93492 396244 93544 396296
rect 231032 396244 231084 396296
rect 233976 396244 234028 396296
rect 247684 396244 247736 396296
rect 253204 396244 253256 396296
rect 261944 396244 261996 396296
rect 269764 396244 269816 396296
rect 315764 396244 315816 396296
rect 58900 396176 58952 396228
rect 83004 396176 83056 396228
rect 222844 396176 222896 396228
rect 277676 396176 277728 396228
rect 59912 396108 59964 396160
rect 80428 396108 80480 396160
rect 106096 396108 106148 396160
rect 115204 396108 115256 396160
rect 237472 396108 237524 396160
rect 248604 396108 248656 396160
rect 255964 396108 256016 396160
rect 260932 396108 260984 396160
rect 316684 396108 316736 396160
rect 342628 396108 342680 396160
rect 102784 396040 102836 396092
rect 106924 396040 106976 396092
rect 108856 396040 108908 396092
rect 119344 396040 119396 396092
rect 163872 395972 163924 396024
rect 219440 395972 219492 396024
rect 251824 395972 251876 396024
rect 256148 395972 256200 396024
rect 118608 395904 118660 395956
rect 189080 395904 189132 395956
rect 113640 395836 113692 395888
rect 184940 395836 184992 395888
rect 195888 395836 195940 395888
rect 262312 395836 262364 395888
rect 154120 395768 154172 395820
rect 227996 395768 228048 395820
rect 171048 395700 171100 395752
rect 250352 395700 250404 395752
rect 184848 395632 184900 395684
rect 268292 395632 268344 395684
rect 136456 395564 136508 395616
rect 227812 395564 227864 395616
rect 118240 395496 118292 395548
rect 224868 395496 224920 395548
rect 233884 395496 233936 395548
rect 247960 395496 248012 395548
rect 61568 395428 61620 395480
rect 278872 395428 278924 395480
rect 56508 395360 56560 395412
rect 290188 395360 290240 395412
rect 54576 395292 54628 395344
rect 298468 395292 298520 395344
rect 62120 394680 62172 394732
rect 66260 394612 66312 394664
rect 238024 394000 238076 394052
rect 251180 394000 251232 394052
rect 177856 393932 177908 393984
rect 237472 393932 237524 393984
rect 240784 392640 240836 392692
rect 258172 392640 258224 392692
rect 193128 392572 193180 392624
rect 253296 392572 253348 392624
rect 258724 392572 258776 392624
rect 277492 392572 277544 392624
rect 66260 389172 66312 389224
rect 68284 389172 68336 389224
rect 84108 378156 84160 378208
rect 580172 378156 580224 378208
rect 68284 378088 68336 378140
rect 69664 378088 69716 378140
rect 43444 373396 43496 373448
rect 136640 373396 136692 373448
rect 39304 373328 39356 373380
rect 133880 373328 133932 373380
rect 3424 373260 3476 373312
rect 142160 373260 142212 373312
rect 195796 373260 195848 373312
rect 287060 373260 287112 373312
rect 69664 372852 69716 372904
rect 70400 372852 70452 372904
rect 3424 371220 3476 371272
rect 143540 371220 143592 371272
rect 70400 369792 70452 369844
rect 75184 369792 75236 369844
rect 85488 364352 85540 364404
rect 579620 364352 579672 364404
rect 75184 358708 75236 358760
rect 76656 358708 76708 358760
rect 3148 357416 3200 357468
rect 144920 357416 144972 357468
rect 76656 357348 76708 357400
rect 78036 357348 78088 357400
rect 56324 356668 56376 356720
rect 145012 356668 145064 356720
rect 78036 353268 78088 353320
rect 80704 353268 80756 353320
rect 82728 351908 82780 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 143632 345040 143684 345092
rect 80704 335996 80756 336048
rect 84200 335996 84252 336048
rect 84200 329740 84252 329792
rect 86224 329740 86276 329792
rect 86224 324572 86276 324624
rect 87972 324572 88024 324624
rect 81348 324300 81400 324352
rect 580172 324300 580224 324352
rect 87972 322940 88024 322992
rect 91744 322872 91796 322924
rect 3424 318792 3476 318844
rect 146300 318792 146352 318844
rect 91744 314236 91796 314288
rect 94596 314236 94648 314288
rect 82636 311856 82688 311908
rect 579988 311856 580040 311908
rect 113088 305600 113140 305652
rect 213184 305600 213236 305652
rect 3240 304988 3292 305040
rect 147680 304988 147732 305040
rect 79968 298120 80020 298172
rect 580172 298120 580224 298172
rect 94596 295332 94648 295384
rect 97264 295332 97316 295384
rect 3424 292544 3476 292596
rect 146392 292544 146444 292596
rect 97264 282888 97316 282940
rect 99472 282820 99524 282872
rect 99472 278672 99524 278724
rect 101496 278672 101548 278724
rect 101496 275204 101548 275256
rect 102140 275204 102192 275256
rect 78588 271872 78640 271924
rect 580172 271872 580224 271924
rect 102140 269084 102192 269136
rect 104164 269084 104216 269136
rect 77208 266976 77260 267028
rect 168472 266976 168524 267028
rect 3056 266364 3108 266416
rect 149060 266364 149112 266416
rect 106924 266296 106976 266348
rect 195980 266296 196032 266348
rect 101956 266228 102008 266280
rect 193220 266228 193272 266280
rect 107476 266160 107528 266212
rect 202880 266160 202932 266212
rect 92296 266092 92348 266144
rect 225880 266092 225932 266144
rect 86868 266024 86920 266076
rect 225604 266024 225656 266076
rect 85396 265956 85448 266008
rect 231124 265956 231176 266008
rect 88248 265888 88300 265940
rect 175280 265888 175332 265940
rect 182088 265888 182140 265940
rect 358912 265888 358964 265940
rect 53196 265820 53248 265872
rect 259552 265820 259604 265872
rect 54300 265752 54352 265804
rect 313280 265752 313332 265804
rect 54208 265684 54260 265736
rect 317420 265684 317472 265736
rect 88248 265616 88300 265668
rect 580264 265616 580316 265668
rect 115204 265548 115256 265600
rect 200120 265548 200172 265600
rect 94504 265480 94556 265532
rect 178040 265480 178092 265532
rect 187608 265480 187660 265532
rect 251916 265480 251968 265532
rect 184756 264936 184808 264988
rect 186964 264936 187016 264988
rect 36544 264868 36596 264920
rect 131120 264868 131172 264920
rect 133788 264868 133840 264920
rect 198096 264868 198148 264920
rect 209596 264868 209648 264920
rect 268476 264868 268528 264920
rect 55864 264800 55916 264852
rect 155960 264800 156012 264852
rect 173808 264800 173860 264852
rect 252560 264800 252612 264852
rect 119988 264732 120040 264784
rect 223672 264732 223724 264784
rect 8208 264664 8260 264716
rect 124220 264664 124272 264716
rect 131028 264664 131080 264716
rect 228548 264664 228600 264716
rect 111524 264596 111576 264648
rect 229468 264596 229520 264648
rect 100668 264528 100720 264580
rect 231308 264528 231360 264580
rect 90916 264460 90968 264512
rect 227904 264460 227956 264512
rect 59544 264392 59596 264444
rect 273352 264392 273404 264444
rect 54392 264324 54444 264376
rect 276112 264324 276164 264376
rect 107568 264256 107620 264308
rect 399484 264256 399536 264308
rect 104808 264188 104860 264240
rect 542360 264188 542412 264240
rect 35164 264120 35216 264172
rect 128360 264120 128412 264172
rect 139308 264120 139360 264172
rect 201592 264120 201644 264172
rect 223488 264120 223540 264172
rect 260104 264120 260156 264172
rect 33784 264052 33836 264104
rect 125600 264052 125652 264104
rect 161388 264052 161440 264104
rect 216404 264052 216456 264104
rect 47584 263984 47636 264036
rect 139400 263984 139452 264036
rect 201408 263984 201460 264036
rect 246304 263984 246356 264036
rect 119344 263916 119396 263968
rect 205640 263916 205692 263968
rect 119988 263848 120040 263900
rect 196532 263848 196584 263900
rect 89536 263780 89588 263832
rect 165712 263780 165764 263832
rect 99288 263508 99340 263560
rect 228364 263508 228416 263560
rect 231400 263508 231452 263560
rect 310520 263508 310572 263560
rect 108948 263440 109000 263492
rect 385684 263440 385736 263492
rect 106096 263372 106148 263424
rect 382924 263372 382976 263424
rect 103428 263304 103480 263356
rect 381544 263304 381596 263356
rect 97816 263236 97868 263288
rect 377404 263236 377456 263288
rect 101956 263168 102008 263220
rect 396724 263168 396776 263220
rect 99288 263100 99340 263152
rect 395344 263100 395396 263152
rect 91008 263032 91060 263084
rect 389824 263032 389876 263084
rect 93768 262964 93820 263016
rect 392584 262964 392636 263016
rect 86868 262896 86920 262948
rect 388444 262896 388496 262948
rect 110328 262828 110380 262880
rect 412640 262828 412692 262880
rect 56048 262760 56100 262812
rect 115940 262760 115992 262812
rect 117228 262760 117280 262812
rect 225512 262760 225564 262812
rect 234252 262760 234304 262812
rect 266452 262760 266504 262812
rect 22744 262692 22796 262744
rect 129740 262692 129792 262744
rect 162124 262692 162176 262744
rect 173900 262692 173952 262744
rect 181996 262692 182048 262744
rect 188344 262692 188396 262744
rect 198556 262692 198608 262744
rect 291844 262692 291896 262744
rect 25504 262624 25556 262676
rect 132500 262624 132552 262676
rect 151728 262624 151780 262676
rect 212540 262624 212592 262676
rect 21364 262556 21416 262608
rect 126980 262556 127032 262608
rect 32404 262488 32456 262540
rect 138020 262488 138072 262540
rect 117228 262420 117280 262472
rect 201500 262420 201552 262472
rect 4804 262148 4856 262200
rect 127072 262148 127124 262200
rect 144828 262148 144880 262200
rect 202972 262148 203024 262200
rect 211068 262148 211120 262200
rect 304264 262148 304316 262200
rect 97908 262080 97960 262132
rect 229652 262080 229704 262132
rect 235448 262080 235500 262132
rect 280160 262080 280212 262132
rect 59452 262012 59504 262064
rect 265072 262012 265124 262064
rect 101864 261944 101916 261996
rect 367744 261944 367796 261996
rect 104716 261876 104768 261928
rect 370504 261876 370556 261928
rect 100668 261808 100720 261860
rect 378784 261808 378836 261860
rect 92388 261740 92440 261792
rect 376024 261740 376076 261792
rect 89628 261672 89680 261724
rect 374644 261672 374696 261724
rect 96436 261604 96488 261656
rect 393964 261604 394016 261656
rect 108856 261536 108908 261588
rect 429200 261536 429252 261588
rect 95148 261468 95200 261520
rect 558184 261468 558236 261520
rect 18604 261400 18656 261452
rect 140872 261400 140924 261452
rect 193036 261400 193088 261452
rect 284944 261400 284996 261452
rect 17224 261332 17276 261384
rect 138112 261332 138164 261384
rect 190368 261332 190420 261384
rect 282184 261332 282236 261384
rect 14464 261264 14516 261316
rect 132592 261264 132644 261316
rect 142068 261264 142120 261316
rect 228640 261264 228692 261316
rect 232504 261264 232556 261316
rect 273444 261264 273496 261316
rect 11704 261196 11756 261248
rect 129832 261196 129884 261248
rect 148968 261196 149020 261248
rect 211252 261196 211304 261248
rect 238208 261196 238260 261248
rect 258080 261196 258132 261248
rect 29644 261128 29696 261180
rect 135260 261128 135312 261180
rect 200856 261128 200908 261180
rect 224776 261128 224828 261180
rect 117136 261060 117188 261112
rect 215944 261060 215996 261112
rect 118608 260992 118660 261044
rect 210424 260992 210476 261044
rect 111524 260924 111576 260976
rect 198004 260924 198056 260976
rect 41328 260856 41380 260908
rect 124312 260856 124364 260908
rect 104164 260788 104216 260840
rect 106648 260788 106700 260840
rect 172428 260788 172480 260840
rect 173164 260788 173216 260840
rect 199660 260788 199712 260840
rect 229560 260788 229612 260840
rect 114468 260720 114520 260772
rect 206284 260720 206336 260772
rect 56140 260652 56192 260704
rect 103520 260652 103572 260704
rect 114376 260652 114428 260704
rect 209044 260652 209096 260704
rect 15844 260584 15896 260636
rect 135352 260584 135404 260636
rect 208308 260584 208360 260636
rect 305000 260584 305052 260636
rect 90916 260516 90968 260568
rect 213368 260516 213420 260568
rect 213644 260516 213696 260568
rect 226892 260516 226944 260568
rect 238300 260516 238352 260568
rect 270592 260516 270644 260568
rect 102048 260448 102100 260500
rect 228456 260448 228508 260500
rect 234160 260448 234212 260500
rect 295340 260448 295392 260500
rect 99196 260380 99248 260432
rect 363604 260380 363656 260432
rect 93676 260312 93728 260364
rect 358084 260312 358136 260364
rect 96344 260244 96396 260296
rect 360844 260244 360896 260296
rect 85396 260176 85448 260228
rect 371884 260176 371936 260228
rect 88156 260108 88208 260160
rect 425704 260108 425756 260160
rect 260748 245556 260800 245608
rect 580172 245556 580224 245608
rect 55772 229100 55824 229152
rect 59820 229100 59872 229152
rect 57428 218016 57480 218068
rect 58532 218016 58584 218068
rect 3056 215228 3108 215280
rect 11704 215228 11756 215280
rect 54208 213868 54260 213920
rect 57520 213868 57572 213920
rect 54300 197276 54352 197328
rect 57520 197276 57572 197328
rect 54668 194488 54720 194540
rect 57520 194488 57572 194540
rect 271144 193128 271196 193180
rect 580172 193128 580224 193180
rect 53288 191768 53340 191820
rect 57520 191768 57572 191820
rect 3332 188844 3384 188896
rect 7564 188844 7616 188896
rect 54760 182112 54812 182164
rect 57520 182112 57572 182164
rect 53380 177964 53432 178016
rect 57520 177964 57572 178016
rect 54576 175176 54628 175228
rect 57520 175176 57572 175228
rect 3056 164160 3108 164212
rect 14464 164160 14516 164212
rect 53472 160012 53524 160064
rect 57428 160012 57480 160064
rect 53196 155864 53248 155916
rect 57520 155864 57572 155916
rect 54852 153144 54904 153196
rect 57520 153144 57572 153196
rect 53564 147568 53616 147620
rect 57428 147568 57480 147620
rect 53656 143488 53708 143540
rect 57520 143488 57572 143540
rect 3056 137912 3108 137964
rect 17224 137912 17276 137964
rect 57520 136552 57572 136604
rect 59820 136552 59872 136604
rect 54392 134716 54444 134768
rect 57428 134716 57480 134768
rect 53748 131044 53800 131096
rect 57612 131044 57664 131096
rect 57704 127916 57756 127968
rect 58716 127916 58768 127968
rect 54944 118600 54996 118652
rect 57612 118600 57664 118652
rect 55036 113092 55088 113144
rect 57612 113092 57664 113144
rect 3332 111732 3384 111784
rect 15844 111732 15896 111784
rect 57704 106224 57756 106276
rect 59820 106224 59872 106276
rect 410524 100648 410576 100700
rect 580172 100648 580224 100700
rect 3240 97928 3292 97980
rect 18604 97928 18656 97980
rect 2964 85484 3016 85536
rect 32404 85484 32456 85536
rect 3332 71680 3384 71732
rect 29644 71680 29696 71732
rect 54484 71680 54536 71732
rect 57612 71680 57664 71732
rect 55128 62024 55180 62076
rect 57060 62024 57112 62076
rect 580172 59916 580224 59968
rect 222108 59848 222160 59900
rect 222568 59780 222620 59832
rect 224132 59780 224184 59832
rect 224316 59780 224368 59832
rect 224224 59712 224276 59764
rect 224776 59712 224828 59764
rect 240876 59848 240928 59900
rect 302240 59848 302292 59900
rect 263692 59780 263744 59832
rect 223580 59440 223632 59492
rect 268384 59440 268436 59492
rect 224500 59372 224552 59424
rect 276020 59372 276072 59424
rect 57796 59304 57848 59356
rect 217048 59304 217100 59356
rect 217968 59304 218020 59356
rect 229100 59304 229152 59356
rect 220912 59236 220964 59288
rect 229376 59236 229428 59288
rect 221556 59168 221608 59220
rect 230480 59168 230532 59220
rect 209872 59100 209924 59152
rect 230664 59100 230716 59152
rect 150624 59032 150676 59084
rect 151452 59032 151504 59084
rect 216772 59032 216824 59084
rect 229284 59032 229336 59084
rect 149428 58964 149480 59016
rect 150256 58964 150308 59016
rect 150716 58964 150768 59016
rect 151728 58964 151780 59016
rect 215852 58964 215904 59016
rect 229192 58964 229244 59016
rect 219164 58896 219216 58948
rect 250444 58896 250496 58948
rect 211344 58828 211396 58880
rect 240140 58828 240192 58880
rect 209228 58760 209280 58812
rect 237380 58760 237432 58812
rect 214380 58692 214432 58744
rect 227720 58692 227772 58744
rect 212264 58624 212316 58676
rect 245660 58624 245712 58676
rect 210700 58556 210752 58608
rect 230572 58556 230624 58608
rect 208952 58488 209004 58540
rect 236000 58488 236052 58540
rect 214932 58420 214984 58472
rect 262864 58420 262916 58472
rect 209504 58352 209556 58404
rect 244372 58352 244424 58404
rect 216404 58284 216456 58336
rect 342352 58284 342404 58336
rect 218520 58216 218572 58268
rect 255412 58216 255464 58268
rect 220636 58148 220688 58200
rect 253204 58148 253256 58200
rect 215576 58080 215628 58132
rect 316684 58080 316736 58132
rect 180800 58012 180852 58064
rect 181168 58012 181220 58064
rect 208676 58012 208728 58064
rect 224960 58012 225012 58064
rect 180708 57944 180760 57996
rect 181720 57944 181772 57996
rect 207756 57944 207808 57996
rect 208308 57944 208360 57996
rect 216588 57944 216640 57996
rect 39948 57876 40000 57928
rect 69940 57876 69992 57928
rect 34428 57808 34480 57860
rect 68468 57808 68520 57860
rect 30288 57740 30340 57792
rect 67548 57740 67600 57792
rect 76840 57876 76892 57928
rect 87880 57876 87932 57928
rect 95332 57876 95384 57928
rect 95424 57876 95476 57928
rect 103980 57876 104032 57928
rect 107108 57876 107160 57928
rect 75092 57808 75144 57860
rect 77392 57808 77444 57860
rect 91836 57808 91888 57860
rect 113732 57808 113784 57860
rect 118148 57808 118200 57860
rect 118608 57808 118660 57860
rect 120908 57808 120960 57860
rect 33048 57672 33100 57724
rect 68100 57672 68152 57724
rect 28908 57604 28960 57656
rect 66904 57604 66956 57656
rect 67548 57604 67600 57656
rect 73068 57672 73120 57724
rect 78312 57740 78364 57792
rect 84292 57740 84344 57792
rect 88984 57740 89036 57792
rect 92664 57740 92716 57792
rect 126244 57740 126296 57792
rect 126428 57808 126480 57860
rect 133788 57876 133840 57928
rect 139492 57876 139544 57928
rect 141792 57876 141844 57928
rect 218888 57876 218940 57928
rect 218980 57876 219032 57928
rect 220360 57876 220412 57928
rect 225328 57876 225380 57928
rect 226984 57876 227036 57928
rect 300124 57876 300176 57928
rect 128452 57740 128504 57792
rect 136272 57808 136324 57860
rect 137376 57808 137428 57860
rect 142528 57740 142580 57792
rect 27528 57536 27580 57588
rect 66628 57536 66680 57588
rect 70308 57536 70360 57588
rect 77760 57672 77812 57724
rect 84660 57672 84712 57724
rect 86316 57672 86368 57724
rect 88800 57672 88852 57724
rect 103888 57672 103940 57724
rect 113824 57672 113876 57724
rect 80704 57604 80756 57656
rect 81256 57604 81308 57656
rect 82176 57604 82228 57656
rect 82636 57604 82688 57656
rect 83096 57604 83148 57656
rect 84108 57604 84160 57656
rect 85212 57604 85264 57656
rect 86224 57604 86276 57656
rect 86408 57604 86460 57656
rect 86868 57604 86920 57656
rect 89996 57604 90048 57656
rect 90732 57604 90784 57656
rect 91468 57604 91520 57656
rect 92388 57604 92440 57656
rect 93308 57604 93360 57656
rect 127900 57604 127952 57656
rect 127992 57604 128044 57656
rect 128176 57604 128228 57656
rect 135536 57672 135588 57724
rect 216588 57740 216640 57792
rect 216680 57740 216732 57792
rect 218244 57740 218296 57792
rect 137192 57604 137244 57656
rect 75828 57536 75880 57588
rect 78956 57536 79008 57588
rect 81900 57536 81952 57588
rect 82728 57536 82780 57588
rect 85856 57536 85908 57588
rect 86776 57536 86828 57588
rect 89720 57536 89772 57588
rect 91008 57536 91060 57588
rect 94504 57536 94556 57588
rect 95148 57536 95200 57588
rect 95976 57536 96028 57588
rect 96528 57536 96580 57588
rect 97172 57536 97224 57588
rect 97724 57536 97776 57588
rect 98920 57536 98972 57588
rect 99288 57536 99340 57588
rect 104256 57536 104308 57588
rect 131856 57536 131908 57588
rect 132040 57536 132092 57588
rect 138664 57604 138716 57656
rect 142712 57604 142764 57656
rect 161848 57672 161900 57724
rect 167644 57672 167696 57724
rect 168104 57672 168156 57724
rect 169300 57672 169352 57724
rect 169668 57672 169720 57724
rect 171232 57672 171284 57724
rect 172244 57672 172296 57724
rect 172704 57672 172756 57724
rect 173808 57672 173860 57724
rect 174452 57672 174504 57724
rect 175188 57672 175240 57724
rect 175556 57672 175608 57724
rect 176568 57672 176620 57724
rect 177212 57672 177264 57724
rect 177948 57672 178000 57724
rect 178040 57672 178092 57724
rect 179328 57672 179380 57724
rect 180708 57672 180760 57724
rect 180984 57672 181036 57724
rect 181076 57672 181128 57724
rect 181720 57672 181772 57724
rect 182548 57672 182600 57724
rect 183100 57672 183152 57724
rect 183744 57672 183796 57724
rect 184756 57672 184808 57724
rect 186780 57672 186832 57724
rect 187424 57672 187476 57724
rect 187700 57672 187752 57724
rect 188896 57672 188948 57724
rect 189080 57672 189132 57724
rect 190092 57672 190144 57724
rect 190644 57672 190696 57724
rect 191656 57672 191708 57724
rect 192024 57672 192076 57724
rect 192760 57672 192812 57724
rect 194876 57672 194928 57724
rect 195704 57672 195756 57724
rect 196348 57672 196400 57724
rect 196992 57672 197044 57724
rect 197636 57672 197688 57724
rect 198464 57672 198516 57724
rect 199016 57672 199068 57724
rect 199752 57672 199804 57724
rect 200856 57672 200908 57724
rect 201316 57672 201368 57724
rect 201776 57672 201828 57724
rect 202512 57672 202564 57724
rect 203524 57672 203576 57724
rect 203984 57672 204036 57724
rect 205088 57672 205140 57724
rect 205548 57672 205600 57724
rect 206284 57672 206336 57724
rect 206836 57672 206888 57724
rect 207112 57672 207164 57724
rect 208216 57672 208268 57724
rect 208308 57672 208360 57724
rect 216864 57672 216916 57724
rect 219440 57808 219492 57860
rect 225420 57808 225472 57860
rect 218428 57740 218480 57792
rect 221648 57740 221700 57792
rect 223304 57740 223356 57792
rect 269764 57808 269816 57860
rect 221464 57672 221516 57724
rect 221832 57672 221884 57724
rect 226984 57672 227036 57724
rect 148692 57604 148744 57656
rect 347136 57604 347188 57656
rect 140964 57536 141016 57588
rect 24768 57468 24820 57520
rect 66076 57468 66128 57520
rect 66168 57468 66220 57520
rect 76564 57468 76616 57520
rect 82820 57468 82872 57520
rect 84016 57468 84068 57520
rect 87328 57468 87380 57520
rect 88156 57468 88208 57520
rect 88524 57468 88576 57520
rect 89536 57468 89588 57520
rect 90640 57468 90692 57520
rect 90916 57468 90968 57520
rect 93032 57468 93084 57520
rect 93676 57468 93728 57520
rect 93860 57468 93912 57520
rect 95056 57468 95108 57520
rect 95700 57468 95752 57520
rect 96344 57468 96396 57520
rect 96620 57468 96672 57520
rect 97632 57468 97684 57520
rect 104164 57468 104216 57520
rect 26148 57400 26200 57452
rect 66352 57400 66404 57452
rect 70216 57400 70268 57452
rect 75092 57400 75144 57452
rect 75184 57400 75236 57452
rect 78588 57400 78640 57452
rect 81624 57400 81676 57452
rect 82452 57400 82504 57452
rect 87604 57400 87656 57452
rect 88248 57400 88300 57452
rect 96896 57400 96948 57452
rect 97816 57400 97868 57452
rect 98092 57400 98144 57452
rect 99288 57400 99340 57452
rect 103980 57400 104032 57452
rect 132040 57400 132092 57452
rect 132960 57468 133012 57520
rect 137284 57468 137336 57520
rect 137376 57468 137428 57520
rect 141608 57468 141660 57520
rect 142528 57468 142580 57520
rect 146852 57468 146904 57520
rect 148416 57536 148468 57588
rect 347044 57536 347096 57588
rect 148324 57468 148376 57520
rect 149612 57468 149664 57520
rect 353300 57468 353352 57520
rect 138020 57400 138072 57452
rect 143632 57400 143684 57452
rect 165712 57400 165764 57452
rect 167184 57400 167236 57452
rect 168196 57400 168248 57452
rect 168840 57400 168892 57452
rect 169576 57400 169628 57452
rect 174176 57400 174228 57452
rect 175096 57400 175148 57452
rect 175372 57400 175424 57452
rect 176476 57400 176528 57452
rect 178132 57400 178184 57452
rect 179236 57400 179288 57452
rect 17868 57332 17920 57384
rect 6828 57264 6880 57316
rect 57612 57264 57664 57316
rect 57796 57332 57848 57384
rect 61568 57332 61620 57384
rect 64236 57332 64288 57384
rect 64788 57332 64840 57384
rect 76196 57332 76248 57384
rect 83372 57332 83424 57384
rect 92664 57332 92716 57384
rect 97540 57332 97592 57384
rect 147772 57332 147824 57384
rect 148140 57332 148192 57384
rect 152556 57332 152608 57384
rect 152648 57332 152700 57384
rect 153108 57332 153160 57384
rect 153844 57332 153896 57384
rect 154304 57332 154356 57384
rect 155040 57332 155092 57384
rect 155684 57332 155736 57384
rect 156512 57332 156564 57384
rect 157064 57332 157116 57384
rect 62028 57264 62080 57316
rect 75644 57264 75696 57316
rect 86132 57264 86184 57316
rect 101312 57264 101364 57316
rect 102600 57264 102652 57316
rect 167000 57264 167052 57316
rect 168196 57264 168248 57316
rect 168472 57332 168524 57384
rect 169484 57332 169536 57384
rect 178684 57332 178736 57384
rect 180340 57332 180392 57384
rect 168748 57264 168800 57316
rect 179604 57264 179656 57316
rect 180708 57264 180760 57316
rect 180800 57264 180852 57316
rect 183560 57264 183612 57316
rect 3976 57196 4028 57248
rect 60648 57196 60700 57248
rect 60832 57196 60884 57248
rect 75000 57196 75052 57248
rect 35808 57128 35860 57180
rect 68744 57128 68796 57180
rect 68928 57128 68980 57180
rect 77116 57196 77168 57248
rect 87052 57196 87104 57248
rect 102968 57196 103020 57248
rect 76564 57128 76616 57180
rect 78036 57128 78088 57180
rect 91192 57128 91244 57180
rect 97264 57128 97316 57180
rect 98368 57128 98420 57180
rect 99012 57128 99064 57180
rect 103520 57128 103572 57180
rect 41328 57060 41380 57112
rect 70124 57060 70176 57112
rect 94964 57060 95016 57112
rect 104164 57060 104216 57112
rect 43444 56992 43496 57044
rect 70492 56992 70544 57044
rect 46848 56924 46900 56976
rect 71688 56924 71740 56976
rect 48228 56856 48280 56908
rect 72056 56856 72108 56908
rect 72148 56856 72200 56908
rect 74172 56856 74224 56908
rect 53748 56788 53800 56840
rect 73528 56788 73580 56840
rect 55128 56720 55180 56772
rect 73804 56720 73856 56772
rect 59268 56652 59320 56704
rect 74724 56992 74776 57044
rect 77208 56992 77260 57044
rect 79232 56992 79284 57044
rect 84936 56992 84988 57044
rect 87604 56992 87656 57044
rect 92296 56992 92348 57044
rect 106188 57060 106240 57112
rect 113824 57060 113876 57112
rect 171600 57196 171652 57248
rect 176844 57196 176896 57248
rect 180432 57196 180484 57248
rect 181352 57196 181404 57248
rect 181996 57196 182048 57248
rect 182272 57196 182324 57248
rect 183284 57196 183336 57248
rect 186504 57400 186556 57452
rect 187516 57400 187568 57452
rect 187608 57400 187660 57452
rect 190368 57400 190420 57452
rect 411904 57400 411956 57452
rect 418804 57332 418856 57384
rect 425704 57264 425756 57316
rect 429844 57196 429896 57248
rect 114284 57128 114336 57180
rect 146392 57128 146444 57180
rect 152004 57128 152056 57180
rect 153016 57128 153068 57180
rect 153476 57128 153528 57180
rect 154212 57128 154264 57180
rect 154764 57128 154816 57180
rect 155868 57128 155920 57180
rect 155960 57128 156012 57180
rect 156880 57128 156932 57180
rect 157340 57128 157392 57180
rect 216680 57128 216732 57180
rect 117596 57060 117648 57112
rect 118516 57060 118568 57112
rect 95332 56924 95384 56976
rect 102784 56924 102836 56976
rect 94228 56856 94280 56908
rect 104256 56856 104308 56908
rect 80980 56788 81032 56840
rect 83096 56788 83148 56840
rect 105268 56720 105320 56772
rect 106188 56720 106240 56772
rect 99564 56652 99616 56704
rect 100668 56652 100720 56704
rect 101128 56652 101180 56704
rect 101864 56652 101916 56704
rect 102324 56652 102376 56704
rect 103060 56652 103112 56704
rect 104348 56652 104400 56704
rect 104808 56652 104860 56704
rect 104992 56652 105044 56704
rect 105820 56652 105872 56704
rect 106464 56652 106516 56704
rect 107568 56652 107620 56704
rect 57244 56584 57296 56636
rect 72148 56584 72200 56636
rect 72424 56584 72476 56636
rect 75920 56584 75972 56636
rect 98736 56584 98788 56636
rect 99196 56584 99248 56636
rect 99932 56584 99984 56636
rect 100392 56584 100444 56636
rect 101680 56584 101732 56636
rect 102048 56584 102100 56636
rect 102876 56584 102928 56636
rect 103428 56584 103480 56636
rect 104072 56584 104124 56636
rect 104532 56584 104584 56636
rect 105544 56584 105596 56636
rect 106096 56584 106148 56636
rect 106740 56584 106792 56636
rect 107476 56584 107528 56636
rect 107660 56584 107712 56636
rect 108488 56584 108540 56636
rect 113364 56924 113416 56976
rect 115480 56856 115532 56908
rect 115848 56856 115900 56908
rect 143540 57060 143592 57112
rect 146300 57060 146352 57112
rect 155132 57060 155184 57112
rect 156236 57060 156288 57112
rect 157248 57060 157300 57112
rect 218704 57128 218756 57180
rect 218980 57128 219032 57180
rect 221556 57128 221608 57180
rect 121736 56992 121788 57044
rect 127716 56992 127768 57044
rect 128452 56992 128504 57044
rect 136640 56992 136692 57044
rect 140044 56992 140096 57044
rect 122656 56924 122708 56976
rect 127808 56924 127860 56976
rect 109500 56788 109552 56840
rect 110236 56788 110288 56840
rect 110696 56788 110748 56840
rect 111708 56788 111760 56840
rect 111892 56788 111944 56840
rect 112904 56788 112956 56840
rect 113732 56788 113784 56840
rect 124864 56856 124916 56908
rect 123576 56788 123628 56840
rect 109776 56720 109828 56772
rect 110328 56720 110380 56772
rect 110420 56720 110472 56772
rect 111432 56720 111484 56772
rect 112168 56720 112220 56772
rect 112996 56720 113048 56772
rect 114560 56720 114612 56772
rect 115480 56720 115532 56772
rect 116676 56720 116728 56772
rect 117044 56720 117096 56772
rect 120264 56720 120316 56772
rect 121276 56720 121328 56772
rect 109224 56652 109276 56704
rect 109960 56652 110012 56704
rect 110972 56652 111024 56704
rect 111524 56652 111576 56704
rect 112720 56652 112772 56704
rect 113088 56652 113140 56704
rect 113640 56652 113692 56704
rect 114468 56652 114520 56704
rect 114836 56652 114888 56704
rect 115572 56652 115624 56704
rect 116400 56652 116452 56704
rect 116860 56652 116912 56704
rect 127716 56788 127768 56840
rect 144184 56924 144236 56976
rect 128360 56856 128412 56908
rect 129372 56856 129424 56908
rect 131856 56856 131908 56908
rect 135352 56856 135404 56908
rect 139124 56856 139176 56908
rect 146116 56856 146168 56908
rect 152556 56992 152608 57044
rect 159364 56992 159416 57044
rect 149152 56924 149204 56976
rect 150164 56924 150216 56976
rect 155316 56924 155368 56976
rect 216864 57060 216916 57112
rect 225696 57060 225748 57112
rect 158812 56856 158864 56908
rect 158904 56856 158956 56908
rect 170312 56924 170364 56976
rect 170864 56924 170916 56976
rect 163412 56856 163464 56908
rect 217140 56924 217192 56976
rect 217416 56992 217468 57044
rect 218980 56992 219032 57044
rect 218612 56924 218664 56976
rect 218796 56924 218848 56976
rect 258724 56924 258776 56976
rect 175004 56856 175056 56908
rect 180524 56856 180576 56908
rect 133144 56788 133196 56840
rect 133788 56788 133840 56840
rect 134064 56788 134116 56840
rect 135076 56788 135128 56840
rect 138572 56788 138624 56840
rect 143632 56788 143684 56840
rect 145472 56788 145524 56840
rect 125968 56720 126020 56772
rect 126796 56720 126848 56772
rect 141884 56720 141936 56772
rect 145104 56720 145156 56772
rect 147680 56720 147732 56772
rect 149060 56720 149112 56772
rect 150256 56720 150308 56772
rect 150808 56788 150860 56840
rect 151636 56788 151688 56840
rect 177304 56788 177356 56840
rect 154120 56720 154172 56772
rect 157340 56720 157392 56772
rect 157432 56720 157484 56772
rect 171508 56720 171560 56772
rect 180892 56788 180944 56840
rect 181904 56788 181956 56840
rect 184112 56788 184164 56840
rect 184664 56788 184716 56840
rect 184940 56788 184992 56840
rect 186044 56788 186096 56840
rect 189448 56788 189500 56840
rect 190276 56788 190328 56840
rect 191288 56788 191340 56840
rect 191564 56788 191616 56840
rect 192208 56788 192260 56840
rect 192944 56788 192996 56840
rect 193404 56788 193456 56840
rect 194232 56788 194284 56840
rect 196900 56788 196952 56840
rect 197268 56788 197320 56840
rect 197820 56788 197872 56840
rect 198648 56788 198700 56840
rect 199660 56788 199712 56840
rect 199936 56788 199988 56840
rect 200580 56856 200632 56908
rect 201408 56856 201460 56908
rect 202328 56856 202380 56908
rect 202696 56856 202748 56908
rect 203248 56856 203300 56908
rect 203892 56856 203944 56908
rect 204444 56856 204496 56908
rect 205364 56856 205416 56908
rect 205640 56856 205692 56908
rect 206652 56856 206704 56908
rect 207480 56856 207532 56908
rect 208308 56856 208360 56908
rect 210424 56856 210476 56908
rect 229560 56856 229612 56908
rect 179880 56720 179932 56772
rect 180524 56720 180576 56772
rect 129832 56652 129884 56704
rect 130936 56652 130988 56704
rect 131396 56652 131448 56704
rect 132316 56652 132368 56704
rect 132592 56652 132644 56704
rect 133604 56652 133656 56704
rect 134616 56652 134668 56704
rect 135168 56652 135220 56704
rect 135260 56652 135312 56704
rect 136088 56652 136140 56704
rect 136272 56652 136324 56704
rect 120540 56584 120592 56636
rect 121368 56584 121420 56636
rect 121460 56584 121512 56636
rect 122748 56584 122800 56636
rect 122932 56584 122984 56636
rect 123760 56584 123812 56636
rect 124772 56584 124824 56636
rect 125416 56584 125468 56636
rect 125692 56584 125744 56636
rect 126428 56584 126480 56636
rect 127164 56584 127216 56636
rect 117872 56516 117924 56568
rect 127256 56516 127308 56568
rect 122012 56448 122064 56500
rect 127440 56584 127492 56636
rect 127992 56584 128044 56636
rect 127900 56516 127952 56568
rect 128912 56584 128964 56636
rect 129464 56584 129516 56636
rect 130108 56584 130160 56636
rect 130660 56584 130712 56636
rect 131120 56584 131172 56636
rect 131672 56584 131724 56636
rect 132408 56584 132460 56636
rect 132868 56584 132920 56636
rect 133328 56584 133380 56636
rect 134340 56584 134392 56636
rect 134892 56584 134944 56636
rect 135812 56584 135864 56636
rect 136548 56584 136600 56636
rect 137008 56584 137060 56636
rect 137744 56584 137796 56636
rect 141424 56652 141476 56704
rect 146668 56652 146720 56704
rect 147404 56652 147456 56704
rect 149888 56652 149940 56704
rect 150348 56652 150400 56704
rect 150716 56652 150768 56704
rect 151360 56652 151412 56704
rect 157984 56652 158036 56704
rect 158444 56652 158496 56704
rect 158536 56652 158588 56704
rect 160744 56652 160796 56704
rect 161388 56652 161440 56704
rect 164332 56652 164384 56704
rect 165068 56652 165120 56704
rect 165804 56652 165856 56704
rect 166816 56652 166868 56704
rect 138204 56584 138256 56636
rect 139308 56584 139360 56636
rect 139768 56584 139820 56636
rect 140504 56584 140556 56636
rect 141516 56584 141568 56636
rect 142068 56584 142120 56636
rect 142436 56584 142488 56636
rect 143172 56584 143224 56636
rect 144276 56584 144328 56636
rect 144644 56584 144696 56636
rect 145748 56584 145800 56636
rect 146208 56584 146260 56636
rect 147220 56584 147272 56636
rect 147588 56584 147640 56636
rect 149336 56584 149388 56636
rect 150072 56584 150124 56636
rect 151084 56584 151136 56636
rect 151544 56584 151596 56636
rect 157708 56584 157760 56636
rect 158260 56584 158312 56636
rect 158352 56584 158404 56636
rect 158720 56584 158772 56636
rect 159180 56584 159232 56636
rect 159732 56584 159784 56636
rect 160376 56584 160428 56636
rect 160928 56584 160980 56636
rect 161572 56584 161624 56636
rect 162676 56584 162728 56636
rect 163136 56584 163188 56636
rect 163872 56584 163924 56636
rect 164884 56584 164936 56636
rect 165344 56584 165396 56636
rect 166080 56584 166132 56636
rect 166632 56584 166684 56636
rect 173256 56584 173308 56636
rect 181168 56652 181220 56704
rect 182088 56652 182140 56704
rect 182916 56652 182968 56704
rect 183376 56652 183428 56704
rect 183560 56652 183612 56704
rect 190368 56652 190420 56704
rect 196072 56652 196124 56704
rect 197176 56652 197228 56704
rect 198740 56652 198792 56704
rect 199660 56652 199712 56704
rect 180984 56584 181036 56636
rect 187608 56584 187660 56636
rect 201500 56652 201552 56704
rect 202420 56652 202472 56704
rect 203156 56788 203208 56840
rect 203800 56788 203852 56840
rect 205916 56788 205968 56840
rect 206928 56788 206980 56840
rect 208124 56788 208176 56840
rect 233884 56788 233936 56840
rect 209044 56652 209096 56704
rect 271144 56720 271196 56772
rect 214012 56652 214064 56704
rect 228272 56652 228324 56704
rect 213460 56584 213512 56636
rect 225788 56584 225840 56636
rect 163688 56516 163740 56568
rect 407764 56516 407816 56568
rect 128176 56448 128228 56500
rect 167276 56448 167328 56500
rect 421564 56448 421616 56500
rect 183468 56380 183520 56432
rect 443644 56380 443696 56432
rect 185308 56312 185360 56364
rect 450544 56312 450596 56364
rect 184388 56244 184440 56296
rect 447784 56244 447836 56296
rect 186228 56176 186280 56228
rect 454684 56176 454736 56228
rect 187976 56108 188028 56160
rect 461584 56108 461636 56160
rect 189172 56040 189224 56092
rect 472624 56040 472676 56092
rect 187056 55972 187108 56024
rect 500960 55972 501012 56024
rect 188988 55904 189040 55956
rect 507860 55904 507912 55956
rect 202972 55836 203024 55888
rect 564440 55836 564492 55888
rect 139400 55768 139452 55820
rect 313280 55768 313332 55820
rect 118792 55700 118844 55752
rect 231860 55700 231912 55752
rect 116032 55632 116084 55684
rect 220820 55632 220872 55684
rect 115204 55564 115256 55616
rect 218060 55564 218112 55616
rect 218612 55564 218664 55616
rect 219072 55564 219124 55616
rect 112444 55496 112496 55548
rect 113088 55496 113140 55548
rect 127256 55496 127308 55548
rect 227720 55496 227772 55548
rect 103796 55428 103848 55480
rect 104716 55428 104768 55480
rect 119344 55428 119396 55480
rect 119896 55428 119948 55480
rect 130752 55428 130804 55480
rect 131028 55428 131080 55480
rect 146392 55428 146444 55480
rect 213920 55428 213972 55480
rect 143540 55360 143592 55412
rect 209780 55360 209832 55412
rect 100760 55292 100812 55344
rect 102048 55292 102100 55344
rect 130476 55292 130528 55344
rect 131028 55292 131080 55344
rect 142160 55156 142212 55208
rect 324320 55156 324372 55208
rect 143080 55088 143132 55140
rect 327080 55088 327132 55140
rect 143908 55020 143960 55072
rect 331220 55020 331272 55072
rect 162768 54952 162820 55004
rect 405740 54952 405792 55004
rect 164608 54884 164660 54936
rect 412640 54884 412692 54936
rect 53656 54816 53708 54868
rect 73252 54816 73304 54868
rect 165528 54816 165580 54868
rect 414664 54816 414716 54868
rect 49608 54748 49660 54800
rect 72332 54748 72384 54800
rect 166448 54748 166500 54800
rect 417424 54748 417476 54800
rect 45468 54680 45520 54732
rect 71412 54680 71464 54732
rect 167184 54680 167236 54732
rect 425796 54680 425848 54732
rect 45376 54612 45428 54664
rect 71136 54612 71188 54664
rect 161020 54612 161072 54664
rect 161296 54612 161348 54664
rect 172060 54612 172112 54664
rect 439504 54612 439556 54664
rect 44088 54544 44140 54596
rect 70860 54544 70912 54596
rect 189080 54544 189132 54596
rect 475384 54544 475436 54596
rect 37188 54476 37240 54528
rect 69296 54476 69348 54528
rect 136088 54476 136140 54528
rect 136456 54476 136508 54528
rect 160100 54476 160152 54528
rect 161296 54476 161348 54528
rect 203156 54476 203208 54528
rect 544384 54476 544436 54528
rect 141240 54408 141292 54460
rect 320180 54408 320232 54460
rect 140320 54340 140372 54392
rect 316040 54340 316092 54392
rect 143632 54272 143684 54324
rect 309140 54272 309192 54324
rect 136732 54204 136784 54256
rect 302240 54204 302292 54256
rect 153200 53728 153252 53780
rect 367100 53728 367152 53780
rect 169116 53660 169168 53712
rect 430580 53660 430632 53712
rect 170036 53592 170088 53644
rect 432604 53592 432656 53644
rect 136180 53524 136232 53576
rect 136364 53524 136416 53576
rect 188252 53524 188304 53576
rect 468484 53524 468536 53576
rect 175648 53456 175700 53508
rect 456800 53456 456852 53508
rect 128636 53388 128688 53440
rect 129556 53388 129608 53440
rect 191012 53388 191064 53440
rect 479524 53388 479576 53440
rect 192024 53320 192076 53372
rect 483664 53320 483716 53372
rect 193680 53252 193732 53304
rect 512644 53252 512696 53304
rect 194600 53184 194652 53236
rect 519544 53184 519596 53236
rect 191840 53116 191892 53168
rect 520280 53116 520332 53168
rect 195428 53048 195480 53100
rect 526444 53048 526496 53100
rect 125324 52980 125376 53032
rect 258080 52980 258132 53032
rect 124496 52912 124548 52964
rect 253940 52912 253992 52964
rect 119068 52844 119120 52896
rect 233240 52844 233292 52896
rect 141884 52776 141936 52828
rect 251180 52776 251232 52828
rect 136640 52708 136692 52760
rect 240140 52708 240192 52760
rect 147680 52368 147732 52420
rect 335360 52368 335412 52420
rect 146024 52300 146076 52352
rect 339500 52300 339552 52352
rect 146944 52232 146996 52284
rect 342260 52232 342312 52284
rect 147864 52164 147916 52216
rect 346400 52164 346452 52216
rect 150440 52096 150492 52148
rect 357440 52096 357492 52148
rect 150532 52028 150584 52080
rect 360200 52028 360252 52080
rect 152280 51960 152332 52012
rect 364340 51960 364392 52012
rect 172980 51892 173032 51944
rect 445760 51892 445812 51944
rect 108028 51824 108080 51876
rect 108856 51824 108908 51876
rect 173900 51824 173952 51876
rect 448520 51824 448572 51876
rect 175556 51756 175608 51808
rect 459560 51756 459612 51808
rect 199384 51688 199436 51740
rect 530584 51688 530636 51740
rect 146116 51008 146168 51060
rect 311900 51008 311952 51060
rect 174820 50940 174872 50992
rect 452660 50940 452712 50992
rect 177488 50872 177540 50924
rect 463700 50872 463752 50924
rect 178408 50804 178460 50856
rect 466460 50804 466512 50856
rect 178040 50736 178092 50788
rect 470600 50736 470652 50788
rect 200212 50668 200264 50720
rect 533344 50668 533396 50720
rect 201132 50600 201184 50652
rect 537484 50600 537536 50652
rect 197544 50532 197596 50584
rect 542360 50532 542412 50584
rect 204720 50464 204772 50516
rect 551284 50464 551336 50516
rect 197636 50396 197688 50448
rect 546500 50396 546552 50448
rect 123300 50328 123352 50380
rect 124128 50328 124180 50380
rect 202052 50328 202104 50380
rect 560300 50328 560352 50380
rect 139492 50260 139544 50312
rect 291200 50260 291252 50312
rect 158720 49104 158772 49156
rect 316132 49104 316184 49156
rect 165712 49036 165764 49088
rect 329840 49036 329892 49088
rect 155132 48968 155184 49020
rect 340880 48968 340932 49020
rect 55772 46180 55824 46232
rect 580356 46180 580408 46232
rect 3332 45500 3384 45552
rect 21364 45500 21416 45552
rect 238116 33056 238168 33108
rect 580172 33056 580224 33108
rect 2780 32852 2832 32904
rect 4804 32852 4856 32904
rect 234068 20612 234120 20664
rect 580080 20612 580132 20664
rect 159364 19932 159416 19984
rect 347780 19932 347832 19984
rect 119804 18640 119856 18692
rect 236000 18640 236052 18692
rect 209044 18572 209096 18624
rect 440240 18572 440292 18624
rect 146944 17892 146996 17944
rect 260840 17892 260892 17944
rect 129372 17824 129424 17876
rect 269120 17824 269172 17876
rect 129280 17756 129332 17808
rect 273260 17756 273312 17808
rect 130660 17688 130712 17740
rect 276020 17688 276072 17740
rect 130752 17620 130804 17672
rect 280160 17620 280212 17672
rect 132132 17552 132184 17604
rect 284300 17552 284352 17604
rect 133512 17484 133564 17536
rect 287060 17484 287112 17536
rect 177304 17416 177356 17468
rect 336740 17416 336792 17468
rect 162124 17348 162176 17400
rect 325700 17348 325752 17400
rect 136272 17280 136324 17332
rect 300860 17280 300912 17332
rect 148324 17212 148376 17264
rect 318800 17212 318852 17264
rect 137284 17144 137336 17196
rect 247040 17144 247092 17196
rect 116952 17076 117004 17128
rect 224960 17076 225012 17128
rect 144184 17008 144236 17060
rect 242900 17008 242952 17060
rect 121276 16532 121328 16584
rect 238116 16532 238168 16584
rect 121184 16464 121236 16516
rect 241704 16464 241756 16516
rect 122564 16396 122616 16448
rect 245200 16396 245252 16448
rect 123852 16328 123904 16380
rect 248788 16328 248840 16380
rect 123944 16260 123996 16312
rect 252376 16260 252428 16312
rect 125416 16192 125468 16244
rect 255872 16192 255924 16244
rect 126612 16124 126664 16176
rect 259460 16124 259512 16176
rect 126704 16056 126756 16108
rect 262956 16056 263008 16108
rect 127992 15988 128044 16040
rect 266544 15988 266596 16040
rect 206652 15920 206704 15972
rect 575112 15920 575164 15972
rect 206744 15852 206796 15904
rect 578608 15852 578660 15904
rect 119896 15784 119948 15836
rect 234620 15784 234672 15836
rect 118424 15716 118476 15768
rect 231032 15716 231084 15768
rect 118516 15648 118568 15700
rect 227536 15648 227588 15700
rect 117044 15580 117096 15632
rect 223948 15580 224000 15632
rect 115664 15512 115716 15564
rect 220452 15512 220504 15564
rect 115572 15444 115624 15496
rect 216864 15444 216916 15496
rect 114376 15376 114428 15428
rect 213368 15376 213420 15428
rect 112720 15308 112772 15360
rect 209872 15308 209924 15360
rect 188896 15104 188948 15156
rect 504180 15104 504232 15156
rect 188712 15036 188764 15088
rect 507676 15036 507728 15088
rect 190276 14968 190328 15020
rect 511264 14968 511316 15020
rect 190184 14900 190236 14952
rect 514760 14900 514812 14952
rect 191564 14832 191616 14884
rect 518348 14832 518400 14884
rect 192944 14764 192996 14816
rect 521844 14764 521896 14816
rect 193036 14696 193088 14748
rect 525432 14696 525484 14748
rect 194324 14628 194376 14680
rect 529020 14628 529072 14680
rect 195704 14560 195756 14612
rect 532516 14560 532568 14612
rect 195796 14492 195848 14544
rect 536104 14492 536156 14544
rect 141516 14424 141568 14476
rect 182548 14424 182600 14476
rect 196900 14424 196952 14476
rect 539600 14424 539652 14476
rect 187424 14356 187476 14408
rect 500592 14356 500644 14408
rect 186136 14288 186188 14340
rect 497096 14288 497148 14340
rect 186044 14220 186096 14272
rect 493508 14220 493560 14272
rect 184664 14152 184716 14204
rect 489920 14152 489972 14204
rect 183192 14084 183244 14136
rect 486424 14084 486476 14136
rect 183284 14016 183336 14068
rect 481640 14016 481692 14068
rect 181720 13948 181772 14000
rect 478144 13948 478196 14000
rect 180524 13880 180576 13932
rect 473360 13880 473412 13932
rect 162492 13744 162544 13796
rect 403624 13744 403676 13796
rect 163964 13676 164016 13728
rect 407212 13676 407264 13728
rect 164056 13608 164108 13660
rect 410800 13608 410852 13660
rect 165344 13540 165396 13592
rect 414296 13540 414348 13592
rect 166816 13472 166868 13524
rect 417424 13472 417476 13524
rect 166724 13404 166776 13456
rect 421380 13404 421432 13456
rect 168104 13336 168156 13388
rect 423772 13336 423824 13388
rect 169484 13268 169536 13320
rect 428464 13268 428516 13320
rect 169392 13200 169444 13252
rect 432052 13200 432104 13252
rect 170864 13132 170916 13184
rect 435548 13132 435600 13184
rect 172244 13064 172296 13116
rect 439136 13064 439188 13116
rect 161020 12996 161072 13048
rect 398840 12996 398892 13048
rect 161112 12928 161164 12980
rect 396540 12928 396592 12980
rect 159824 12860 159876 12912
rect 393044 12860 393096 12912
rect 158352 12792 158404 12844
rect 389456 12792 389508 12844
rect 158260 12724 158312 12776
rect 385960 12724 386012 12776
rect 156972 12656 157024 12708
rect 382372 12656 382424 12708
rect 156880 12588 156932 12640
rect 378876 12588 378928 12640
rect 155684 12520 155736 12572
rect 374000 12520 374052 12572
rect 137744 12384 137796 12436
rect 304356 12384 304408 12436
rect 137836 12316 137888 12368
rect 307944 12316 307996 12368
rect 139216 12248 139268 12300
rect 311440 12248 311492 12300
rect 140504 12180 140556 12232
rect 315028 12180 315080 12232
rect 140596 12112 140648 12164
rect 318524 12112 318576 12164
rect 142068 12044 142120 12096
rect 322112 12044 322164 12096
rect 143172 11976 143224 12028
rect 325608 11976 325660 12028
rect 143356 11908 143408 11960
rect 329196 11908 329248 11960
rect 144644 11840 144696 11892
rect 332692 11840 332744 11892
rect 175096 11772 175148 11824
rect 450452 11772 450504 11824
rect 177856 11704 177908 11756
rect 465172 11704 465224 11756
rect 136364 11636 136416 11688
rect 299480 11636 299532 11688
rect 136456 11568 136508 11620
rect 297272 11568 297324 11620
rect 134892 11500 134944 11552
rect 293684 11500 293736 11552
rect 133696 11432 133748 11484
rect 290188 11432 290240 11484
rect 133604 11364 133656 11416
rect 286600 11364 286652 11416
rect 130844 11296 130896 11348
rect 279516 11296 279568 11348
rect 130936 11228 130988 11280
rect 276112 11228 276164 11280
rect 128084 11160 128136 11212
rect 268844 11160 268896 11212
rect 128176 11092 128228 11144
rect 265348 11092 265400 11144
rect 209780 11024 209832 11076
rect 210976 11024 211028 11076
rect 197084 10956 197136 11008
rect 541992 10956 542044 11008
rect 108672 10888 108724 10940
rect 188528 10888 188580 10940
rect 198556 10888 198608 10940
rect 545488 10888 545540 10940
rect 108580 10820 108632 10872
rect 190828 10820 190880 10872
rect 199752 10820 199804 10872
rect 547880 10820 547932 10872
rect 108764 10752 108816 10804
rect 192024 10752 192076 10804
rect 199844 10752 199896 10804
rect 552664 10752 552716 10804
rect 110052 10684 110104 10736
rect 193220 10684 193272 10736
rect 201316 10684 201368 10736
rect 556160 10684 556212 10736
rect 110236 10616 110288 10668
rect 195428 10616 195480 10668
rect 202512 10616 202564 10668
rect 559748 10616 559800 10668
rect 110144 10548 110196 10600
rect 197912 10548 197964 10600
rect 202604 10548 202656 10600
rect 563244 10548 563296 10600
rect 111432 10480 111484 10532
rect 199108 10480 199160 10532
rect 203984 10480 204036 10532
rect 566832 10480 566884 10532
rect 111524 10412 111576 10464
rect 201592 10412 201644 10464
rect 205364 10412 205416 10464
rect 570328 10412 570380 10464
rect 111340 10344 111392 10396
rect 201500 10344 201552 10396
rect 205456 10344 205508 10396
rect 572720 10344 572772 10396
rect 112904 10276 112956 10328
rect 205088 10276 205140 10328
rect 206836 10276 206888 10328
rect 577412 10276 577464 10328
rect 196992 10208 197044 10260
rect 538404 10208 538456 10260
rect 118608 10140 118660 10192
rect 229836 10140 229888 10192
rect 117136 10072 117188 10124
rect 226432 10072 226484 10124
rect 116860 10004 116912 10056
rect 222752 10004 222804 10056
rect 115756 9936 115808 9988
rect 218612 9936 218664 9988
rect 115480 9868 115532 9920
rect 215668 9868 215720 9920
rect 114468 9800 114520 9852
rect 212172 9800 212224 9852
rect 112812 9732 112864 9784
rect 208584 9732 208636 9784
rect 173716 9596 173768 9648
rect 448612 9596 448664 9648
rect 175188 9528 175240 9580
rect 452108 9528 452160 9580
rect 176476 9460 176528 9512
rect 455696 9460 455748 9512
rect 101680 9392 101732 9444
rect 163688 9392 163740 9444
rect 176384 9392 176436 9444
rect 459192 9392 459244 9444
rect 103244 9324 103296 9376
rect 167184 9324 167236 9376
rect 177948 9324 178000 9376
rect 462780 9324 462832 9376
rect 103336 9256 103388 9308
rect 170680 9256 170732 9308
rect 179236 9256 179288 9308
rect 466276 9256 466328 9308
rect 104532 9188 104584 9240
rect 174268 9188 174320 9240
rect 179328 9188 179380 9240
rect 469864 9188 469916 9240
rect 105912 9120 105964 9172
rect 177856 9120 177908 9172
rect 180616 9120 180668 9172
rect 473452 9120 473504 9172
rect 106004 9052 106056 9104
rect 181444 9052 181496 9104
rect 181904 9052 181956 9104
rect 476948 9052 477000 9104
rect 107476 8984 107528 9036
rect 184940 8984 184992 9036
rect 185952 8984 186004 9036
rect 495900 8984 495952 9036
rect 107384 8916 107436 8968
rect 187332 8916 187384 8968
rect 187516 8916 187568 8968
rect 499396 8916 499448 8968
rect 172336 8848 172388 8900
rect 443828 8848 443880 8900
rect 173808 8780 173860 8832
rect 445024 8780 445076 8832
rect 172152 8712 172204 8764
rect 441528 8712 441580 8764
rect 170956 8644 171008 8696
rect 437940 8644 437992 8696
rect 168196 8576 168248 8628
rect 422576 8576 422628 8628
rect 166632 8508 166684 8560
rect 418988 8508 419040 8560
rect 97264 8440 97316 8492
rect 103704 8440 103756 8492
rect 162584 8440 162636 8492
rect 404820 8440 404872 8492
rect 162676 8372 162728 8424
rect 401324 8372 401376 8424
rect 158444 8304 158496 8356
rect 387156 8304 387208 8356
rect 152924 8236 152976 8288
rect 367008 8236 367060 8288
rect 154304 8168 154356 8220
rect 370596 8168 370648 8220
rect 155868 8100 155920 8152
rect 374092 8100 374144 8152
rect 155776 8032 155828 8084
rect 377680 8032 377732 8084
rect 157064 7964 157116 8016
rect 381176 7964 381228 8016
rect 94964 7896 95016 7948
rect 137652 7896 137704 7948
rect 158536 7896 158588 7948
rect 384764 7896 384816 7948
rect 96344 7828 96396 7880
rect 141240 7828 141292 7880
rect 158628 7828 158680 7880
rect 388260 7828 388312 7880
rect 97632 7760 97684 7812
rect 144736 7760 144788 7812
rect 159916 7760 159968 7812
rect 391848 7760 391900 7812
rect 99012 7692 99064 7744
rect 151820 7692 151872 7744
rect 161296 7692 161348 7744
rect 395344 7692 395396 7744
rect 86316 7624 86368 7676
rect 97448 7624 97500 7676
rect 98920 7624 98972 7676
rect 155408 7624 155460 7676
rect 161204 7624 161256 7676
rect 398932 7624 398984 7676
rect 85488 7556 85540 7608
rect 98828 7556 98880 7608
rect 100392 7556 100444 7608
rect 158904 7556 158956 7608
rect 162400 7556 162452 7608
rect 402520 7556 402572 7608
rect 153016 7488 153068 7540
rect 363512 7488 363564 7540
rect 151544 7420 151596 7472
rect 359924 7420 359976 7472
rect 150072 7352 150124 7404
rect 356336 7352 356388 7404
rect 150164 7284 150216 7336
rect 352840 7284 352892 7336
rect 147496 7216 147548 7268
rect 345756 7216 345808 7268
rect 147404 7148 147456 7200
rect 342168 7148 342220 7200
rect 146208 7080 146260 7132
rect 338672 7080 338724 7132
rect 144828 7012 144880 7064
rect 335084 7012 335136 7064
rect 128268 6808 128320 6860
rect 267740 6808 267792 6860
rect 129464 6740 129516 6792
rect 270408 6740 270460 6792
rect 129648 6672 129700 6724
rect 274824 6672 274876 6724
rect 131028 6604 131080 6656
rect 278320 6604 278372 6656
rect 132316 6536 132368 6588
rect 281908 6536 281960 6588
rect 132224 6468 132276 6520
rect 285404 6468 285456 6520
rect 133788 6400 133840 6452
rect 288992 6400 289044 6452
rect 135076 6332 135128 6384
rect 292580 6332 292632 6384
rect 93676 6264 93728 6316
rect 130568 6264 130620 6316
rect 134984 6264 135036 6316
rect 296076 6264 296128 6316
rect 95056 6196 95108 6248
rect 134156 6196 134208 6248
rect 136548 6196 136600 6248
rect 299664 6196 299716 6248
rect 83832 6128 83884 6180
rect 93952 6128 94004 6180
rect 129556 6128 129608 6180
rect 271236 6128 271288 6180
rect 126888 6060 126940 6112
rect 264152 6060 264204 6112
rect 271144 6060 271196 6112
rect 447416 6128 447468 6180
rect 126796 5992 126848 6044
rect 260656 5992 260708 6044
rect 125232 5924 125284 5976
rect 257068 5924 257120 5976
rect 124036 5856 124088 5908
rect 253480 5856 253532 5908
rect 124128 5788 124180 5840
rect 249984 5788 250036 5840
rect 122656 5720 122708 5772
rect 246396 5720 246448 5772
rect 122748 5652 122800 5704
rect 242992 5652 243044 5704
rect 121368 5584 121420 5636
rect 239312 5584 239364 5636
rect 119712 5516 119764 5568
rect 235816 5516 235868 5568
rect 101772 5448 101824 5500
rect 166080 5448 166132 5500
rect 197268 5448 197320 5500
rect 540796 5448 540848 5500
rect 103428 5380 103480 5432
rect 169576 5380 169628 5432
rect 198648 5380 198700 5432
rect 544292 5380 544344 5432
rect 104716 5312 104768 5364
rect 173164 5312 173216 5364
rect 199660 5312 199712 5364
rect 547972 5312 548024 5364
rect 102784 5244 102836 5296
rect 103428 5244 103480 5296
rect 104624 5244 104676 5296
rect 176660 5244 176712 5296
rect 199936 5244 199988 5296
rect 551468 5244 551520 5296
rect 106096 5176 106148 5228
rect 180248 5176 180300 5228
rect 202420 5176 202472 5228
rect 107568 5108 107620 5160
rect 183744 5108 183796 5160
rect 202696 5108 202748 5160
rect 205824 5176 205876 5228
rect 554964 5176 555016 5228
rect 108856 5040 108908 5092
rect 189724 5040 189776 5092
rect 203892 5040 203944 5092
rect 558552 5108 558604 5160
rect 108948 4972 109000 5024
rect 193312 4972 193364 5024
rect 194232 4972 194284 5024
rect 204996 4972 205048 5024
rect 562048 5040 562100 5092
rect 565636 4972 565688 5024
rect 110328 4904 110380 4956
rect 196808 4904 196860 4956
rect 204076 4904 204128 4956
rect 569132 4904 569184 4956
rect 111708 4836 111760 4888
rect 200304 4836 200356 4888
rect 201408 4836 201460 4888
rect 111616 4768 111668 4820
rect 203892 4768 203944 4820
rect 205548 4836 205600 4888
rect 572812 4836 572864 4888
rect 205824 4768 205876 4820
rect 206928 4768 206980 4820
rect 576308 4768 576360 4820
rect 101864 4700 101916 4752
rect 162492 4700 162544 4752
rect 197176 4700 197228 4752
rect 537208 4700 537260 4752
rect 100484 4632 100536 4684
rect 157800 4632 157852 4684
rect 99104 4564 99156 4616
rect 154212 4564 154264 4616
rect 195520 4564 195572 4616
rect 533712 4632 533764 4684
rect 97724 4496 97776 4548
rect 147128 4496 147180 4548
rect 194508 4496 194560 4548
rect 530124 4564 530176 4616
rect 204996 4496 205048 4548
rect 526628 4496 526680 4548
rect 96436 4428 96488 4480
rect 143540 4428 143592 4480
rect 192760 4428 192812 4480
rect 523040 4428 523092 4480
rect 95148 4360 95200 4412
rect 136456 4360 136508 4412
rect 141424 4360 141476 4412
rect 186136 4360 186188 4412
rect 191472 4360 191524 4412
rect 519544 4360 519596 4412
rect 93768 4292 93820 4344
rect 132960 4292 133012 4344
rect 191656 4292 191708 4344
rect 515956 4292 516008 4344
rect 92296 4224 92348 4276
rect 126980 4224 127032 4276
rect 190092 4224 190144 4276
rect 512460 4224 512512 4276
rect 276020 4156 276072 4208
rect 277124 4156 277176 4208
rect 28908 4088 28960 4140
rect 52460 4088 52512 4140
rect 52552 4088 52604 4140
rect 53656 4088 53708 4140
rect 56048 4088 56100 4140
rect 57244 4088 57296 4140
rect 58440 4088 58492 4140
rect 59268 4088 59320 4140
rect 59636 4088 59688 4140
rect 60648 4088 60700 4140
rect 82452 4088 82504 4140
rect 85672 4088 85724 4140
rect 91008 4088 91060 4140
rect 117596 4088 117648 4140
rect 139308 4088 139360 4140
rect 309048 4088 309100 4140
rect 421564 4088 421616 4140
rect 423680 4088 423732 4140
rect 439504 4088 439556 4140
rect 442632 4088 442684 4140
rect 472624 4088 472676 4140
rect 510068 4088 510120 4140
rect 23020 4020 23072 4072
rect 65708 4020 65760 4072
rect 71504 4020 71556 4072
rect 76564 4020 76616 4072
rect 90732 4020 90784 4072
rect 118792 4020 118844 4072
rect 144552 4020 144604 4072
rect 333888 4020 333940 4072
rect 479524 4020 479576 4072
rect 517152 4020 517204 4072
rect 19432 3952 19484 4004
rect 27620 3952 27672 4004
rect 20628 3884 20680 3936
rect 65156 3952 65208 4004
rect 88064 3952 88116 4004
rect 111616 3952 111668 4004
rect 113088 3952 113140 4004
rect 201408 3952 201460 4004
rect 201500 3952 201552 4004
rect 202696 3952 202748 4004
rect 218980 3952 219032 4004
rect 408408 3952 408460 4004
rect 468484 3952 468536 4004
rect 506480 3952 506532 4004
rect 27804 3884 27856 3936
rect 64972 3884 65024 3936
rect 89628 3884 89680 3936
rect 116400 3884 116452 3936
rect 147588 3884 147640 3936
rect 344560 3884 344612 3936
rect 447784 3884 447836 3936
rect 491116 3884 491168 3936
rect 18236 3816 18288 3868
rect 52368 3816 52420 3868
rect 52460 3816 52512 3868
rect 15936 3748 15988 3800
rect 56140 3816 56192 3868
rect 61844 3816 61896 3868
rect 90640 3816 90692 3868
rect 119896 3816 119948 3868
rect 150256 3816 150308 3868
rect 351644 3816 351696 3868
rect 425704 3816 425756 3868
rect 468668 3816 468720 3868
rect 475384 3816 475436 3868
rect 513564 3816 513616 3868
rect 12256 3680 12308 3732
rect 55496 3680 55548 3732
rect 67272 3748 67324 3800
rect 82636 3748 82688 3800
rect 87972 3748 88024 3800
rect 90916 3748 90968 3800
rect 121092 3748 121144 3800
rect 122104 3748 122156 3800
rect 128176 3748 128228 3800
rect 150348 3748 150400 3800
rect 355232 3748 355284 3800
rect 418804 3748 418856 3800
rect 461584 3748 461636 3800
rect 461676 3748 461728 3800
rect 505376 3748 505428 3800
rect 63960 3680 64012 3732
rect 84016 3680 84068 3732
rect 90364 3680 90416 3732
rect 90824 3680 90876 3732
rect 122288 3680 122340 3732
rect 160008 3680 160060 3732
rect 394240 3680 394292 3732
rect 411996 3680 412048 3732
rect 454500 3680 454552 3732
rect 454684 3680 454736 3732
rect 498200 3680 498252 3732
rect 537484 3680 537536 3732
rect 557356 3680 557408 3732
rect 7656 3612 7708 3664
rect 56140 3612 56192 3664
rect 1676 3544 1728 3596
rect 2872 3476 2924 3528
rect 3976 3476 4028 3528
rect 5264 3544 5316 3596
rect 61292 3612 61344 3664
rect 82544 3612 82596 3664
rect 89168 3612 89220 3664
rect 92388 3612 92440 3664
rect 124680 3612 124732 3664
rect 138664 3612 138716 3664
rect 140044 3612 140096 3664
rect 161388 3612 161440 3664
rect 397736 3612 397788 3664
rect 443644 3612 443696 3664
rect 64328 3544 64380 3596
rect 64788 3544 64840 3596
rect 55220 3476 55272 3528
rect 55496 3476 55548 3528
rect 60004 3476 60056 3528
rect 63224 3476 63276 3528
rect 72424 3544 72476 3596
rect 75000 3544 75052 3596
rect 75828 3544 75880 3596
rect 81348 3544 81400 3596
rect 65524 3476 65576 3528
rect 66168 3476 66220 3528
rect 66720 3476 66772 3528
rect 67548 3476 67600 3528
rect 67916 3476 67968 3528
rect 68928 3476 68980 3528
rect 69112 3476 69164 3528
rect 70216 3476 70268 3528
rect 72608 3476 72660 3528
rect 73068 3476 73120 3528
rect 572 3408 624 3460
rect 59360 3408 59412 3460
rect 60832 3408 60884 3460
rect 75368 3476 75420 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 79692 3476 79744 3528
rect 80336 3476 80388 3528
rect 80428 3476 80480 3528
rect 80888 3476 80940 3528
rect 81256 3476 81308 3528
rect 82084 3476 82136 3528
rect 84108 3544 84160 3596
rect 91560 3544 91612 3596
rect 97816 3544 97868 3596
rect 84476 3476 84528 3528
rect 73804 3408 73856 3460
rect 75184 3408 75236 3460
rect 83924 3408 83976 3460
rect 95148 3476 95200 3528
rect 96528 3476 96580 3528
rect 98460 3476 98512 3528
rect 98828 3476 98880 3528
rect 100668 3544 100720 3596
rect 8760 3340 8812 3392
rect 9588 3340 9640 3392
rect 9956 3340 10008 3392
rect 10968 3340 11020 3392
rect 11152 3340 11204 3392
rect 12348 3340 12400 3392
rect 17040 3340 17092 3392
rect 17868 3340 17920 3392
rect 25320 3340 25372 3392
rect 26148 3340 26200 3392
rect 27712 3340 27764 3392
rect 28816 3340 28868 3392
rect 32404 3340 32456 3392
rect 33048 3340 33100 3392
rect 33600 3340 33652 3392
rect 34428 3340 34480 3392
rect 34796 3340 34848 3392
rect 35808 3340 35860 3392
rect 40684 3340 40736 3392
rect 41328 3340 41380 3392
rect 43076 3340 43128 3392
rect 44088 3340 44140 3392
rect 31300 3272 31352 3324
rect 67824 3340 67876 3392
rect 78588 3340 78640 3392
rect 79784 3340 79836 3392
rect 86224 3340 86276 3392
rect 99196 3408 99248 3460
rect 99564 3408 99616 3460
rect 100116 3408 100168 3460
rect 89444 3340 89496 3392
rect 101220 3476 101272 3528
rect 100300 3408 100352 3460
rect 101404 3544 101456 3596
rect 103336 3544 103388 3596
rect 103428 3544 103480 3596
rect 106832 3544 106884 3596
rect 101496 3476 101548 3528
rect 107476 3544 107528 3596
rect 142436 3544 142488 3596
rect 165252 3544 165304 3596
rect 415492 3544 415544 3596
rect 429844 3544 429896 3596
rect 145932 3476 145984 3528
rect 168012 3476 168064 3528
rect 48964 3272 49016 3324
rect 49608 3272 49660 3324
rect 41880 3204 41932 3256
rect 43444 3204 43496 3256
rect 38384 3136 38436 3188
rect 44272 3136 44324 3188
rect 45376 3136 45428 3188
rect 55772 3136 55824 3188
rect 35992 3068 36044 3120
rect 69204 3272 69256 3324
rect 88984 3272 89036 3324
rect 96252 3272 96304 3324
rect 101036 3340 101088 3392
rect 102324 3408 102376 3460
rect 102876 3408 102928 3460
rect 106924 3408 106976 3460
rect 110144 3408 110196 3460
rect 156604 3408 156656 3460
rect 169668 3408 169720 3460
rect 107016 3340 107068 3392
rect 107108 3340 107160 3392
rect 110512 3340 110564 3392
rect 110604 3340 110656 3392
rect 123484 3340 123536 3392
rect 124864 3340 124916 3392
rect 125876 3340 125928 3392
rect 137744 3340 137796 3392
rect 306748 3340 306800 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 347044 3340 347096 3392
rect 349252 3340 349304 3392
rect 374000 3340 374052 3392
rect 375288 3340 375340 3392
rect 398840 3340 398892 3392
rect 400128 3340 400180 3392
rect 407764 3340 407816 3392
rect 409604 3340 409656 3392
rect 414664 3408 414716 3460
rect 416688 3408 416740 3460
rect 423772 3476 423824 3528
rect 424968 3476 425020 3528
rect 425796 3476 425848 3528
rect 427268 3476 427320 3528
rect 448520 3544 448572 3596
rect 449808 3544 449860 3596
rect 450544 3612 450596 3664
rect 494704 3612 494756 3664
rect 519636 3612 519688 3664
rect 531320 3612 531372 3664
rect 533344 3612 533396 3664
rect 553768 3612 553820 3664
rect 487620 3544 487672 3596
rect 512644 3544 512696 3596
rect 527824 3544 527876 3596
rect 530584 3544 530636 3596
rect 550272 3544 550324 3596
rect 551284 3544 551336 3596
rect 571524 3544 571576 3596
rect 426164 3408 426216 3460
rect 432604 3408 432656 3460
rect 434444 3408 434496 3460
rect 436836 3408 436888 3460
rect 429660 3340 429712 3392
rect 115204 3272 115256 3324
rect 135168 3272 135220 3324
rect 294880 3272 294932 3324
rect 299480 3272 299532 3324
rect 300768 3272 300820 3324
rect 347136 3272 347188 3324
rect 350448 3272 350500 3324
rect 473360 3476 473412 3528
rect 474556 3476 474608 3528
rect 481640 3476 481692 3528
rect 482836 3476 482888 3528
rect 483664 3476 483716 3528
rect 524236 3476 524288 3528
rect 526444 3476 526496 3528
rect 534908 3476 534960 3528
rect 544384 3476 544436 3528
rect 568028 3476 568080 3528
rect 572720 3476 572772 3528
rect 573916 3476 573968 3528
rect 475752 3340 475804 3392
rect 581000 3408 581052 3460
rect 547880 3340 547932 3392
rect 549076 3340 549128 3392
rect 55956 3204 56008 3256
rect 69664 3204 69716 3256
rect 89536 3204 89588 3256
rect 112812 3204 112864 3256
rect 112996 3204 113048 3256
rect 206192 3204 206244 3256
rect 218704 3204 218756 3256
rect 376484 3204 376536 3256
rect 72516 3136 72568 3188
rect 77392 3136 77444 3188
rect 79508 3136 79560 3188
rect 88248 3136 88300 3188
rect 109316 3136 109368 3188
rect 55956 3068 56008 3120
rect 56140 3068 56192 3120
rect 72976 3068 73028 3120
rect 86684 3068 86736 3120
rect 105728 3068 105780 3120
rect 106188 3068 106240 3120
rect 126336 3136 126388 3188
rect 129372 3136 129424 3188
rect 132408 3136 132460 3188
rect 283104 3136 283156 3188
rect 179052 3068 179104 3120
rect 193220 3068 193272 3120
rect 194416 3068 194468 3120
rect 201408 3068 201460 3120
rect 207388 3068 207440 3120
rect 221648 3068 221700 3120
rect 371700 3068 371752 3120
rect 24216 3000 24268 3052
rect 24768 3000 24820 3052
rect 57244 3000 57296 3052
rect 74448 3000 74500 3052
rect 88156 3000 88208 3052
rect 108120 3000 108172 3052
rect 26516 2932 26568 2984
rect 27528 2932 27580 2984
rect 50160 2932 50212 2984
rect 55864 2932 55916 2984
rect 52368 2864 52420 2916
rect 64512 2932 64564 2984
rect 86868 2932 86920 2984
rect 104532 2932 104584 2984
rect 104624 2932 104676 2984
rect 219348 3000 219400 3052
rect 323308 3000 323360 3052
rect 417516 3000 417568 3052
rect 420184 3000 420236 3052
rect 114008 2932 114060 2984
rect 221464 2932 221516 2984
rect 305552 2932 305604 2984
rect 86776 2864 86828 2916
rect 102232 2864 102284 2916
rect 102324 2864 102376 2916
rect 103612 2864 103664 2916
rect 103704 2864 103756 2916
rect 110604 2864 110656 2916
rect 221556 2864 221608 2916
rect 298468 2864 298520 2916
rect 55220 2796 55272 2848
rect 59452 2796 59504 2848
rect 82728 2796 82780 2848
rect 86868 2796 86920 2848
rect 87604 2796 87656 2848
rect 98644 2796 98696 2848
rect 98460 2728 98512 2780
rect 99380 2796 99432 2848
rect 103888 2796 103940 2848
rect 110144 2796 110196 2848
rect 242900 2796 242952 2848
rect 244096 2796 244148 2848
rect 270408 2796 270460 2848
rect 272432 2796 272484 2848
rect 154304 2116 154356 2168
rect 369400 2116 369452 2168
rect 154396 2048 154448 2100
rect 372896 2048 372948 2100
rect 99196 960 99248 1012
rect 99840 960 99892 1012
rect 51356 688 51408 740
rect 56140 688 56192 740
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 3422 410544 3478 410553
rect 3422 410479 3478 410488
rect 3436 373318 3464 410479
rect 3516 397520 3568 397526
rect 3514 397488 3516 397497
rect 3568 397488 3570 397497
rect 3514 397423 3570 397432
rect 3424 373312 3476 373318
rect 3424 373254 3476 373260
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 4816 262206 4844 683674
rect 8220 264722 8248 702406
rect 24320 700330 24348 703520
rect 40512 700398 40540 703520
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 33784 700324 33836 700330
rect 33784 700266 33836 700272
rect 21364 656940 21416 656946
rect 21364 656882 21416 656888
rect 11704 632120 11756 632126
rect 11704 632062 11756 632068
rect 8208 264716 8260 264722
rect 8208 264658 8260 264664
rect 4804 262200 4856 262206
rect 4804 262142 4856 262148
rect 11716 261254 11744 632062
rect 14464 579692 14516 579698
rect 14464 579634 14516 579640
rect 14476 261322 14504 579634
rect 15844 527196 15896 527202
rect 15844 527138 15896 527144
rect 14464 261316 14516 261322
rect 14464 261258 14516 261264
rect 11704 261248 11756 261254
rect 11704 261190 11756 261196
rect 15856 260642 15884 527138
rect 17224 474768 17276 474774
rect 17224 474710 17276 474716
rect 17236 261390 17264 474710
rect 18604 422340 18656 422346
rect 18604 422282 18656 422288
rect 18616 261458 18644 422282
rect 21376 262614 21404 656882
rect 22744 605872 22796 605878
rect 22744 605814 22796 605820
rect 22756 262750 22784 605814
rect 25504 553444 25556 553450
rect 25504 553386 25556 553392
rect 22744 262744 22796 262750
rect 22744 262686 22796 262692
rect 25516 262682 25544 553386
rect 29644 501016 29696 501022
rect 29644 500958 29696 500964
rect 25504 262676 25556 262682
rect 25504 262618 25556 262624
rect 21364 262608 21416 262614
rect 21364 262550 21416 262556
rect 18604 261452 18656 261458
rect 18604 261394 18656 261400
rect 17224 261384 17276 261390
rect 17224 261326 17276 261332
rect 29656 261186 29684 500958
rect 32404 448588 32456 448594
rect 32404 448530 32456 448536
rect 32416 262546 32444 448530
rect 33796 264110 33824 700266
rect 35164 670744 35216 670750
rect 35164 670686 35216 670692
rect 35176 264178 35204 670686
rect 36544 618316 36596 618322
rect 36544 618258 36596 618264
rect 36556 264926 36584 618258
rect 39304 565888 39356 565894
rect 39304 565830 39356 565836
rect 39316 373386 39344 565830
rect 39304 373380 39356 373386
rect 39304 373322 39356 373328
rect 36544 264920 36596 264926
rect 36544 264862 36596 264868
rect 35164 264172 35216 264178
rect 35164 264114 35216 264120
rect 33784 264104 33836 264110
rect 33784 264046 33836 264052
rect 32404 262540 32456 262546
rect 32404 262482 32456 262488
rect 29644 261180 29696 261186
rect 29644 261122 29696 261128
rect 41340 260914 41368 700334
rect 72988 700330 73016 703520
rect 58900 700324 58952 700330
rect 58900 700266 58952 700272
rect 72976 700324 73028 700330
rect 72976 700266 73028 700272
rect 43444 514820 43496 514826
rect 43444 514762 43496 514768
rect 43456 373454 43484 514762
rect 53654 488744 53710 488753
rect 53654 488679 53710 488688
rect 53286 488608 53342 488617
rect 53286 488543 53342 488552
rect 47584 462392 47636 462398
rect 47584 462334 47636 462340
rect 43444 373448 43496 373454
rect 43444 373390 43496 373396
rect 47596 264042 47624 462334
rect 53196 265872 53248 265878
rect 53196 265814 53248 265820
rect 47584 264036 47636 264042
rect 47584 263978 47636 263984
rect 41328 260908 41380 260914
rect 41328 260850 41380 260856
rect 15844 260636 15896 260642
rect 15844 260578 15896 260584
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 236745 3464 254079
rect 4066 241088 4122 241097
rect 4122 241046 4200 241074
rect 4066 241023 4122 241032
rect 3422 236736 3478 236745
rect 3422 236671 3478 236680
rect 4172 233889 4200 241046
rect 4158 233880 4214 233889
rect 4158 233815 4214 233824
rect 17222 233472 17278 233481
rect 17222 233407 17278 233416
rect 3514 232248 3570 232257
rect 3514 232183 3570 232192
rect 3422 228304 3478 228313
rect 3422 228239 3478 228248
rect 3056 215280 3108 215286
rect 3056 215222 3108 215228
rect 3068 214985 3096 215222
rect 3054 214976 3110 214985
rect 3054 214911 3110 214920
rect 3332 188896 3384 188902
rect 3330 188864 3332 188873
rect 3384 188864 3386 188873
rect 3330 188799 3386 188808
rect 3056 164212 3108 164218
rect 3056 164154 3108 164160
rect 3068 162897 3096 164154
rect 3054 162888 3110 162897
rect 3054 162823 3110 162832
rect 3056 137964 3108 137970
rect 3056 137906 3108 137912
rect 3068 136785 3096 137906
rect 3054 136776 3110 136785
rect 3054 136711 3110 136720
rect 3332 111784 3384 111790
rect 3332 111726 3384 111732
rect 3344 110673 3372 111726
rect 3330 110664 3386 110673
rect 3330 110599 3386 110608
rect 3240 97980 3292 97986
rect 3240 97922 3292 97928
rect 3252 97617 3280 97922
rect 3238 97608 3294 97617
rect 3238 97543 3294 97552
rect 2964 85536 3016 85542
rect 2964 85478 3016 85484
rect 2976 84697 3004 85478
rect 2962 84688 3018 84697
rect 2962 84623 3018 84632
rect 3332 71732 3384 71738
rect 3332 71674 3384 71680
rect 3344 71641 3372 71674
rect 3330 71632 3386 71641
rect 3330 71567 3386 71576
rect 3332 45552 3384 45558
rect 3330 45520 3332 45529
rect 3384 45520 3386 45529
rect 3330 45455 3386 45464
rect 2780 32904 2832 32910
rect 2780 32846 2832 32852
rect 2792 32473 2820 32846
rect 2778 32464 2834 32473
rect 2778 32399 2834 32408
rect 3436 6497 3464 228239
rect 3528 19417 3556 232183
rect 4802 232112 4858 232121
rect 4802 232047 4858 232056
rect 3606 228576 3662 228585
rect 3606 228511 3662 228520
rect 3620 58585 3648 228511
rect 3790 228440 3846 228449
rect 3790 228375 3846 228384
rect 3698 227080 3754 227089
rect 3698 227015 3754 227024
rect 3712 149841 3740 227015
rect 3804 201929 3832 228375
rect 3790 201920 3846 201929
rect 3790 201855 3846 201864
rect 3698 149832 3754 149841
rect 3698 149767 3754 149776
rect 3606 58576 3662 58585
rect 3606 58511 3662 58520
rect 3976 57248 4028 57254
rect 3976 57190 4028 57196
rect 4066 57216 4122 57225
rect 3514 19408 3570 19417
rect 3514 19343 3570 19352
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 1676 3596 1728 3602
rect 1676 3538 1728 3544
rect 572 3460 624 3466
rect 572 3402 624 3408
rect 584 480 612 3402
rect 1688 480 1716 3538
rect 3988 3534 4016 57190
rect 4066 57151 4122 57160
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 3976 3528 4028 3534
rect 3976 3470 4028 3476
rect 2884 480 2912 3470
rect 4080 480 4108 57151
rect 4816 32910 4844 232047
rect 11702 231296 11758 231305
rect 11702 231231 11758 231240
rect 7562 229120 7618 229129
rect 7562 229055 7618 229064
rect 7576 188902 7604 229055
rect 11716 215286 11744 231231
rect 14462 231160 14518 231169
rect 14462 231095 14518 231104
rect 11704 215280 11756 215286
rect 11704 215222 11756 215228
rect 7564 188896 7616 188902
rect 7564 188838 7616 188844
rect 14476 164218 14504 231095
rect 15842 231024 15898 231033
rect 15842 230959 15898 230968
rect 14464 164212 14516 164218
rect 14464 164154 14516 164160
rect 15856 111790 15884 230959
rect 17236 137970 17264 233407
rect 21362 233336 21418 233345
rect 21362 233271 21418 233280
rect 18602 229256 18658 229265
rect 18602 229191 18658 229200
rect 17224 137964 17276 137970
rect 17224 137906 17276 137912
rect 15844 111784 15896 111790
rect 15844 111726 15896 111732
rect 18616 97986 18644 229191
rect 18604 97980 18656 97986
rect 18604 97922 18656 97928
rect 12346 57624 12402 57633
rect 12346 57559 12402 57568
rect 10966 57488 11022 57497
rect 10966 57423 11022 57432
rect 9586 57352 9642 57361
rect 6828 57316 6880 57322
rect 9586 57287 9642 57296
rect 6828 57258 6880 57264
rect 4804 32904 4856 32910
rect 4804 32846 4856 32852
rect 6840 6914 6868 57258
rect 6472 6886 6868 6914
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5276 480 5304 3538
rect 6472 480 6500 6886
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7668 480 7696 3606
rect 9600 3398 9628 57287
rect 10980 3398 11008 57423
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 8772 480 8800 3334
rect 9968 480 9996 3334
rect 11164 480 11192 3334
rect 12268 1850 12296 3674
rect 12360 3398 12388 57559
rect 17868 57384 17920 57390
rect 17868 57326 17920 57332
rect 15106 57080 15162 57089
rect 15106 57015 15162 57024
rect 13726 56944 13782 56953
rect 13726 56879 13782 56888
rect 13740 6914 13768 56879
rect 15120 6914 15148 57015
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12268 1822 12388 1850
rect 12360 480 12388 1822
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 15936 3800 15988 3806
rect 15936 3742 15988 3748
rect 15948 480 15976 3742
rect 17880 3398 17908 57326
rect 21376 45558 21404 233271
rect 32402 232520 32458 232529
rect 32402 232455 32458 232464
rect 29642 232384 29698 232393
rect 29642 232319 29698 232328
rect 29656 71738 29684 232319
rect 32416 85542 32444 232455
rect 53208 155922 53236 265814
rect 53300 191826 53328 488543
rect 53470 486568 53526 486577
rect 53470 486503 53526 486512
rect 53378 483304 53434 483313
rect 53378 483239 53434 483248
rect 53288 191820 53340 191826
rect 53288 191762 53340 191768
rect 53392 178022 53420 483239
rect 53380 178016 53432 178022
rect 53380 177958 53432 177964
rect 53484 160070 53512 486503
rect 53562 483440 53618 483449
rect 53562 483375 53618 483384
rect 53472 160064 53524 160070
rect 53472 160006 53524 160012
rect 53196 155916 53248 155922
rect 53196 155858 53248 155864
rect 53576 147626 53604 483375
rect 53564 147620 53616 147626
rect 53564 147562 53616 147568
rect 53668 143546 53696 488679
rect 58806 487928 58862 487937
rect 58806 487863 58862 487872
rect 54758 487792 54814 487801
rect 54758 487727 54814 487736
rect 54666 487248 54722 487257
rect 54666 487183 54722 487192
rect 53746 485888 53802 485897
rect 53746 485823 53802 485832
rect 53656 143540 53708 143546
rect 53656 143482 53708 143488
rect 53760 131102 53788 485823
rect 54576 395344 54628 395350
rect 54576 395286 54628 395292
rect 54300 265804 54352 265810
rect 54300 265746 54352 265752
rect 54208 265736 54260 265742
rect 54208 265678 54260 265684
rect 54220 213926 54248 265678
rect 54208 213920 54260 213926
rect 54208 213862 54260 213868
rect 54312 197334 54340 265746
rect 54392 264376 54444 264382
rect 54392 264318 54444 264324
rect 54300 197328 54352 197334
rect 54300 197270 54352 197276
rect 54404 134774 54432 264318
rect 54482 242176 54538 242185
rect 54482 242111 54538 242120
rect 54392 134768 54444 134774
rect 54392 134710 54444 134716
rect 53748 131096 53800 131102
rect 53748 131038 53800 131044
rect 32404 85536 32456 85542
rect 32404 85478 32456 85484
rect 54496 71738 54524 242111
rect 54588 175234 54616 395286
rect 54680 194546 54708 487183
rect 54668 194540 54720 194546
rect 54668 194482 54720 194488
rect 54772 182170 54800 487727
rect 58714 487656 58770 487665
rect 58714 487591 58770 487600
rect 54942 487520 54998 487529
rect 54942 487455 54998 487464
rect 54850 485616 54906 485625
rect 54850 485551 54906 485560
rect 54760 182164 54812 182170
rect 54760 182106 54812 182112
rect 54576 175228 54628 175234
rect 54576 175170 54628 175176
rect 54864 153202 54892 485551
rect 54852 153196 54904 153202
rect 54852 153138 54904 153144
rect 54956 118658 54984 487455
rect 56874 487384 56930 487393
rect 56874 487319 56930 487328
rect 55126 484800 55182 484809
rect 55126 484735 55182 484744
rect 55034 484528 55090 484537
rect 55034 484463 55090 484472
rect 54944 118652 54996 118658
rect 54944 118594 54996 118600
rect 55048 113150 55076 484463
rect 55036 113144 55088 113150
rect 55036 113086 55088 113092
rect 29644 71732 29696 71738
rect 29644 71674 29696 71680
rect 54484 71732 54536 71738
rect 54484 71674 54536 71680
rect 55140 62082 55168 484735
rect 56598 432304 56654 432313
rect 56598 432239 56654 432248
rect 56508 395412 56560 395418
rect 56508 395354 56560 395360
rect 56324 356720 56376 356726
rect 56324 356662 56376 356668
rect 55864 264852 55916 264858
rect 55864 264794 55916 264800
rect 55772 229152 55824 229158
rect 55772 229094 55824 229100
rect 55128 62076 55180 62082
rect 55128 62018 55180 62024
rect 39948 57928 40000 57934
rect 39948 57870 40000 57876
rect 34428 57860 34480 57866
rect 34428 57802 34480 57808
rect 30288 57792 30340 57798
rect 30288 57734 30340 57740
rect 28908 57656 28960 57662
rect 28908 57598 28960 57604
rect 27528 57588 27580 57594
rect 27528 57530 27580 57536
rect 24768 57520 24820 57526
rect 24768 57462 24820 57468
rect 22006 56808 22062 56817
rect 22006 56743 22062 56752
rect 21364 45552 21416 45558
rect 21364 45494 21416 45500
rect 22020 6914 22048 56743
rect 21836 6886 22048 6914
rect 19432 4004 19484 4010
rect 19432 3946 19484 3952
rect 18236 3868 18288 3874
rect 18236 3810 18288 3816
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17052 480 17080 3334
rect 18248 480 18276 3810
rect 19444 480 19472 3946
rect 20628 3936 20680 3942
rect 20628 3878 20680 3884
rect 20640 480 20668 3878
rect 21836 480 21864 6886
rect 23020 4072 23072 4078
rect 23020 4014 23072 4020
rect 23032 480 23060 4014
rect 24780 3058 24808 57462
rect 26148 57452 26200 57458
rect 26148 57394 26200 57400
rect 26160 3398 26188 57394
rect 25320 3392 25372 3398
rect 25320 3334 25372 3340
rect 26148 3392 26200 3398
rect 26148 3334 26200 3340
rect 24216 3052 24268 3058
rect 24216 2994 24268 3000
rect 24768 3052 24820 3058
rect 24768 2994 24820 3000
rect 24228 480 24256 2994
rect 25332 480 25360 3334
rect 27540 2990 27568 57530
rect 28920 6914 28948 57598
rect 30300 6914 30328 57734
rect 33048 57724 33100 57730
rect 33048 57666 33100 57672
rect 28828 6886 28948 6914
rect 30116 6886 30328 6914
rect 27620 4004 27672 4010
rect 27620 3946 27672 3952
rect 27632 3890 27660 3946
rect 27804 3936 27856 3942
rect 27632 3884 27804 3890
rect 27632 3878 27856 3884
rect 27632 3862 27844 3878
rect 28828 3398 28856 6886
rect 28908 4140 28960 4146
rect 28908 4082 28960 4088
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 28816 3392 28868 3398
rect 28816 3334 28868 3340
rect 26516 2984 26568 2990
rect 26516 2926 26568 2932
rect 27528 2984 27580 2990
rect 27528 2926 27580 2932
rect 26528 480 26556 2926
rect 27724 480 27752 3334
rect 28920 480 28948 4082
rect 30116 480 30144 6886
rect 33060 3398 33088 57666
rect 34440 3398 34468 57802
rect 35808 57180 35860 57186
rect 35808 57122 35860 57128
rect 35820 3398 35848 57122
rect 37188 54528 37240 54534
rect 37188 54470 37240 54476
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 34428 3392 34480 3398
rect 34428 3334 34480 3340
rect 34796 3392 34848 3398
rect 34796 3334 34848 3340
rect 35808 3392 35860 3398
rect 35808 3334 35860 3340
rect 31300 3324 31352 3330
rect 31300 3266 31352 3272
rect 31312 480 31340 3266
rect 32416 480 32444 3334
rect 33612 480 33640 3334
rect 34808 480 34836 3334
rect 35992 3120 36044 3126
rect 35992 3062 36044 3068
rect 36004 480 36032 3062
rect 37200 480 37228 54470
rect 39960 6914 39988 57870
rect 41328 57112 41380 57118
rect 41328 57054 41380 57060
rect 39592 6886 39988 6914
rect 38384 3188 38436 3194
rect 38384 3130 38436 3136
rect 38396 480 38424 3130
rect 39592 480 39620 6886
rect 41340 3398 41368 57054
rect 43444 57044 43496 57050
rect 43444 56986 43496 56992
rect 40684 3392 40736 3398
rect 40684 3334 40736 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 43076 3392 43128 3398
rect 43076 3334 43128 3340
rect 40696 480 40724 3334
rect 41880 3256 41932 3262
rect 41880 3198 41932 3204
rect 41892 480 41920 3198
rect 43088 480 43116 3334
rect 43456 3262 43484 56986
rect 46848 56976 46900 56982
rect 46848 56918 46900 56924
rect 45468 54732 45520 54738
rect 45468 54674 45520 54680
rect 45376 54664 45428 54670
rect 45376 54606 45428 54612
rect 44088 54596 44140 54602
rect 44088 54538 44140 54544
rect 44100 3398 44128 54538
rect 44088 3392 44140 3398
rect 44088 3334 44140 3340
rect 43444 3256 43496 3262
rect 43444 3198 43496 3204
rect 45388 3194 45416 54606
rect 44272 3188 44324 3194
rect 44272 3130 44324 3136
rect 45376 3188 45428 3194
rect 45376 3130 45428 3136
rect 44284 480 44312 3130
rect 45480 480 45508 54674
rect 46860 6914 46888 56918
rect 48228 56908 48280 56914
rect 48228 56850 48280 56856
rect 48240 6914 48268 56850
rect 53748 56840 53800 56846
rect 53748 56782 53800 56788
rect 53656 54868 53708 54874
rect 53656 54810 53708 54816
rect 49608 54800 49660 54806
rect 49608 54742 49660 54748
rect 46676 6886 46888 6914
rect 47872 6886 48268 6914
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 49620 3330 49648 54742
rect 53668 4146 53696 54810
rect 52460 4140 52512 4146
rect 52460 4082 52512 4088
rect 52552 4140 52604 4146
rect 52552 4082 52604 4088
rect 53656 4140 53708 4146
rect 53656 4082 53708 4088
rect 52472 3874 52500 4082
rect 52368 3868 52420 3874
rect 52368 3810 52420 3816
rect 52460 3868 52512 3874
rect 52460 3810 52512 3816
rect 48964 3324 49016 3330
rect 48964 3266 49016 3272
rect 49608 3324 49660 3330
rect 49608 3266 49660 3272
rect 48976 480 49004 3266
rect 50160 2984 50212 2990
rect 50160 2926 50212 2932
rect 50172 480 50200 2926
rect 52380 2922 52408 3810
rect 52368 2916 52420 2922
rect 52368 2858 52420 2864
rect 51356 740 51408 746
rect 51356 682 51408 688
rect 51368 480 51396 682
rect 52564 480 52592 4082
rect 53760 480 53788 56782
rect 55128 56772 55180 56778
rect 55128 56714 55180 56720
rect 55140 2774 55168 56714
rect 55784 46238 55812 229094
rect 55876 206281 55904 264794
rect 56048 262812 56100 262818
rect 56048 262754 56100 262760
rect 55954 235376 56010 235385
rect 55954 235311 56010 235320
rect 55862 206272 55918 206281
rect 55862 206207 55918 206216
rect 55968 121281 55996 235311
rect 56060 137057 56088 262754
rect 56140 260704 56192 260710
rect 56140 260646 56192 260652
rect 56046 137048 56102 137057
rect 56046 136983 56102 136992
rect 55954 121272 56010 121281
rect 55954 121207 56010 121216
rect 56152 108769 56180 260646
rect 56230 239592 56286 239601
rect 56230 239527 56286 239536
rect 56138 108760 56194 108769
rect 56138 108695 56194 108704
rect 56244 83609 56272 239527
rect 56336 184249 56364 356662
rect 56414 236600 56470 236609
rect 56414 236535 56470 236544
rect 56428 215801 56456 236535
rect 56414 215792 56470 215801
rect 56414 215727 56470 215736
rect 56322 184240 56378 184249
rect 56322 184175 56378 184184
rect 56520 165345 56548 395354
rect 56506 165336 56562 165345
rect 56506 165271 56562 165280
rect 56612 105641 56640 432239
rect 56782 227216 56838 227225
rect 56782 227151 56838 227160
rect 56690 226672 56746 226681
rect 56690 226607 56746 226616
rect 56598 105632 56654 105641
rect 56598 105567 56654 105576
rect 56230 83600 56286 83609
rect 56230 83535 56286 83544
rect 56704 77217 56732 226607
rect 56796 149705 56824 227151
rect 56782 149696 56838 149705
rect 56782 149631 56838 149640
rect 56690 77208 56746 77217
rect 56690 77143 56746 77152
rect 56888 64705 56916 487319
rect 58438 485344 58494 485353
rect 58438 485279 58494 485288
rect 57518 483984 57574 483993
rect 57518 483919 57574 483928
rect 57334 435432 57390 435441
rect 57334 435367 57390 435376
rect 57242 433392 57298 433401
rect 57242 433327 57298 433336
rect 57150 429448 57206 429457
rect 57150 429383 57206 429392
rect 57058 407552 57114 407561
rect 57058 407487 57114 407496
rect 57072 399702 57100 407487
rect 57060 399696 57112 399702
rect 57060 399638 57112 399644
rect 57164 399566 57192 429383
rect 57256 399634 57284 433327
rect 57244 399628 57296 399634
rect 57244 399570 57296 399576
rect 57152 399560 57204 399566
rect 57152 399502 57204 399508
rect 57348 399498 57376 435367
rect 57426 427952 57482 427961
rect 57426 427887 57482 427896
rect 57336 399492 57388 399498
rect 57336 399434 57388 399440
rect 57242 243672 57298 243681
rect 57242 243607 57298 243616
rect 57150 243536 57206 243545
rect 57150 243471 57206 243480
rect 57058 226264 57114 226273
rect 57058 226199 57114 226208
rect 57072 187513 57100 226199
rect 57058 187504 57114 187513
rect 57058 187439 57114 187448
rect 57164 102377 57192 243471
rect 57150 102368 57206 102377
rect 57150 102303 57206 102312
rect 57256 96121 57284 243607
rect 57334 239456 57390 239465
rect 57334 239391 57390 239400
rect 57242 96112 57298 96121
rect 57242 96047 57298 96056
rect 57348 89865 57376 239391
rect 57440 218074 57468 427887
rect 57532 222057 57560 483919
rect 57794 436384 57850 436393
rect 57794 436319 57850 436328
rect 57610 430672 57666 430681
rect 57610 430607 57666 430616
rect 57518 222048 57574 222057
rect 57518 221983 57574 221992
rect 57428 218068 57480 218074
rect 57428 218010 57480 218016
rect 57520 213920 57572 213926
rect 57520 213862 57572 213868
rect 57532 212673 57560 213862
rect 57518 212664 57574 212673
rect 57518 212599 57574 212608
rect 57520 197328 57572 197334
rect 57520 197270 57572 197276
rect 57532 196897 57560 197270
rect 57518 196888 57574 196897
rect 57518 196823 57574 196832
rect 57520 194540 57572 194546
rect 57520 194482 57572 194488
rect 57532 193769 57560 194482
rect 57518 193760 57574 193769
rect 57518 193695 57574 193704
rect 57520 191820 57572 191826
rect 57520 191762 57572 191768
rect 57532 190641 57560 191762
rect 57518 190632 57574 190641
rect 57518 190567 57574 190576
rect 57520 182164 57572 182170
rect 57520 182106 57572 182112
rect 57532 181121 57560 182106
rect 57518 181112 57574 181121
rect 57518 181047 57574 181056
rect 57520 178016 57572 178022
rect 57518 177984 57520 177993
rect 57572 177984 57574 177993
rect 57518 177919 57574 177928
rect 57520 175228 57572 175234
rect 57520 175170 57572 175176
rect 57532 174865 57560 175170
rect 57518 174856 57574 174865
rect 57518 174791 57574 174800
rect 57428 160064 57480 160070
rect 57428 160006 57480 160012
rect 57440 159089 57468 160006
rect 57426 159080 57482 159089
rect 57426 159015 57482 159024
rect 57518 155952 57574 155961
rect 57518 155887 57520 155896
rect 57572 155887 57574 155896
rect 57520 155858 57572 155864
rect 57520 153196 57572 153202
rect 57520 153138 57572 153144
rect 57532 152833 57560 153138
rect 57518 152824 57574 152833
rect 57518 152759 57574 152768
rect 57428 147620 57480 147626
rect 57428 147562 57480 147568
rect 57440 146577 57468 147562
rect 57426 146568 57482 146577
rect 57426 146503 57482 146512
rect 57520 143540 57572 143546
rect 57520 143482 57572 143488
rect 57532 143313 57560 143482
rect 57518 143304 57574 143313
rect 57518 143239 57574 143248
rect 57520 136604 57572 136610
rect 57520 136546 57572 136552
rect 57428 134768 57480 134774
rect 57428 134710 57480 134716
rect 57440 133929 57468 134710
rect 57426 133920 57482 133929
rect 57426 133855 57482 133864
rect 57532 122834 57560 136546
rect 57624 132494 57652 430607
rect 57624 132466 57744 132494
rect 57612 131096 57664 131102
rect 57612 131038 57664 131044
rect 57624 130801 57652 131038
rect 57610 130792 57666 130801
rect 57610 130727 57666 130736
rect 57716 127974 57744 132466
rect 57704 127968 57756 127974
rect 57704 127910 57756 127916
rect 57440 122806 57560 122834
rect 57334 89856 57390 89865
rect 57334 89791 57390 89800
rect 57440 86737 57468 122806
rect 57612 118652 57664 118658
rect 57612 118594 57664 118600
rect 57624 118153 57652 118594
rect 57610 118144 57666 118153
rect 57610 118079 57666 118088
rect 57612 113144 57664 113150
rect 57612 113086 57664 113092
rect 57624 111897 57652 113086
rect 57610 111888 57666 111897
rect 57610 111823 57666 111832
rect 57704 106276 57756 106282
rect 57704 106218 57756 106224
rect 57426 86728 57482 86737
rect 57426 86663 57482 86672
rect 57716 74089 57744 106218
rect 57702 74080 57758 74089
rect 57702 74015 57758 74024
rect 57612 71732 57664 71738
rect 57612 71674 57664 71680
rect 57624 70961 57652 71674
rect 57610 70952 57666 70961
rect 57610 70887 57666 70896
rect 56874 64696 56930 64705
rect 56874 64631 56930 64640
rect 57060 62076 57112 62082
rect 57060 62018 57112 62024
rect 57072 61577 57100 62018
rect 57058 61568 57114 61577
rect 57058 61503 57114 61512
rect 57808 59362 57836 436319
rect 57886 410000 57942 410009
rect 57886 409935 57942 409944
rect 57900 398138 57928 409935
rect 57888 398132 57940 398138
rect 57888 398074 57940 398080
rect 58346 250472 58402 250481
rect 58346 250407 58402 250416
rect 58254 240816 58310 240825
rect 58254 240751 58310 240760
rect 58070 238096 58126 238105
rect 58070 238031 58126 238040
rect 57886 226400 57942 226409
rect 57886 226335 57942 226344
rect 57900 209545 57928 226335
rect 57886 209536 57942 209545
rect 57886 209471 57942 209480
rect 58084 162217 58112 238031
rect 58162 235240 58218 235249
rect 58162 235175 58218 235184
rect 58176 218929 58204 235175
rect 58162 218920 58218 218929
rect 58162 218855 58218 218864
rect 58070 162208 58126 162217
rect 58070 162143 58126 162152
rect 58268 124545 58296 240751
rect 58254 124536 58310 124545
rect 58254 124471 58310 124480
rect 58360 115025 58388 250407
rect 58452 229945 58480 485279
rect 58530 485208 58586 485217
rect 58530 485143 58586 485152
rect 58544 230081 58572 485143
rect 58624 396636 58676 396642
rect 58624 396578 58676 396584
rect 58530 230072 58586 230081
rect 58530 230007 58586 230016
rect 58438 229936 58494 229945
rect 58438 229871 58494 229880
rect 58532 218068 58584 218074
rect 58532 218010 58584 218016
rect 58346 115016 58402 115025
rect 58346 114951 58402 114960
rect 57796 59356 57848 59362
rect 57796 59298 57848 59304
rect 57796 57384 57848 57390
rect 57624 57332 57796 57338
rect 57624 57326 57848 57332
rect 57624 57322 57836 57326
rect 57612 57316 57836 57322
rect 57664 57310 57836 57316
rect 57612 57258 57664 57264
rect 58544 57089 58572 218010
rect 58636 140185 58664 396578
rect 58728 200025 58756 487591
rect 58714 200016 58770 200025
rect 58714 199951 58770 199960
rect 58820 168609 58848 487863
rect 58912 399838 58940 700266
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 88340 699712 88392 699718
rect 88340 699654 88392 699660
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 104900 699712 104952 699718
rect 104900 699654 104952 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 77208 647896 77260 647902
rect 77208 647838 77260 647844
rect 77220 645930 77248 647838
rect 74540 645924 74592 645930
rect 74540 645866 74592 645872
rect 77208 645924 77260 645930
rect 77208 645866 77260 645872
rect 74552 638994 74580 645866
rect 74540 638988 74592 638994
rect 74540 638930 74592 638936
rect 71780 638920 71832 638926
rect 71780 638862 71832 638868
rect 71792 636274 71820 638862
rect 71780 636268 71832 636274
rect 71780 636210 71832 636216
rect 69020 636200 69072 636206
rect 69020 636142 69072 636148
rect 69032 632126 69060 636142
rect 69020 632120 69072 632126
rect 69020 632062 69072 632068
rect 65524 632052 65576 632058
rect 65524 631994 65576 632000
rect 65536 604518 65564 631994
rect 64144 604512 64196 604518
rect 64144 604454 64196 604460
rect 65524 604512 65576 604518
rect 65524 604454 65576 604460
rect 64156 572762 64184 604454
rect 62764 572756 62816 572762
rect 62764 572698 62816 572704
rect 64144 572756 64196 572762
rect 64144 572698 64196 572704
rect 62776 561066 62804 572698
rect 61384 561060 61436 561066
rect 61384 561002 61436 561008
rect 62764 561060 62816 561066
rect 62764 561002 62816 561008
rect 61396 553450 61424 561002
rect 60004 553444 60056 553450
rect 60004 553386 60056 553392
rect 61384 553444 61436 553450
rect 61384 553386 61436 553392
rect 59082 489968 59138 489977
rect 59082 489903 59138 489912
rect 58990 484664 59046 484673
rect 58990 484599 59046 484608
rect 58900 399832 58952 399838
rect 58900 399774 58952 399780
rect 58900 396228 58952 396234
rect 58900 396170 58952 396176
rect 58806 168600 58862 168609
rect 58806 168535 58862 168544
rect 58622 140176 58678 140185
rect 58622 140111 58678 140120
rect 58716 127968 58768 127974
rect 58716 127910 58768 127916
rect 58728 57905 58756 127910
rect 58912 67833 58940 396170
rect 59004 127673 59032 484599
rect 58990 127664 59046 127673
rect 58990 127599 59046 127608
rect 59096 99249 59124 489903
rect 59266 489016 59322 489025
rect 59266 488951 59322 488960
rect 59174 488880 59230 488889
rect 59174 488815 59230 488824
rect 59082 99240 59138 99249
rect 59082 99175 59138 99184
rect 59188 92993 59216 488815
rect 59174 92984 59230 92993
rect 59174 92919 59230 92928
rect 59280 80345 59308 488951
rect 59358 408232 59414 408241
rect 59358 408167 59414 408176
rect 59372 398818 59400 408167
rect 60016 398886 60044 553386
rect 88352 485353 88380 699654
rect 104256 674756 104308 674762
rect 104256 674698 104308 674704
rect 104268 667418 104296 674698
rect 102784 667412 102836 667418
rect 102784 667354 102836 667360
rect 104256 667412 104308 667418
rect 104256 667354 104308 667360
rect 102796 662454 102824 667354
rect 100760 662448 100812 662454
rect 100760 662390 100812 662396
rect 102784 662448 102836 662454
rect 102784 662390 102836 662396
rect 100772 659734 100800 662390
rect 100760 659728 100812 659734
rect 100760 659670 100812 659676
rect 96528 659660 96580 659666
rect 96528 659602 96580 659608
rect 96540 658034 96568 659602
rect 94504 658028 94556 658034
rect 94504 657970 94556 657976
rect 96528 658028 96580 658034
rect 96528 657970 96580 657976
rect 94516 650146 94544 657970
rect 92480 650140 92532 650146
rect 92480 650082 92532 650088
rect 94504 650140 94556 650146
rect 94504 650082 94556 650088
rect 92492 647902 92520 650082
rect 92480 647896 92532 647902
rect 92480 647838 92532 647844
rect 88338 485344 88394 485353
rect 88338 485279 88394 485288
rect 104912 485217 104940 699654
rect 137848 698630 137876 703520
rect 154132 700330 154160 703520
rect 170324 700398 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 170312 700392 170364 700398
rect 170312 700334 170364 700340
rect 196532 700392 196584 700398
rect 196532 700334 196584 700340
rect 154120 700324 154172 700330
rect 154120 700266 154172 700272
rect 134156 698624 134208 698630
rect 134156 698566 134208 698572
rect 137836 698624 137888 698630
rect 137836 698566 137888 698572
rect 134168 696998 134196 698566
rect 134156 696992 134208 696998
rect 134156 696934 134208 696940
rect 128912 696924 128964 696930
rect 128912 696866 128964 696872
rect 128924 693802 128952 696866
rect 126520 693796 126572 693802
rect 126520 693738 126572 693744
rect 128912 693796 128964 693802
rect 128912 693738 128964 693744
rect 126532 690198 126560 693738
rect 124588 690192 124640 690198
rect 124588 690134 124640 690140
rect 126520 690192 126572 690198
rect 126520 690134 126572 690140
rect 124600 688702 124628 690134
rect 121460 688696 121512 688702
rect 121460 688638 121512 688644
rect 124588 688696 124640 688702
rect 124588 688638 124640 688644
rect 121472 684418 121500 688638
rect 114560 684412 114612 684418
rect 114560 684354 114612 684360
rect 121460 684412 121512 684418
rect 121460 684354 121512 684360
rect 114572 681766 114600 684354
rect 114560 681760 114612 681766
rect 114560 681702 114612 681708
rect 106280 681692 106332 681698
rect 106280 681634 106332 681640
rect 106292 677634 106320 681634
rect 106200 677606 106320 677634
rect 106200 674762 106228 677606
rect 106188 674756 106240 674762
rect 106188 674698 106240 674704
rect 118606 490104 118662 490113
rect 118606 490039 118662 490048
rect 118620 486441 118648 490039
rect 158534 488064 158590 488073
rect 158534 487999 158590 488008
rect 133602 487928 133658 487937
rect 133602 487863 133658 487872
rect 118606 486432 118662 486441
rect 118606 486367 118662 486376
rect 133616 485897 133644 487863
rect 138570 487792 138626 487801
rect 138570 487727 138626 487736
rect 143722 487792 143778 487801
rect 143722 487727 143778 487736
rect 138584 485897 138612 487727
rect 143736 485897 143764 487727
rect 153934 487656 153990 487665
rect 153934 487591 153990 487600
rect 153948 485897 153976 487591
rect 158548 485897 158576 487999
rect 133602 485888 133658 485897
rect 133602 485823 133658 485832
rect 138570 485888 138626 485897
rect 138570 485823 138626 485832
rect 143722 485888 143778 485897
rect 143722 485823 143778 485832
rect 153934 485888 153990 485897
rect 153934 485823 153990 485832
rect 158534 485888 158590 485897
rect 158534 485823 158590 485832
rect 104898 485208 104954 485217
rect 104898 485143 104954 485152
rect 121460 399832 121512 399838
rect 121460 399774 121512 399780
rect 177948 399832 178000 399838
rect 177948 399774 178000 399780
rect 111708 399764 111760 399770
rect 111708 399706 111760 399712
rect 60004 398880 60056 398886
rect 60004 398822 60056 398828
rect 62028 398880 62080 398886
rect 62028 398822 62080 398828
rect 59360 398812 59412 398818
rect 59360 398754 59412 398760
rect 59266 80336 59322 80345
rect 59266 80271 59322 80280
rect 59372 74534 59400 398754
rect 62040 397338 62068 398822
rect 85486 398168 85542 398177
rect 85486 398103 85542 398112
rect 92294 398168 92350 398177
rect 92294 398103 92350 398112
rect 95882 398168 95938 398177
rect 95882 398103 95938 398112
rect 76194 397352 76250 397361
rect 62040 397310 62160 397338
rect 61476 396976 61528 396982
rect 61476 396918 61528 396924
rect 61384 396568 61436 396574
rect 61384 396510 61436 396516
rect 60004 396364 60056 396370
rect 60004 396306 60056 396312
rect 59912 396160 59964 396166
rect 59912 396102 59964 396108
rect 59544 264444 59596 264450
rect 59544 264386 59596 264392
rect 59452 262064 59504 262070
rect 59452 262006 59504 262012
rect 59464 171737 59492 262006
rect 59556 203153 59584 264386
rect 59820 229152 59872 229158
rect 59820 229094 59872 229100
rect 59832 226817 59860 229094
rect 59818 226808 59874 226817
rect 59818 226743 59874 226752
rect 59542 203144 59598 203153
rect 59542 203079 59598 203088
rect 59450 171728 59506 171737
rect 59450 171663 59506 171672
rect 59924 142154 59952 396102
rect 59832 142126 59952 142154
rect 59832 136610 59860 142126
rect 59820 136604 59872 136610
rect 59820 136546 59872 136552
rect 60016 113174 60044 396306
rect 61396 227225 61424 396510
rect 61382 227216 61438 227225
rect 61382 227151 61438 227160
rect 61488 227066 61516 396918
rect 61568 395480 61620 395486
rect 61568 395422 61620 395428
rect 61580 229094 61608 395422
rect 62132 394738 62160 397310
rect 76194 397287 76250 397296
rect 78310 397352 78366 397361
rect 78310 397287 78366 397296
rect 79598 397352 79654 397361
rect 79598 397287 79654 397296
rect 80426 397352 80482 397361
rect 80426 397287 80482 397296
rect 82358 397352 82414 397361
rect 82358 397287 82414 397296
rect 83002 397352 83058 397361
rect 85500 397322 85528 398103
rect 89350 397352 89406 397361
rect 83002 397287 83058 397296
rect 85488 397316 85540 397322
rect 62948 397248 63000 397254
rect 62948 397190 63000 397196
rect 62764 397044 62816 397050
rect 62764 396986 62816 396992
rect 62120 394732 62172 394738
rect 62120 394674 62172 394680
rect 61580 229066 62068 229094
rect 61120 227038 61516 227066
rect 60186 226808 60242 226817
rect 60242 226766 60490 226794
rect 60186 226743 60242 226752
rect 61120 226273 61148 227038
rect 61750 226536 61806 226545
rect 61410 226494 61750 226522
rect 61750 226471 61806 226480
rect 62040 226273 62068 229066
rect 62670 226808 62726 226817
rect 62330 226766 62670 226794
rect 62670 226743 62726 226752
rect 62776 226409 62804 396986
rect 62960 226681 62988 397190
rect 76208 396370 76236 397287
rect 78324 396846 78352 397287
rect 79612 397186 79640 397287
rect 79600 397180 79652 397186
rect 79600 397122 79652 397128
rect 78312 396840 78364 396846
rect 77206 396808 77262 396817
rect 78312 396782 78364 396788
rect 77206 396743 77262 396752
rect 76196 396364 76248 396370
rect 76196 396306 76248 396312
rect 66260 394664 66312 394670
rect 66260 394606 66312 394612
rect 66272 389230 66300 394606
rect 66260 389224 66312 389230
rect 66260 389166 66312 389172
rect 68284 389224 68336 389230
rect 68284 389166 68336 389172
rect 68296 378146 68324 389166
rect 68284 378140 68336 378146
rect 68284 378082 68336 378088
rect 69664 378140 69716 378146
rect 69664 378082 69716 378088
rect 69676 372910 69704 378082
rect 69664 372904 69716 372910
rect 69664 372846 69716 372852
rect 70400 372904 70452 372910
rect 70400 372846 70452 372852
rect 70412 369850 70440 372846
rect 70400 369844 70452 369850
rect 70400 369786 70452 369792
rect 75184 369844 75236 369850
rect 75184 369786 75236 369792
rect 75196 358766 75224 369786
rect 75184 358760 75236 358766
rect 75184 358702 75236 358708
rect 76656 358760 76708 358766
rect 76656 358702 76708 358708
rect 76668 357406 76696 358702
rect 76656 357400 76708 357406
rect 76656 357342 76708 357348
rect 77220 267034 77248 396743
rect 80440 396166 80468 397287
rect 82372 396914 82400 397287
rect 82360 396908 82412 396914
rect 82360 396850 82412 396856
rect 83016 396234 83044 397287
rect 89350 397287 89406 397296
rect 90086 397352 90142 397361
rect 90086 397287 90142 397296
rect 91466 397352 91522 397361
rect 91466 397287 91522 397296
rect 85488 397258 85540 397264
rect 89364 397118 89392 397287
rect 89352 397112 89404 397118
rect 89352 397054 89404 397060
rect 85394 396808 85450 396817
rect 85394 396743 85450 396752
rect 86866 396808 86922 396817
rect 86866 396743 86922 396752
rect 88246 396808 88302 396817
rect 88246 396743 88302 396752
rect 89534 396808 89590 396817
rect 89534 396743 89590 396752
rect 83004 396228 83056 396234
rect 83004 396170 83056 396176
rect 80428 396160 80480 396166
rect 80428 396102 80480 396108
rect 84108 378208 84160 378214
rect 84108 378150 84160 378156
rect 78036 357400 78088 357406
rect 78036 357342 78088 357348
rect 78048 353326 78076 357342
rect 78036 353320 78088 353326
rect 78036 353262 78088 353268
rect 80704 353320 80756 353326
rect 80704 353262 80756 353268
rect 80716 336054 80744 353262
rect 82728 351960 82780 351966
rect 82728 351902 82780 351908
rect 80704 336048 80756 336054
rect 80704 335990 80756 335996
rect 81348 324352 81400 324358
rect 81348 324294 81400 324300
rect 79968 298172 80020 298178
rect 79968 298114 80020 298120
rect 78588 271924 78640 271930
rect 78588 271866 78640 271872
rect 77208 267028 77260 267034
rect 77208 266970 77260 266976
rect 77206 245712 77262 245721
rect 77206 245647 77262 245656
rect 67362 234696 67418 234705
rect 67362 234631 67418 234640
rect 65982 230752 66038 230761
rect 65982 230687 66038 230696
rect 63222 229800 63278 229809
rect 63222 229735 63278 229744
rect 63236 226780 63264 229735
rect 64142 229392 64198 229401
rect 64142 229327 64198 229336
rect 64156 226780 64184 229327
rect 65062 227896 65118 227905
rect 65062 227831 65118 227840
rect 65076 226780 65104 227831
rect 65996 226780 66024 230687
rect 67376 226794 67404 234631
rect 75642 231976 75698 231985
rect 75642 231911 75698 231920
rect 68742 230888 68798 230897
rect 68742 230823 68798 230832
rect 66930 226766 67404 226794
rect 68756 226780 68784 230823
rect 70398 230616 70454 230625
rect 70398 230551 70454 230560
rect 70412 229809 70440 230551
rect 70398 229800 70454 229809
rect 70398 229735 70454 229744
rect 74538 229800 74594 229809
rect 74538 229735 74594 229744
rect 70306 229664 70362 229673
rect 70306 229599 70362 229608
rect 70320 227089 70348 229599
rect 71686 229528 71742 229537
rect 71686 229463 71742 229472
rect 71700 228585 71728 229463
rect 71686 228576 71742 228585
rect 71686 228511 71742 228520
rect 74552 228449 74580 229735
rect 74538 228440 74594 228449
rect 74538 228375 74594 228384
rect 73342 228168 73398 228177
rect 73342 228103 73398 228112
rect 70582 228032 70638 228041
rect 70582 227967 70638 227976
rect 70306 227080 70362 227089
rect 70306 227015 70362 227024
rect 70030 226944 70086 226953
rect 70030 226879 70086 226888
rect 70044 226794 70072 226879
rect 69690 226766 70072 226794
rect 70596 226780 70624 227967
rect 72422 227760 72478 227769
rect 72422 227695 72478 227704
rect 72436 226780 72464 227695
rect 73356 226780 73384 228103
rect 74262 227080 74318 227089
rect 74262 227015 74318 227024
rect 74276 226780 74304 227015
rect 75656 226794 75684 231911
rect 76194 228440 76250 228449
rect 76194 228375 76250 228384
rect 75210 226766 75684 226794
rect 76208 226780 76236 228375
rect 77220 226794 77248 245647
rect 78600 229094 78628 271866
rect 79322 237960 79378 237969
rect 79322 237895 79378 237904
rect 78416 229066 78628 229094
rect 78416 226794 78444 229066
rect 79336 226794 79364 237895
rect 79980 226794 80008 298114
rect 81360 234614 81388 324294
rect 82636 311908 82688 311914
rect 82636 311850 82688 311856
rect 82648 234614 82676 311850
rect 81176 234586 81388 234614
rect 82096 234586 82676 234614
rect 81176 226794 81204 234586
rect 82096 226794 82124 234586
rect 82740 226794 82768 351902
rect 84120 234614 84148 378150
rect 84200 336048 84252 336054
rect 84200 335990 84252 335996
rect 84212 329798 84240 335990
rect 84200 329792 84252 329798
rect 84200 329734 84252 329740
rect 85408 266014 85436 396743
rect 85488 364404 85540 364410
rect 85488 364346 85540 364352
rect 85396 266008 85448 266014
rect 85396 265950 85448 265956
rect 85396 260228 85448 260234
rect 85396 260170 85448 260176
rect 85408 234614 85436 260170
rect 83936 234586 84148 234614
rect 85316 234586 85436 234614
rect 83936 226794 83964 234586
rect 84474 228984 84530 228993
rect 84474 228919 84530 228928
rect 77142 226766 77248 226794
rect 78062 226766 78444 226794
rect 78982 226766 79364 226794
rect 79902 226766 80008 226794
rect 80822 226766 81204 226794
rect 81742 226766 82124 226794
rect 82662 226766 82768 226794
rect 83582 226766 83964 226794
rect 84488 226780 84516 228919
rect 85316 226794 85344 234586
rect 85500 228993 85528 364346
rect 86224 329792 86276 329798
rect 86224 329734 86276 329740
rect 86236 324630 86264 329734
rect 86224 324624 86276 324630
rect 86224 324566 86276 324572
rect 86880 266082 86908 396743
rect 87972 324624 88024 324630
rect 87972 324566 88024 324572
rect 87984 322998 88012 324566
rect 87972 322992 88024 322998
rect 87972 322934 88024 322940
rect 86868 266076 86920 266082
rect 86868 266018 86920 266024
rect 88260 265946 88288 396743
rect 88248 265940 88300 265946
rect 88248 265882 88300 265888
rect 88248 265668 88300 265674
rect 88248 265610 88300 265616
rect 86868 262948 86920 262954
rect 86868 262890 86920 262896
rect 86880 234614 86908 262890
rect 88156 260160 88208 260166
rect 88156 260102 88208 260108
rect 88168 234614 88196 260102
rect 86696 234586 86908 234614
rect 88076 234586 88196 234614
rect 85486 228984 85542 228993
rect 85486 228919 85542 228928
rect 86696 226794 86724 234586
rect 87234 228984 87290 228993
rect 87234 228919 87290 228928
rect 85316 226766 85422 226794
rect 86342 226766 86724 226794
rect 87248 226780 87276 228919
rect 88076 226794 88104 234586
rect 88260 228993 88288 265610
rect 89548 263838 89576 396743
rect 90100 396438 90128 397287
rect 90914 396808 90970 396817
rect 90914 396743 90970 396752
rect 90088 396432 90140 396438
rect 90088 396374 90140 396380
rect 90928 264518 90956 396743
rect 91480 396370 91508 397287
rect 91468 396364 91520 396370
rect 91468 396306 91520 396312
rect 91744 322924 91796 322930
rect 91744 322866 91796 322872
rect 91756 314294 91784 322866
rect 91744 314288 91796 314294
rect 91744 314230 91796 314236
rect 92308 266150 92336 398103
rect 93490 397352 93546 397361
rect 93490 397287 93546 397296
rect 95054 397352 95110 397361
rect 95054 397287 95110 397296
rect 92478 396808 92534 396817
rect 92478 396743 92534 396752
rect 92296 266144 92348 266150
rect 92296 266086 92348 266092
rect 90916 264512 90968 264518
rect 90916 264454 90968 264460
rect 89536 263832 89588 263838
rect 89536 263774 89588 263780
rect 91008 263084 91060 263090
rect 91008 263026 91060 263032
rect 89628 261724 89680 261730
rect 89628 261666 89680 261672
rect 89640 234614 89668 261666
rect 90916 260568 90968 260574
rect 90916 260510 90968 260516
rect 90928 234614 90956 260510
rect 89456 234586 89668 234614
rect 90836 234586 90956 234614
rect 88246 228984 88302 228993
rect 88246 228919 88302 228928
rect 89456 226794 89484 234586
rect 90270 230480 90326 230489
rect 90270 230415 90326 230424
rect 90284 226794 90312 230415
rect 88076 226766 88182 226794
rect 89102 226766 89484 226794
rect 90022 226766 90312 226794
rect 90836 226794 90864 234586
rect 91020 230489 91048 263026
rect 92388 261792 92440 261798
rect 92388 261734 92440 261740
rect 91006 230480 91062 230489
rect 91006 230415 91062 230424
rect 92400 226794 92428 261734
rect 92492 239601 92520 396743
rect 93504 396302 93532 397287
rect 94504 397112 94556 397118
rect 94504 397054 94556 397060
rect 93492 396296 93544 396302
rect 93492 396238 93544 396244
rect 94516 265538 94544 397054
rect 95068 396506 95096 397287
rect 95896 396642 95924 398103
rect 98090 397352 98146 397361
rect 98090 397287 98146 397296
rect 102782 397352 102838 397361
rect 102782 397287 102838 397296
rect 104806 397352 104862 397361
rect 104806 397287 104862 397296
rect 106094 397352 106150 397361
rect 106094 397287 106150 397296
rect 106922 397352 106978 397361
rect 106922 397287 106978 397296
rect 108854 397352 108910 397361
rect 108854 397287 108910 397296
rect 109130 397352 109186 397361
rect 109130 397287 109186 397296
rect 96526 396808 96582 396817
rect 96526 396743 96582 396752
rect 97906 396808 97962 396817
rect 97906 396743 97962 396752
rect 95884 396636 95936 396642
rect 95884 396578 95936 396584
rect 95056 396500 95108 396506
rect 95056 396442 95108 396448
rect 94596 314288 94648 314294
rect 94596 314230 94648 314236
rect 94608 295390 94636 314230
rect 94596 295384 94648 295390
rect 94596 295326 94648 295332
rect 94504 265532 94556 265538
rect 94504 265474 94556 265480
rect 93768 263016 93820 263022
rect 93768 262958 93820 262964
rect 93676 260364 93728 260370
rect 93676 260306 93728 260312
rect 92478 239592 92534 239601
rect 92478 239527 92534 239536
rect 93688 234614 93716 260306
rect 93596 234586 93716 234614
rect 93214 230480 93270 230489
rect 93214 230415 93270 230424
rect 93228 226794 93256 230415
rect 90836 226766 91034 226794
rect 91954 226766 92428 226794
rect 92874 226766 93256 226794
rect 93596 226794 93624 234586
rect 93780 230489 93808 262958
rect 96436 261656 96488 261662
rect 96436 261598 96488 261604
rect 95148 261520 95200 261526
rect 95148 261462 95200 261468
rect 93766 230480 93822 230489
rect 93766 230415 93822 230424
rect 95160 226794 95188 261462
rect 96344 260296 96396 260302
rect 96344 260238 96396 260244
rect 95606 228984 95662 228993
rect 95606 228919 95662 228928
rect 93596 226766 93794 226794
rect 94714 226766 95188 226794
rect 95620 226780 95648 228919
rect 96356 226794 96384 260238
rect 96448 228993 96476 261598
rect 96540 234025 96568 396743
rect 97264 295384 97316 295390
rect 97264 295326 97316 295332
rect 97276 282946 97304 295326
rect 97264 282940 97316 282946
rect 97264 282882 97316 282888
rect 97816 263288 97868 263294
rect 97816 263230 97868 263236
rect 96526 234016 96582 234025
rect 96526 233951 96582 233960
rect 96434 228984 96490 228993
rect 96434 228919 96490 228928
rect 97828 226794 97856 263230
rect 97920 262138 97948 396743
rect 98104 396574 98132 397287
rect 101954 396944 102010 396953
rect 101954 396879 102010 396888
rect 99286 396808 99342 396817
rect 99286 396743 99342 396752
rect 100666 396808 100722 396817
rect 100666 396743 100722 396752
rect 98092 396568 98144 396574
rect 98092 396510 98144 396516
rect 99300 263566 99328 396743
rect 99472 282872 99524 282878
rect 99472 282814 99524 282820
rect 99484 278730 99512 282814
rect 99472 278724 99524 278730
rect 99472 278666 99524 278672
rect 100680 264586 100708 396743
rect 100758 396672 100814 396681
rect 100758 396607 100814 396616
rect 100668 264580 100720 264586
rect 100668 264522 100720 264528
rect 99288 263560 99340 263566
rect 99288 263502 99340 263508
rect 99288 263152 99340 263158
rect 99288 263094 99340 263100
rect 97908 262132 97960 262138
rect 97908 262074 97960 262080
rect 99196 260432 99248 260438
rect 99196 260374 99248 260380
rect 99208 234614 99236 260374
rect 99116 234586 99236 234614
rect 98734 230480 98790 230489
rect 98734 230415 98790 230424
rect 98748 226794 98776 230415
rect 96356 226766 96554 226794
rect 97474 226766 97856 226794
rect 98394 226766 98776 226794
rect 99116 226794 99144 234586
rect 99300 230489 99328 263094
rect 100668 261860 100720 261866
rect 100668 261802 100720 261808
rect 99286 230480 99342 230489
rect 99286 230415 99342 230424
rect 100680 226794 100708 261802
rect 100772 238105 100800 396607
rect 101496 278724 101548 278730
rect 101496 278666 101548 278672
rect 101508 275262 101536 278666
rect 101496 275256 101548 275262
rect 101496 275198 101548 275204
rect 101968 266286 101996 396879
rect 102046 396808 102102 396817
rect 102046 396743 102102 396752
rect 101956 266280 102008 266286
rect 101956 266222 102008 266228
rect 101956 263220 102008 263226
rect 101956 263162 102008 263168
rect 101864 261996 101916 262002
rect 101864 261938 101916 261944
rect 101876 246401 101904 261938
rect 101862 246392 101918 246401
rect 101862 246327 101918 246336
rect 101968 244066 101996 263162
rect 102060 260506 102088 396743
rect 102796 396098 102824 397287
rect 103518 396808 103574 396817
rect 103518 396743 103574 396752
rect 102784 396092 102836 396098
rect 102784 396034 102836 396040
rect 102140 275256 102192 275262
rect 102140 275198 102192 275204
rect 102152 269142 102180 275198
rect 102140 269136 102192 269142
rect 102140 269078 102192 269084
rect 103428 263356 103480 263362
rect 103428 263298 103480 263304
rect 102048 260500 102100 260506
rect 102048 260442 102100 260448
rect 102046 246392 102102 246401
rect 102046 246327 102102 246336
rect 101876 244038 101996 244066
rect 101876 241514 101904 244038
rect 101876 241486 101996 241514
rect 100758 238096 100814 238105
rect 100758 238031 100814 238040
rect 101968 227066 101996 241486
rect 101600 227038 101996 227066
rect 101600 226794 101628 227038
rect 99116 226766 99314 226794
rect 100234 226766 100708 226794
rect 101154 226766 101628 226794
rect 102060 226780 102088 246327
rect 103440 226794 103468 263298
rect 103532 260710 103560 396743
rect 104820 396574 104848 397287
rect 106002 396808 106058 396817
rect 106002 396743 106058 396752
rect 104808 396568 104860 396574
rect 104808 396510 104860 396516
rect 104164 269136 104216 269142
rect 104164 269078 104216 269084
rect 104176 260846 104204 269078
rect 104808 264240 104860 264246
rect 104808 264182 104860 264188
rect 104716 261928 104768 261934
rect 104716 261870 104768 261876
rect 104164 260840 104216 260846
rect 104164 260782 104216 260788
rect 103520 260704 103572 260710
rect 103520 260646 103572 260652
rect 104728 234614 104756 261870
rect 104636 234586 104756 234614
rect 104254 230480 104310 230489
rect 104254 230415 104310 230424
rect 104268 226794 104296 230415
rect 102994 226766 103468 226794
rect 103914 226766 104296 226794
rect 104636 226794 104664 234586
rect 104820 230489 104848 264182
rect 106016 240961 106044 396743
rect 106108 396166 106136 397287
rect 106936 396642 106964 397287
rect 107474 396808 107530 396817
rect 107474 396743 107530 396752
rect 106924 396636 106976 396642
rect 106924 396578 106976 396584
rect 106096 396160 106148 396166
rect 106096 396102 106148 396108
rect 106924 396092 106976 396098
rect 106924 396034 106976 396040
rect 106936 266354 106964 396034
rect 106924 266348 106976 266354
rect 106924 266290 106976 266296
rect 107488 266218 107516 396743
rect 107658 396672 107714 396681
rect 107658 396607 107714 396616
rect 107476 266212 107528 266218
rect 107476 266154 107528 266160
rect 107568 264308 107620 264314
rect 107568 264250 107620 264256
rect 106096 263424 106148 263430
rect 106096 263366 106148 263372
rect 106002 240952 106058 240961
rect 106002 240887 106058 240896
rect 104806 230480 104862 230489
rect 104806 230415 104862 230424
rect 106108 226794 106136 263366
rect 106648 260840 106700 260846
rect 106648 260782 106700 260788
rect 106660 254017 106688 260782
rect 106646 254008 106702 254017
rect 106646 253943 106702 253952
rect 107580 234614 107608 264250
rect 107672 235385 107700 396607
rect 108868 396098 108896 397287
rect 109144 396982 109172 397287
rect 109132 396976 109184 396982
rect 109132 396918 109184 396924
rect 111614 396808 111670 396817
rect 111614 396743 111670 396752
rect 111522 396672 111578 396681
rect 111522 396607 111578 396616
rect 108856 396092 108908 396098
rect 108856 396034 108908 396040
rect 111536 264654 111564 396607
rect 111524 264648 111576 264654
rect 111524 264590 111576 264596
rect 108948 263492 109000 263498
rect 108948 263434 109000 263440
rect 108856 261588 108908 261594
rect 108856 261530 108908 261536
rect 107658 235376 107714 235385
rect 107658 235311 107714 235320
rect 108868 234614 108896 261530
rect 107120 234586 107608 234614
rect 108040 234586 108896 234614
rect 107120 226794 107148 234586
rect 108040 226794 108068 234586
rect 108960 226794 108988 263434
rect 110328 262880 110380 262886
rect 110328 262822 110380 262828
rect 110340 229094 110368 262822
rect 111524 260976 111576 260982
rect 111524 260918 111576 260924
rect 110418 253872 110474 253881
rect 110418 253807 110474 253816
rect 110432 251841 110460 253807
rect 110418 251832 110474 251841
rect 110418 251767 110474 251776
rect 111536 229094 111564 260918
rect 111628 239601 111656 396743
rect 111614 239592 111670 239601
rect 111614 239527 111670 239536
rect 109880 229066 110368 229094
rect 110800 229066 111564 229094
rect 109880 226794 109908 229066
rect 110800 226794 110828 229066
rect 111720 226794 111748 399706
rect 121368 398268 121420 398274
rect 121368 398210 121420 398216
rect 115848 398200 115900 398206
rect 113638 398168 113694 398177
rect 115848 398142 115900 398148
rect 113638 398103 113694 398112
rect 112350 397352 112406 397361
rect 112350 397287 112406 397296
rect 113362 397352 113418 397361
rect 113362 397287 113418 397296
rect 112364 396710 112392 397287
rect 113376 396778 113404 397287
rect 113364 396772 113416 396778
rect 113364 396714 113416 396720
rect 112352 396704 112404 396710
rect 112352 396646 112404 396652
rect 113652 395894 113680 398103
rect 113822 397352 113878 397361
rect 113822 397287 113878 397296
rect 113836 397050 113864 397287
rect 113824 397044 113876 397050
rect 113824 396986 113876 396992
rect 115754 396808 115810 396817
rect 115754 396743 115810 396752
rect 115204 396160 115256 396166
rect 115204 396102 115256 396108
rect 113640 395888 113692 395894
rect 113640 395830 113692 395836
rect 113088 305652 113140 305658
rect 113088 305594 113140 305600
rect 113100 229094 113128 305594
rect 115216 265606 115244 396102
rect 115204 265600 115256 265606
rect 115204 265542 115256 265548
rect 114468 260772 114520 260778
rect 114468 260714 114520 260720
rect 114376 260704 114428 260710
rect 114376 260646 114428 260652
rect 112640 229066 113128 229094
rect 112640 226794 112668 229066
rect 113454 227624 113510 227633
rect 113454 227559 113510 227568
rect 113468 226794 113496 227559
rect 114388 226794 114416 260646
rect 114480 227633 114508 260714
rect 115768 236881 115796 396743
rect 115754 236872 115810 236881
rect 115754 236807 115810 236816
rect 115860 229094 115888 398142
rect 118238 397352 118294 397361
rect 118238 397287 118294 397296
rect 118606 397352 118662 397361
rect 118606 397287 118662 397296
rect 117226 396808 117282 396817
rect 117226 396743 117282 396752
rect 115938 396672 115994 396681
rect 115938 396607 115994 396616
rect 115952 262818 115980 396607
rect 117240 262818 117268 396743
rect 118252 395554 118280 397287
rect 118620 395962 118648 397287
rect 119986 396808 120042 396817
rect 119986 396743 120042 396752
rect 121274 396808 121330 396817
rect 121274 396743 121330 396752
rect 119344 396092 119396 396098
rect 119344 396034 119396 396040
rect 118608 395956 118660 395962
rect 118608 395898 118660 395904
rect 118240 395548 118292 395554
rect 118240 395490 118292 395496
rect 119356 263974 119384 396034
rect 120000 264790 120028 396743
rect 119988 264784 120040 264790
rect 119988 264726 120040 264732
rect 119344 263968 119396 263974
rect 119344 263910 119396 263916
rect 119988 263900 120040 263906
rect 119988 263842 120040 263848
rect 115940 262812 115992 262818
rect 115940 262754 115992 262760
rect 117228 262812 117280 262818
rect 117228 262754 117280 262760
rect 117228 262472 117280 262478
rect 117228 262414 117280 262420
rect 117136 261112 117188 261118
rect 117136 261054 117188 261060
rect 117148 229094 117176 261054
rect 115400 229066 115888 229094
rect 116320 229066 117176 229094
rect 114466 227624 114522 227633
rect 114466 227559 114522 227568
rect 115400 226794 115428 229066
rect 116320 226794 116348 229066
rect 117240 226794 117268 262414
rect 118608 261044 118660 261050
rect 118608 260986 118660 260992
rect 118620 229094 118648 260986
rect 118698 251832 118754 251841
rect 118698 251767 118754 251776
rect 118712 248414 118740 251767
rect 118712 248386 119200 248414
rect 118160 229066 118648 229094
rect 118160 226794 118188 229066
rect 118974 227624 119030 227633
rect 118974 227559 119030 227568
rect 118988 226794 119016 227559
rect 104636 226766 104834 226794
rect 105846 226766 106136 226794
rect 106766 226766 107148 226794
rect 107686 226766 108068 226794
rect 108606 226766 108988 226794
rect 109526 226766 109908 226794
rect 110446 226766 110828 226794
rect 111366 226766 111748 226794
rect 112286 226766 112668 226794
rect 113206 226766 113496 226794
rect 114126 226766 114416 226794
rect 115046 226766 115428 226794
rect 115966 226766 116348 226794
rect 116886 226766 117268 226794
rect 117806 226766 118188 226794
rect 118726 226766 119016 226794
rect 119172 226794 119200 248386
rect 120000 227633 120028 263842
rect 121288 247625 121316 396743
rect 121274 247616 121330 247625
rect 121274 247551 121330 247560
rect 121380 229094 121408 398210
rect 121472 248414 121500 399774
rect 165620 398132 165672 398138
rect 165620 398074 165672 398080
rect 140780 397520 140832 397526
rect 140780 397462 140832 397468
rect 136454 397352 136510 397361
rect 136454 397287 136510 397296
rect 124126 396808 124182 396817
rect 124126 396743 124182 396752
rect 126886 396808 126942 396817
rect 126886 396743 126942 396752
rect 129646 396808 129702 396817
rect 129646 396743 129702 396752
rect 131026 396808 131082 396817
rect 131026 396743 131082 396752
rect 133786 396808 133842 396817
rect 133786 396743 133842 396752
rect 121472 248386 122144 248414
rect 121550 230072 121606 230081
rect 121550 230007 121606 230016
rect 121104 229066 121408 229094
rect 119986 227624 120042 227633
rect 119986 227559 120042 227568
rect 121104 226794 121132 229066
rect 119172 226766 119646 226794
rect 120658 226766 121132 226794
rect 121564 226780 121592 230007
rect 122116 226794 122144 248386
rect 124140 238105 124168 396743
rect 124220 264716 124272 264722
rect 124220 264658 124272 264664
rect 124126 238096 124182 238105
rect 124126 238031 124182 238040
rect 124232 233753 124260 264658
rect 125600 264104 125652 264110
rect 125600 264046 125652 264052
rect 124312 260908 124364 260914
rect 124312 260850 124364 260856
rect 124218 233744 124274 233753
rect 124218 233679 124274 233688
rect 123390 229936 123446 229945
rect 123390 229871 123446 229880
rect 122116 226766 122498 226794
rect 123404 226780 123432 229871
rect 124324 226780 124352 260850
rect 125612 248414 125640 264046
rect 125612 248386 125824 248414
rect 124862 233744 124918 233753
rect 124862 233679 124918 233688
rect 124876 226794 124904 233679
rect 125796 226794 125824 248386
rect 126900 235385 126928 396743
rect 128360 264172 128412 264178
rect 128360 264114 128412 264120
rect 126980 262608 127032 262614
rect 126980 262550 127032 262556
rect 126886 235376 126942 235385
rect 126886 235311 126942 235320
rect 126992 233753 127020 262550
rect 127072 262200 127124 262206
rect 127072 262142 127124 262148
rect 126978 233744 127034 233753
rect 126978 233679 127034 233688
rect 124876 226766 125258 226794
rect 125796 226766 126178 226794
rect 127084 226780 127112 262142
rect 128372 248414 128400 264114
rect 129660 249121 129688 396743
rect 131040 264722 131068 396743
rect 133800 264926 133828 396743
rect 136468 395622 136496 397287
rect 139306 396808 139362 396817
rect 139306 396743 139362 396752
rect 136456 395616 136508 395622
rect 136456 395558 136508 395564
rect 136640 373448 136692 373454
rect 136640 373390 136692 373396
rect 133880 373380 133932 373386
rect 133880 373322 133932 373328
rect 131120 264920 131172 264926
rect 131120 264862 131172 264868
rect 133788 264920 133840 264926
rect 133788 264862 133840 264868
rect 131028 264716 131080 264722
rect 131028 264658 131080 264664
rect 129740 262744 129792 262750
rect 129740 262686 129792 262692
rect 129646 249112 129702 249121
rect 129646 249047 129702 249056
rect 128372 248386 128584 248414
rect 127622 233744 127678 233753
rect 127622 233679 127678 233688
rect 127636 226794 127664 233679
rect 128556 226794 128584 248386
rect 129752 233753 129780 262686
rect 129832 261248 129884 261254
rect 129832 261190 129884 261196
rect 129738 233744 129794 233753
rect 129738 233679 129794 233688
rect 127636 226766 128018 226794
rect 128556 226766 128938 226794
rect 129844 226780 129872 261190
rect 131132 248414 131160 264862
rect 132500 262676 132552 262682
rect 132500 262618 132552 262624
rect 131132 248386 131344 248414
rect 130382 233744 130438 233753
rect 130382 233679 130438 233688
rect 130396 226794 130424 233679
rect 131316 226794 131344 248386
rect 132512 233753 132540 262618
rect 132592 261316 132644 261322
rect 132592 261258 132644 261264
rect 132498 233744 132554 233753
rect 132498 233679 132554 233688
rect 130396 226766 130778 226794
rect 131316 226766 131698 226794
rect 132604 226780 132632 261258
rect 133892 248414 133920 373322
rect 135260 261180 135312 261186
rect 135260 261122 135312 261128
rect 133892 248386 134104 248414
rect 133142 233744 133198 233753
rect 133142 233679 133198 233688
rect 133156 226794 133184 233679
rect 134076 226794 134104 248386
rect 135272 233753 135300 261122
rect 135352 260636 135404 260642
rect 135352 260578 135404 260584
rect 135258 233744 135314 233753
rect 135258 233679 135314 233688
rect 135364 226794 135392 260578
rect 136652 248414 136680 373390
rect 139320 264178 139348 396743
rect 139308 264172 139360 264178
rect 139308 264114 139360 264120
rect 139400 264036 139452 264042
rect 139400 263978 139452 263984
rect 138020 262540 138072 262546
rect 138020 262482 138072 262488
rect 136652 248386 136864 248414
rect 135902 233744 135958 233753
rect 135902 233679 135958 233688
rect 135916 226794 135944 233679
rect 136836 226794 136864 248386
rect 138032 233753 138060 262482
rect 138112 261384 138164 261390
rect 138112 261326 138164 261332
rect 138018 233744 138074 233753
rect 138018 233679 138074 233688
rect 138124 226794 138152 261326
rect 139412 248414 139440 263978
rect 139412 248386 139624 248414
rect 138662 233744 138718 233753
rect 138662 233679 138718 233688
rect 138676 226794 138704 233679
rect 139596 226794 139624 248386
rect 140792 233753 140820 397462
rect 154118 397352 154174 397361
rect 154118 397287 154174 397296
rect 163870 397352 163926 397361
rect 163870 397287 163926 397296
rect 142066 396808 142122 396817
rect 142066 396743 142122 396752
rect 144826 396808 144882 396817
rect 144826 396743 144882 396752
rect 145010 396808 145066 396817
rect 145010 396743 145066 396752
rect 148966 396808 149022 396817
rect 148966 396743 149022 396752
rect 151726 396808 151782 396817
rect 151726 396743 151782 396752
rect 140872 261452 140924 261458
rect 140872 261394 140924 261400
rect 140778 233744 140834 233753
rect 140778 233679 140834 233688
rect 140884 226794 140912 261394
rect 142080 261322 142108 396743
rect 142160 373312 142212 373318
rect 142160 373254 142212 373260
rect 142068 261316 142120 261322
rect 142068 261258 142120 261264
rect 142172 248414 142200 373254
rect 143540 371272 143592 371278
rect 143540 371214 143592 371220
rect 142172 248386 142384 248414
rect 141422 233744 141478 233753
rect 141422 233679 141478 233688
rect 141436 226794 141464 233679
rect 142356 226794 142384 248386
rect 143552 226794 143580 371214
rect 143632 345092 143684 345098
rect 143632 345034 143684 345040
rect 143644 248414 143672 345034
rect 144840 262206 144868 396743
rect 144920 357468 144972 357474
rect 144920 357410 144972 357416
rect 144828 262200 144880 262206
rect 144828 262142 144880 262148
rect 144932 248414 144960 357410
rect 145024 356726 145052 396743
rect 145012 356720 145064 356726
rect 145012 356662 145064 356668
rect 146300 318844 146352 318850
rect 146300 318786 146352 318792
rect 143644 248386 144224 248414
rect 144932 248386 145144 248414
rect 144196 226794 144224 248386
rect 145116 226794 145144 248386
rect 146312 226794 146340 318786
rect 147680 305040 147732 305046
rect 147680 304982 147732 304988
rect 146392 292596 146444 292602
rect 146392 292538 146444 292544
rect 146404 248414 146432 292538
rect 147692 248414 147720 304982
rect 148980 261254 149008 396743
rect 149060 266416 149112 266422
rect 149060 266358 149112 266364
rect 148968 261248 149020 261254
rect 148968 261190 149020 261196
rect 146404 248386 146984 248414
rect 147692 248386 147904 248414
rect 146956 226794 146984 248386
rect 147876 226794 147904 248386
rect 149072 226794 149100 266358
rect 151740 262682 151768 396743
rect 154132 395826 154160 397287
rect 162124 396908 162176 396914
rect 162124 396850 162176 396856
rect 155958 396808 156014 396817
rect 155958 396743 156014 396752
rect 158626 396808 158682 396817
rect 158626 396743 158682 396752
rect 161386 396808 161442 396817
rect 161386 396743 161442 396752
rect 154120 395820 154172 395826
rect 154120 395762 154172 395768
rect 155972 264858 156000 396743
rect 155960 264852 156012 264858
rect 155960 264794 156012 264800
rect 151728 262676 151780 262682
rect 151728 262618 151780 262624
rect 150806 236736 150862 236745
rect 150806 236671 150862 236680
rect 149702 233880 149758 233889
rect 149702 233815 149758 233824
rect 149716 226794 149744 233815
rect 150820 226794 150848 236671
rect 155406 233472 155462 233481
rect 155406 233407 155462 233416
rect 152094 231296 152150 231305
rect 152094 231231 152150 231240
rect 133156 226766 133538 226794
rect 134076 226766 134458 226794
rect 135364 226766 135470 226794
rect 135916 226766 136390 226794
rect 136836 226766 137310 226794
rect 138124 226766 138230 226794
rect 138676 226766 139150 226794
rect 139596 226766 140070 226794
rect 140884 226766 140990 226794
rect 141436 226766 141910 226794
rect 142356 226766 142830 226794
rect 143552 226766 143750 226794
rect 144196 226766 144670 226794
rect 145116 226766 145590 226794
rect 146312 226766 146510 226794
rect 146956 226766 147430 226794
rect 147876 226766 148350 226794
rect 149072 226766 149270 226794
rect 149716 226766 150190 226794
rect 150820 226766 151202 226794
rect 152108 226780 152136 231231
rect 154854 231160 154910 231169
rect 154854 231095 154910 231104
rect 153934 229800 153990 229809
rect 153934 229735 153990 229744
rect 153014 229120 153070 229129
rect 153014 229055 153070 229064
rect 153028 226780 153056 229055
rect 153948 226780 153976 229735
rect 154868 226780 154896 231095
rect 155420 226794 155448 233407
rect 158640 232529 158668 396743
rect 161400 264110 161428 396743
rect 161388 264104 161440 264110
rect 161388 264046 161440 264052
rect 162136 262750 162164 396850
rect 163884 396030 163912 397287
rect 163872 396024 163924 396030
rect 163872 395966 163924 395972
rect 162124 262744 162176 262750
rect 162124 262686 162176 262692
rect 161018 233336 161074 233345
rect 161018 233271 161074 233280
rect 158166 232520 158222 232529
rect 158166 232455 158222 232464
rect 158626 232520 158682 232529
rect 158626 232455 158682 232464
rect 157614 231024 157670 231033
rect 157614 230959 157670 230968
rect 156694 229664 156750 229673
rect 156694 229599 156750 229608
rect 155866 229256 155922 229265
rect 155866 229191 155922 229200
rect 155880 228313 155908 229191
rect 155866 228304 155922 228313
rect 155866 228239 155922 228248
rect 155420 226766 155802 226794
rect 156708 226780 156736 229599
rect 157628 226780 157656 230959
rect 158180 226794 158208 232455
rect 160190 232384 160246 232393
rect 160190 232319 160246 232328
rect 158718 232248 158774 232257
rect 158718 232183 158774 232192
rect 158732 229809 158760 232183
rect 158718 229800 158774 229809
rect 158718 229735 158774 229744
rect 159454 229120 159510 229129
rect 159454 229055 159510 229064
rect 158180 226766 158562 226794
rect 159468 226780 159496 229055
rect 160204 226794 160232 232319
rect 161032 226794 161060 233271
rect 162858 232112 162914 232121
rect 162858 232047 162914 232056
rect 162214 229528 162270 229537
rect 162214 229463 162270 229472
rect 160204 226766 160402 226794
rect 161032 226766 161322 226794
rect 162228 226780 162256 229463
rect 162872 226794 162900 232047
rect 164974 229800 165030 229809
rect 164974 229735 165030 229744
rect 164054 229256 164110 229265
rect 164054 229191 164110 229200
rect 162872 226766 163162 226794
rect 164068 226780 164096 229191
rect 164988 226780 165016 229735
rect 165632 226794 165660 398074
rect 173164 396908 173216 396914
rect 173164 396850 173216 396856
rect 168380 396840 168432 396846
rect 166906 396808 166962 396817
rect 168380 396782 168432 396788
rect 166906 396743 166962 396752
rect 165712 263832 165764 263838
rect 165712 263774 165764 263780
rect 165724 248414 165752 263774
rect 165724 248386 166488 248414
rect 166460 226794 166488 248386
rect 166920 233753 166948 396743
rect 168392 233889 168420 396782
rect 171048 395752 171100 395758
rect 171048 395694 171100 395700
rect 168472 267028 168524 267034
rect 168472 266970 168524 266976
rect 168378 233880 168434 233889
rect 168378 233815 168434 233824
rect 166906 233744 166962 233753
rect 166906 233679 166962 233688
rect 167826 229800 167882 229809
rect 167826 229735 167882 229744
rect 165632 226766 166014 226794
rect 166460 226766 166934 226794
rect 167840 226780 167868 229735
rect 168484 226794 168512 266970
rect 169298 233880 169354 233889
rect 169298 233815 169354 233824
rect 169312 226794 169340 233815
rect 171060 229094 171088 395694
rect 173176 260846 173204 396850
rect 177856 393984 177908 393990
rect 177856 393926 177908 393932
rect 175280 265940 175332 265946
rect 175280 265882 175332 265888
rect 173808 264852 173860 264858
rect 173808 264794 173860 264800
rect 172428 260840 172480 260846
rect 172428 260782 172480 260788
rect 173164 260840 173216 260846
rect 173164 260782 173216 260788
rect 171506 229936 171562 229945
rect 171506 229871 171562 229880
rect 170968 229066 171088 229094
rect 170968 226794 170996 229066
rect 168484 226766 168774 226794
rect 169312 226766 169694 226794
rect 170614 226766 170996 226794
rect 171520 226780 171548 229871
rect 172440 226780 172468 260782
rect 173820 229094 173848 264794
rect 173900 262744 173952 262750
rect 173900 262686 173952 262692
rect 173912 248414 173940 262686
rect 175292 248414 175320 265882
rect 173912 248386 174768 248414
rect 175292 248386 175688 248414
rect 174266 230072 174322 230081
rect 174266 230007 174322 230016
rect 173728 229066 173848 229094
rect 173728 226794 173756 229066
rect 173374 226766 173756 226794
rect 174280 226780 174308 230007
rect 174740 226794 174768 248386
rect 175660 226794 175688 248386
rect 177302 233744 177358 233753
rect 177302 233679 177358 233688
rect 177316 226794 177344 233679
rect 174740 226766 175214 226794
rect 175660 226766 176134 226794
rect 177054 226766 177344 226794
rect 177868 226794 177896 393926
rect 177960 233753 177988 399774
rect 183466 397352 183522 397361
rect 183466 397287 183522 397296
rect 183480 397118 183508 397287
rect 183468 397112 183520 397118
rect 183468 397054 183520 397060
rect 188344 396976 188396 396982
rect 188344 396918 188396 396924
rect 186964 396840 187016 396846
rect 182178 396808 182234 396817
rect 186964 396782 187016 396788
rect 182178 396743 182234 396752
rect 182088 265940 182140 265946
rect 182088 265882 182140 265888
rect 178040 265532 178092 265538
rect 178040 265474 178092 265480
rect 178052 248414 178080 265474
rect 181996 262744 182048 262750
rect 181996 262686 182048 262692
rect 178052 248386 178448 248414
rect 177946 233744 178002 233753
rect 177946 233679 178002 233688
rect 178420 226794 178448 248386
rect 181166 233744 181222 233753
rect 181166 233679 181222 233688
rect 179786 230344 179842 230353
rect 179786 230279 179842 230288
rect 177868 226766 177974 226794
rect 178420 226766 178894 226794
rect 179800 226780 179828 230279
rect 181180 226794 181208 233679
rect 182008 226794 182036 262686
rect 182100 233753 182128 265882
rect 182192 250481 182220 396743
rect 184940 395888 184992 395894
rect 184940 395830 184992 395836
rect 184848 395684 184900 395690
rect 184848 395626 184900 395632
rect 184756 264988 184808 264994
rect 184756 264930 184808 264936
rect 182178 250472 182234 250481
rect 182178 250407 182234 250416
rect 182086 233744 182142 233753
rect 182086 233679 182142 233688
rect 183926 233744 183982 233753
rect 183926 233679 183982 233688
rect 182638 230208 182694 230217
rect 182638 230143 182694 230152
rect 182178 229392 182234 229401
rect 182178 229327 182234 229336
rect 182192 228313 182220 229327
rect 182178 228304 182234 228313
rect 182178 228239 182234 228248
rect 180826 226766 181208 226794
rect 181746 226766 182036 226794
rect 182652 226780 182680 230143
rect 183940 226794 183968 233679
rect 184768 226794 184796 264930
rect 184860 233753 184888 395626
rect 184952 248414 184980 395830
rect 186976 264994 187004 396782
rect 187608 265532 187660 265538
rect 187608 265474 187660 265480
rect 186964 264988 187016 264994
rect 186964 264930 187016 264936
rect 184952 248386 185072 248414
rect 184846 233744 184902 233753
rect 184846 233679 184902 233688
rect 183586 226766 183968 226794
rect 184506 226766 184796 226794
rect 185044 226794 185072 248386
rect 186318 229664 186374 229673
rect 186318 229599 186374 229608
rect 185044 226766 185426 226794
rect 186332 226780 186360 229599
rect 187620 226794 187648 265474
rect 188356 262750 188384 396918
rect 189080 395956 189132 395962
rect 189080 395898 189132 395904
rect 188344 262744 188396 262750
rect 188344 262686 188396 262692
rect 188158 230480 188214 230489
rect 188158 230415 188214 230424
rect 187266 226766 187648 226794
rect 188172 226780 188200 230415
rect 189092 226780 189120 395898
rect 195888 395888 195940 395894
rect 195888 395830 195940 395836
rect 193128 392624 193180 392630
rect 193128 392566 193180 392572
rect 193036 261452 193088 261458
rect 193036 261394 193088 261400
rect 190368 261384 190420 261390
rect 190368 261326 190420 261332
rect 190380 226794 190408 261326
rect 192206 233744 192262 233753
rect 192206 233679 192262 233688
rect 190734 230344 190790 230353
rect 190918 230344 190974 230353
rect 190790 230302 190868 230330
rect 190734 230279 190790 230288
rect 190840 230081 190868 230302
rect 190918 230279 190974 230288
rect 190826 230072 190882 230081
rect 190826 230007 190882 230016
rect 190458 229936 190514 229945
rect 190514 229894 190684 229922
rect 190458 229871 190514 229880
rect 190656 229809 190684 229894
rect 190458 229800 190514 229809
rect 190458 229735 190514 229744
rect 190642 229800 190698 229809
rect 190642 229735 190698 229744
rect 190472 229537 190500 229735
rect 190458 229528 190514 229537
rect 190458 229463 190514 229472
rect 190026 226766 190408 226794
rect 190932 226780 190960 230279
rect 192220 226794 192248 233679
rect 193048 226794 193076 261394
rect 193140 233753 193168 392566
rect 195796 373312 195848 373318
rect 195796 373254 195848 373260
rect 193220 266280 193272 266286
rect 193220 266222 193272 266228
rect 193232 248414 193260 266222
rect 193232 248386 193352 248414
rect 193126 233744 193182 233753
rect 193126 233679 193182 233688
rect 191866 226766 192248 226794
rect 192786 226766 193076 226794
rect 193324 226794 193352 248386
rect 195808 229094 195836 373254
rect 195072 229066 195836 229094
rect 195072 226794 195100 229066
rect 195900 226794 195928 395830
rect 195980 266348 196032 266354
rect 195980 266290 196032 266296
rect 195992 248414 196020 266290
rect 196544 263906 196572 700334
rect 196624 700324 196676 700330
rect 196624 700266 196676 700272
rect 198004 700324 198056 700330
rect 198004 700266 198056 700272
rect 196636 398274 196664 700266
rect 197450 485480 197506 485489
rect 197450 485415 197506 485424
rect 196806 485072 196862 485081
rect 196806 485007 196862 485016
rect 196714 484936 196770 484945
rect 196714 484871 196770 484880
rect 196624 398268 196676 398274
rect 196624 398210 196676 398216
rect 196532 263900 196584 263906
rect 196532 263842 196584 263848
rect 195992 248386 196112 248414
rect 193324 226766 193706 226794
rect 194626 226766 195100 226794
rect 195638 226766 195928 226794
rect 196084 226794 196112 248386
rect 196728 229673 196756 484871
rect 196820 230353 196848 485007
rect 197358 484800 197414 484809
rect 197358 484735 197414 484744
rect 196806 230344 196862 230353
rect 196806 230279 196862 230288
rect 197372 230081 197400 484735
rect 197358 230072 197414 230081
rect 197358 230007 197414 230016
rect 197464 229945 197492 485415
rect 197634 484120 197690 484129
rect 197634 484055 197690 484064
rect 197542 483984 197598 483993
rect 197542 483919 197598 483928
rect 197450 229936 197506 229945
rect 197450 229871 197506 229880
rect 197556 229809 197584 483919
rect 197542 229800 197598 229809
rect 197542 229735 197598 229744
rect 196714 229664 196770 229673
rect 196714 229599 196770 229608
rect 197648 229537 197676 484055
rect 197726 417752 197782 417761
rect 197726 417687 197782 417696
rect 197740 239465 197768 417687
rect 198016 260982 198044 700266
rect 201038 486296 201094 486305
rect 201038 486231 201094 486240
rect 200854 485888 200910 485897
rect 200854 485823 200910 485832
rect 200762 485072 200818 485081
rect 200762 485007 200818 485016
rect 198646 484936 198702 484945
rect 198646 484871 198702 484880
rect 198096 264920 198148 264926
rect 198096 264862 198148 264868
rect 198004 260976 198056 260982
rect 198004 260918 198056 260924
rect 197726 239456 197782 239465
rect 197726 239391 197782 239400
rect 198108 230353 198136 264862
rect 198556 262744 198608 262750
rect 198556 262686 198608 262692
rect 198094 230344 198150 230353
rect 198094 230279 198150 230288
rect 197634 229528 197690 229537
rect 197634 229463 197690 229472
rect 198568 229094 198596 262686
rect 197832 229066 198596 229094
rect 197832 226794 197860 229066
rect 198660 226794 198688 484871
rect 199382 479224 199438 479233
rect 199382 479159 199438 479168
rect 198738 416392 198794 416401
rect 198738 416327 198794 416336
rect 198752 243681 198780 416327
rect 198738 243672 198794 243681
rect 198738 243607 198794 243616
rect 199396 234161 199424 479159
rect 199658 419384 199714 419393
rect 199658 419319 199714 419328
rect 199474 414896 199530 414905
rect 199474 414831 199530 414840
rect 199382 234152 199438 234161
rect 199382 234087 199438 234096
rect 199290 230344 199346 230353
rect 199290 230279 199346 230288
rect 196084 226766 196558 226794
rect 197478 226766 197860 226794
rect 198398 226766 198688 226794
rect 199304 226780 199332 230279
rect 199488 228585 199516 414831
rect 199566 413672 199622 413681
rect 199566 413607 199622 413616
rect 199580 232665 199608 413607
rect 199672 260846 199700 419319
rect 200120 265600 200172 265606
rect 200120 265542 200172 265548
rect 199660 260840 199712 260846
rect 199660 260782 199712 260788
rect 200132 248414 200160 265542
rect 200132 248386 200712 248414
rect 200486 233744 200542 233753
rect 200486 233679 200542 233688
rect 199566 232656 199622 232665
rect 199566 232591 199622 232600
rect 199474 228576 199530 228585
rect 199474 228511 199530 228520
rect 200500 226794 200528 233679
rect 200238 226766 200528 226794
rect 200684 226794 200712 248386
rect 200776 230489 200804 485007
rect 200868 261186 200896 485823
rect 201052 322153 201080 486231
rect 201038 322144 201094 322153
rect 201038 322079 201094 322088
rect 201408 264036 201460 264042
rect 201408 263978 201460 263984
rect 200856 261180 200908 261186
rect 200856 261122 200908 261128
rect 201420 233753 201448 263978
rect 201512 262478 201540 702986
rect 215944 700732 215996 700738
rect 215944 700674 215996 700680
rect 209044 700664 209096 700670
rect 209044 700606 209096 700612
rect 206376 700596 206428 700602
rect 206376 700538 206428 700544
rect 206284 700528 206336 700534
rect 206284 700470 206336 700476
rect 204904 700460 204956 700466
rect 204904 700402 204956 700408
rect 202142 487928 202198 487937
rect 202142 487863 202198 487872
rect 201592 264172 201644 264178
rect 201592 264114 201644 264120
rect 201500 262472 201552 262478
rect 201500 262414 201552 262420
rect 201406 233744 201462 233753
rect 201406 233679 201462 233688
rect 200762 230480 200818 230489
rect 200762 230415 200818 230424
rect 201604 226794 201632 264114
rect 202156 230217 202184 487863
rect 204258 487792 204314 487801
rect 204258 487727 204314 487736
rect 202880 266212 202932 266218
rect 202880 266154 202932 266160
rect 202142 230208 202198 230217
rect 202142 230143 202198 230152
rect 202892 226794 202920 266154
rect 202972 262200 203024 262206
rect 202972 262142 203024 262148
rect 202984 248414 203012 262142
rect 204272 248414 204300 487727
rect 204916 399770 204944 700402
rect 204904 399764 204956 399770
rect 204904 399706 204956 399712
rect 205640 263968 205692 263974
rect 205640 263910 205692 263916
rect 205652 248414 205680 263910
rect 206296 260778 206324 700470
rect 206388 398206 206416 700538
rect 206376 398200 206428 398206
rect 206376 398142 206428 398148
rect 206928 397044 206980 397050
rect 206928 396986 206980 396992
rect 206284 260772 206336 260778
rect 206284 260714 206336 260720
rect 202984 248386 203472 248414
rect 204272 248386 204392 248414
rect 205652 248386 206232 248414
rect 203444 226794 203472 248386
rect 204364 226794 204392 248386
rect 206006 230480 206062 230489
rect 206006 230415 206062 230424
rect 206020 226794 206048 230415
rect 200684 226766 201158 226794
rect 201604 226766 202078 226794
rect 202892 226766 202998 226794
rect 203444 226766 203918 226794
rect 204364 226766 204838 226794
rect 205758 226766 206048 226794
rect 206204 226794 206232 248386
rect 206940 230489 206968 396986
rect 209056 260710 209084 700606
rect 213184 700392 213236 700398
rect 213184 700334 213236 700340
rect 210424 699712 210476 699718
rect 210424 699654 210476 699660
rect 209134 486976 209190 486985
rect 209134 486911 209190 486920
rect 209044 260704 209096 260710
rect 209044 260646 209096 260652
rect 208308 260636 208360 260642
rect 208308 260578 208360 260584
rect 208320 234614 208348 260578
rect 209148 239465 209176 486911
rect 209318 486160 209374 486169
rect 209318 486095 209374 486104
rect 209228 430636 209280 430642
rect 209228 430578 209280 430584
rect 209240 399838 209268 430578
rect 209228 399832 209280 399838
rect 209228 399774 209280 399780
rect 209332 260137 209360 486095
rect 209686 484800 209742 484809
rect 209686 484735 209742 484744
rect 209596 264920 209648 264926
rect 209596 264862 209648 264868
rect 209318 260128 209374 260137
rect 209318 260063 209374 260072
rect 209134 239456 209190 239465
rect 209134 239391 209190 239400
rect 207952 234586 208348 234614
rect 206926 230480 206982 230489
rect 206926 230415 206982 230424
rect 207952 226794 207980 234586
rect 208766 230480 208822 230489
rect 208766 230415 208822 230424
rect 208780 226794 208808 230415
rect 209608 226794 209636 264862
rect 209700 230489 209728 484735
rect 210436 261050 210464 699654
rect 210514 486704 210570 486713
rect 210514 486639 210570 486648
rect 210424 261044 210476 261050
rect 210424 260986 210476 260992
rect 209686 230480 209742 230489
rect 209686 230415 209742 230424
rect 210528 229809 210556 486639
rect 211158 485208 211214 485217
rect 211158 485143 211214 485152
rect 211068 262200 211120 262206
rect 211068 262142 211120 262148
rect 211080 234614 211108 262142
rect 210896 234586 211108 234614
rect 210514 229800 210570 229809
rect 210514 229735 210570 229744
rect 210896 226794 210924 234586
rect 211172 230489 211200 485143
rect 213196 305658 213224 700334
rect 213368 510672 213420 510678
rect 213368 510614 213420 510620
rect 213274 486840 213330 486849
rect 213274 486775 213330 486784
rect 213184 305652 213236 305658
rect 213184 305594 213236 305600
rect 212540 262676 212592 262682
rect 212540 262618 212592 262624
rect 211252 261248 211304 261254
rect 211252 261190 211304 261196
rect 211158 230480 211214 230489
rect 211158 230415 211214 230424
rect 206204 226766 206678 226794
rect 207598 226766 207980 226794
rect 208518 226766 208808 226794
rect 209438 226766 209636 226794
rect 210450 226766 210924 226794
rect 211264 226794 211292 261190
rect 212552 248414 212580 262618
rect 212552 248386 212856 248414
rect 211986 230480 212042 230489
rect 211986 230415 212042 230424
rect 212000 226794 212028 230415
rect 212828 226794 212856 248386
rect 213288 234297 213316 486775
rect 213380 260574 213408 510614
rect 214562 487248 214618 487257
rect 214562 487183 214618 487192
rect 213458 486568 213514 486577
rect 213458 486503 213514 486512
rect 213368 260568 213420 260574
rect 213368 260510 213420 260516
rect 213472 250481 213500 486503
rect 213642 486432 213698 486441
rect 213642 486367 213698 486376
rect 213656 260574 213684 486367
rect 213918 485344 213974 485353
rect 213918 485279 213974 485288
rect 213644 260568 213696 260574
rect 213644 260510 213696 260516
rect 213458 250472 213514 250481
rect 213458 250407 213514 250416
rect 213932 248414 213960 485279
rect 214576 484537 214604 487183
rect 214562 484528 214618 484537
rect 214562 484463 214618 484472
rect 215206 484528 215262 484537
rect 215206 484463 215262 484472
rect 214576 408406 214604 484463
rect 214564 408400 214616 408406
rect 214564 408342 214616 408348
rect 214576 398818 214604 408342
rect 214564 398812 214616 398818
rect 214564 398754 214616 398760
rect 213932 248386 214696 248414
rect 213274 234288 213330 234297
rect 213274 234223 213330 234232
rect 214470 230480 214526 230489
rect 214470 230415 214526 230424
rect 214484 226794 214512 230415
rect 211264 226766 211370 226794
rect 212000 226766 212290 226794
rect 212828 226766 213210 226794
rect 214130 226766 214512 226794
rect 214668 226794 214696 248386
rect 215220 230489 215248 484463
rect 215956 261118 215984 700674
rect 218992 699718 219020 703520
rect 235184 700738 235212 703520
rect 235172 700732 235224 700738
rect 235172 700674 235224 700680
rect 267660 700670 267688 703520
rect 267648 700664 267700 700670
rect 267648 700606 267700 700612
rect 283852 700602 283880 703520
rect 283840 700596 283892 700602
rect 283840 700538 283892 700544
rect 300136 700534 300164 703520
rect 300124 700528 300176 700534
rect 300124 700470 300176 700476
rect 332520 700466 332548 703520
rect 332508 700460 332560 700466
rect 332508 700402 332560 700408
rect 348804 700398 348832 703520
rect 348792 700392 348844 700398
rect 348792 700334 348844 700340
rect 364996 700330 365024 703520
rect 397472 700602 397500 703520
rect 385684 700596 385736 700602
rect 385684 700538 385736 700544
rect 397460 700596 397512 700602
rect 397460 700538 397512 700544
rect 399484 700596 399536 700602
rect 399484 700538 399536 700544
rect 382924 700528 382976 700534
rect 382924 700470 382976 700476
rect 370504 700460 370556 700466
rect 370504 700402 370556 700408
rect 364984 700324 365036 700330
rect 364984 700266 365036 700272
rect 367744 700324 367796 700330
rect 367744 700266 367796 700272
rect 218980 699712 219032 699718
rect 218980 699654 219032 699660
rect 363604 670744 363656 670750
rect 363604 670686 363656 670692
rect 360844 616888 360896 616894
rect 360844 616830 360896 616836
rect 358084 563100 358136 563106
rect 358084 563042 358136 563048
rect 218702 490104 218758 490113
rect 218702 490039 218758 490048
rect 217966 487656 218022 487665
rect 217966 487591 218022 487600
rect 216310 487112 216366 487121
rect 216310 487047 216366 487056
rect 216034 486024 216090 486033
rect 216034 485959 216090 485968
rect 215944 261112 215996 261118
rect 215944 261054 215996 261060
rect 215206 230480 215262 230489
rect 215206 230415 215262 230424
rect 216048 229945 216076 485959
rect 216218 483712 216274 483721
rect 216218 483647 216274 483656
rect 216232 230353 216260 483647
rect 216324 232801 216352 487047
rect 217506 436928 217562 436937
rect 217506 436863 217562 436872
rect 216678 431080 216734 431089
rect 216678 431015 216734 431024
rect 216692 430642 216720 431015
rect 216680 430636 216732 430642
rect 216680 430578 216732 430584
rect 217414 429992 217470 430001
rect 217414 429927 217470 429936
rect 217230 410000 217286 410009
rect 217230 409935 217286 409944
rect 216680 408400 216732 408406
rect 216678 408368 216680 408377
rect 216732 408368 216734 408377
rect 216678 408303 216734 408312
rect 217138 408096 217194 408105
rect 217138 408031 217194 408040
rect 216588 397384 216640 397390
rect 216588 397326 216640 397332
rect 216404 264104 216456 264110
rect 216404 264046 216456 264052
rect 216310 232792 216366 232801
rect 216310 232727 216366 232736
rect 216416 230489 216444 264046
rect 216600 234614 216628 397326
rect 216508 234586 216628 234614
rect 216402 230480 216458 230489
rect 216402 230415 216458 230424
rect 216218 230344 216274 230353
rect 216218 230279 216274 230288
rect 216034 229936 216090 229945
rect 216034 229871 216090 229880
rect 216508 226794 216536 234586
rect 217152 228721 217180 408031
rect 217244 242321 217272 409935
rect 217428 399770 217456 429927
rect 217416 399764 217468 399770
rect 217416 399706 217468 399712
rect 217520 398138 217548 436863
rect 217690 435976 217746 435985
rect 217690 435911 217746 435920
rect 217598 428224 217654 428233
rect 217598 428159 217654 428168
rect 217612 399906 217640 428159
rect 217600 399900 217652 399906
rect 217600 399842 217652 399848
rect 217704 399838 217732 435911
rect 217782 433800 217838 433809
rect 217782 433735 217838 433744
rect 217692 399832 217744 399838
rect 217692 399774 217744 399780
rect 217508 398132 217560 398138
rect 217508 398074 217560 398080
rect 217230 242312 217286 242321
rect 217230 242247 217286 242256
rect 217796 238241 217824 433735
rect 217874 432848 217930 432857
rect 217874 432783 217930 432792
rect 217782 238232 217838 238241
rect 217782 238167 217838 238176
rect 217888 231169 217916 432783
rect 217874 231160 217930 231169
rect 217874 231095 217930 231104
rect 217980 230602 218008 487591
rect 218150 486704 218206 486713
rect 218150 486639 218206 486648
rect 218058 483848 218114 483857
rect 218058 483783 218114 483792
rect 218072 398206 218100 483783
rect 218164 400042 218192 486639
rect 218426 486568 218482 486577
rect 218426 486503 218482 486512
rect 218242 486296 218298 486305
rect 218242 486231 218298 486240
rect 218152 400036 218204 400042
rect 218152 399978 218204 399984
rect 218256 399974 218284 486231
rect 218334 483576 218390 483585
rect 218334 483511 218390 483520
rect 218244 399968 218296 399974
rect 218244 399910 218296 399916
rect 218060 398200 218112 398206
rect 218060 398142 218112 398148
rect 218348 231577 218376 483511
rect 218440 399430 218468 486503
rect 218610 486024 218666 486033
rect 218610 485959 218666 485968
rect 218518 484256 218574 484265
rect 218518 484191 218574 484200
rect 218428 399424 218480 399430
rect 218428 399366 218480 399372
rect 218334 231568 218390 231577
rect 218334 231503 218390 231512
rect 218532 231033 218560 484191
rect 218624 400110 218652 485959
rect 218612 400104 218664 400110
rect 218612 400046 218664 400052
rect 218716 231305 218744 490039
rect 260838 489968 260894 489977
rect 260838 489903 260894 489912
rect 218978 489288 219034 489297
rect 218978 489223 219034 489232
rect 218886 488064 218942 488073
rect 218886 487999 218942 488008
rect 218794 486976 218850 486985
rect 218794 486911 218850 486920
rect 218808 398177 218836 486911
rect 218794 398168 218850 398177
rect 218794 398103 218850 398112
rect 218900 231441 218928 487999
rect 218992 398041 219020 489223
rect 219898 489152 219954 489161
rect 219898 489087 219954 489096
rect 219806 487792 219862 487801
rect 219806 487727 219862 487736
rect 219346 486432 219402 486441
rect 219346 486367 219402 486376
rect 219254 485888 219310 485897
rect 219254 485823 219310 485832
rect 219162 485344 219218 485353
rect 219162 485279 219218 485288
rect 219070 483576 219126 483585
rect 219070 483511 219126 483520
rect 218978 398032 219034 398041
rect 218978 397967 219034 397976
rect 218886 231432 218942 231441
rect 218886 231367 218942 231376
rect 218702 231296 218758 231305
rect 218702 231231 218758 231240
rect 218518 231024 218574 231033
rect 218518 230959 218574 230968
rect 217336 230574 218008 230602
rect 217138 228712 217194 228721
rect 217138 228647 217194 228656
rect 217336 226794 217364 230574
rect 219084 230489 219112 483511
rect 217782 230480 217838 230489
rect 217782 230415 217838 230424
rect 219070 230480 219126 230489
rect 219070 230415 219126 230424
rect 214668 226766 215050 226794
rect 215970 226766 216536 226794
rect 216890 226766 217364 226794
rect 217796 226780 217824 230415
rect 219176 226794 219204 485279
rect 219268 227225 219296 485823
rect 219254 227216 219310 227225
rect 219254 227151 219310 227160
rect 218730 226766 219204 226794
rect 62946 226672 63002 226681
rect 71686 226672 71742 226681
rect 71530 226630 71686 226658
rect 62946 226607 63002 226616
rect 71686 226607 71742 226616
rect 62762 226400 62818 226409
rect 68190 226400 68246 226409
rect 67850 226358 68190 226386
rect 62762 226335 62818 226344
rect 68190 226335 68246 226344
rect 219360 226273 219388 486367
rect 219714 485208 219770 485217
rect 219714 485143 219770 485152
rect 219530 483984 219586 483993
rect 219530 483919 219586 483928
rect 219544 398750 219572 483919
rect 219622 483712 219678 483721
rect 219622 483647 219678 483656
rect 219532 398744 219584 398750
rect 219532 398686 219584 398692
rect 219636 398614 219664 483647
rect 219624 398608 219676 398614
rect 219624 398550 219676 398556
rect 219728 398206 219756 485143
rect 219716 398200 219768 398206
rect 219820 398177 219848 487727
rect 219912 398546 219940 489087
rect 253386 489016 253442 489025
rect 253386 488951 253442 488960
rect 219990 486160 220046 486169
rect 219990 486095 220046 486104
rect 219900 398540 219952 398546
rect 219900 398482 219952 398488
rect 219716 398142 219768 398148
rect 219806 398168 219862 398177
rect 219806 398103 219862 398112
rect 219440 396024 219492 396030
rect 219440 395966 219492 395972
rect 219452 226794 219480 395966
rect 220004 227361 220032 486095
rect 253400 485897 253428 488951
rect 258354 488880 258410 488889
rect 258354 488815 258410 488824
rect 258368 485897 258396 488815
rect 260852 486577 260880 489903
rect 288530 489288 288586 489297
rect 288530 489223 288586 489232
rect 278410 488744 278466 488753
rect 278410 488679 278466 488688
rect 266082 487928 266138 487937
rect 266082 487863 266138 487872
rect 260838 486568 260894 486577
rect 260838 486503 260894 486512
rect 266096 485897 266124 487863
rect 273258 486432 273314 486441
rect 273258 486367 273314 486376
rect 253386 485888 253442 485897
rect 253386 485823 253442 485832
rect 258354 485888 258410 485897
rect 258354 485823 258410 485832
rect 266082 485888 266138 485897
rect 266082 485823 266138 485832
rect 273272 485353 273300 486367
rect 278424 485897 278452 488679
rect 288544 486305 288572 489223
rect 295890 489152 295946 489161
rect 295890 489087 295946 489096
rect 288530 486296 288586 486305
rect 288530 486231 288586 486240
rect 295904 486169 295932 489087
rect 310978 488608 311034 488617
rect 310978 488543 311034 488552
rect 301502 487384 301558 487393
rect 301502 487319 301558 487328
rect 301516 486577 301544 487319
rect 301502 486568 301558 486577
rect 301502 486503 301558 486512
rect 295890 486160 295946 486169
rect 295890 486095 295946 486104
rect 310992 485897 311020 488543
rect 313554 487792 313610 487801
rect 313554 487727 313610 487736
rect 313568 485897 313596 487727
rect 320270 487656 320326 487665
rect 320270 487591 320326 487600
rect 320284 485897 320312 487591
rect 340142 487248 340198 487257
rect 340142 487183 340198 487192
rect 340156 486441 340184 487183
rect 340142 486432 340198 486441
rect 340142 486367 340198 486376
rect 278410 485888 278466 485897
rect 278410 485823 278466 485832
rect 310978 485888 311034 485897
rect 310978 485823 311034 485832
rect 313554 485888 313610 485897
rect 313554 485823 313610 485832
rect 320270 485888 320326 485897
rect 320270 485823 320326 485832
rect 273258 485344 273314 485353
rect 273258 485279 273314 485288
rect 356518 484528 356574 484537
rect 356518 484463 356574 484472
rect 226340 400036 226392 400042
rect 226340 399978 226392 399984
rect 226708 400036 226760 400042
rect 226708 399978 226760 399984
rect 224960 398744 225012 398750
rect 224960 398686 225012 398692
rect 222844 396228 222896 396234
rect 222844 396170 222896 396176
rect 222856 251161 222884 396170
rect 224868 395548 224920 395554
rect 224868 395490 224920 395496
rect 223672 264784 223724 264790
rect 223672 264726 223724 264732
rect 223488 264172 223540 264178
rect 223488 264114 223540 264120
rect 222106 251152 222162 251161
rect 222106 251087 222162 251096
rect 222842 251152 222898 251161
rect 222842 251087 222898 251096
rect 222120 234614 222148 251087
rect 223500 238754 223528 264114
rect 221936 234586 222148 234614
rect 222856 238726 223528 238754
rect 220542 230344 220598 230353
rect 220542 230279 220598 230288
rect 219990 227352 220046 227361
rect 219990 227287 220046 227296
rect 219452 226766 219650 226794
rect 220556 226780 220584 230279
rect 221936 226794 221964 234586
rect 222856 226794 222884 238726
rect 223302 230480 223358 230489
rect 223302 230415 223358 230424
rect 221490 226766 221964 226794
rect 222410 226766 222884 226794
rect 223316 226780 223344 230415
rect 223684 228857 223712 264726
rect 224776 261180 224828 261186
rect 224776 261122 224828 261128
rect 224222 233880 224278 233889
rect 224222 233815 224278 233824
rect 223670 228848 223726 228857
rect 223670 228783 223726 228792
rect 224236 226780 224264 233815
rect 61106 226264 61162 226273
rect 61106 226199 61162 226208
rect 62026 226264 62082 226273
rect 62026 226199 62082 226208
rect 219346 226264 219402 226273
rect 219346 226199 219402 226208
rect 59832 113146 60044 113174
rect 59832 106282 59860 113146
rect 59820 106276 59872 106282
rect 59820 106218 59872 106224
rect 59372 74506 59768 74534
rect 58898 67824 58954 67833
rect 58898 67759 58954 67768
rect 59740 60058 59768 74506
rect 59740 60030 60122 60058
rect 59740 59922 59768 60030
rect 59372 59894 59768 59922
rect 58714 57896 58770 57905
rect 58714 57831 58770 57840
rect 58622 57760 58678 57769
rect 58622 57695 58678 57704
rect 58636 57361 58664 57695
rect 58622 57352 58678 57361
rect 58622 57287 58678 57296
rect 58530 57080 58586 57089
rect 58530 57015 58586 57024
rect 58254 56944 58310 56953
rect 58254 56879 58310 56888
rect 58268 56681 58296 56879
rect 59268 56704 59320 56710
rect 58254 56672 58310 56681
rect 57244 56636 57296 56642
rect 59268 56646 59320 56652
rect 58254 56607 58310 56616
rect 57244 56578 57296 56584
rect 55772 46232 55824 46238
rect 55772 46174 55824 46180
rect 57256 4146 57284 56578
rect 59280 4146 59308 56646
rect 56048 4140 56100 4146
rect 56048 4082 56100 4088
rect 57244 4140 57296 4146
rect 57244 4082 57296 4088
rect 58440 4140 58492 4146
rect 58440 4082 58492 4088
rect 59268 4140 59320 4146
rect 59268 4082 59320 4088
rect 55496 3732 55548 3738
rect 55496 3674 55548 3680
rect 55508 3534 55536 3674
rect 55220 3528 55272 3534
rect 55220 3470 55272 3476
rect 55496 3528 55548 3534
rect 55496 3470 55548 3476
rect 55232 2854 55260 3470
rect 55956 3256 56008 3262
rect 55784 3204 55956 3210
rect 55784 3198 56008 3204
rect 55784 3194 55996 3198
rect 55772 3188 55996 3194
rect 55824 3182 55996 3188
rect 55772 3130 55824 3136
rect 55956 3120 56008 3126
rect 55876 3068 55956 3074
rect 55876 3062 56008 3068
rect 55876 3046 55996 3062
rect 55876 2990 55904 3046
rect 55864 2984 55916 2990
rect 55864 2926 55916 2932
rect 55220 2848 55272 2854
rect 55220 2790 55272 2796
rect 54956 2746 55168 2774
rect 54956 480 54984 2746
rect 56060 480 56088 4082
rect 56140 3868 56192 3874
rect 56140 3810 56192 3816
rect 56152 3670 56180 3810
rect 56140 3664 56192 3670
rect 56140 3606 56192 3612
rect 56140 3120 56192 3126
rect 56140 3062 56192 3068
rect 56152 746 56180 3062
rect 57244 3052 57296 3058
rect 57244 2994 57296 3000
rect 56140 740 56192 746
rect 56140 682 56192 688
rect 57256 480 57284 2994
rect 58452 480 58480 4082
rect 59372 3466 59400 59894
rect 60384 57610 60412 60044
rect 59464 57582 60412 57610
rect 59360 3460 59412 3466
rect 59360 3402 59412 3408
rect 59464 2854 59492 57582
rect 60002 57488 60058 57497
rect 60002 57423 60058 57432
rect 59636 4140 59688 4146
rect 59636 4082 59688 4088
rect 59452 2848 59504 2854
rect 59452 2790 59504 2796
rect 59648 480 59676 4082
rect 60016 3534 60044 57423
rect 60660 57254 60688 60044
rect 60648 57248 60700 57254
rect 60832 57248 60884 57254
rect 60648 57190 60700 57196
rect 60752 57196 60832 57202
rect 60936 57225 60964 60044
rect 60752 57190 60884 57196
rect 60922 57216 60978 57225
rect 60752 57174 60872 57190
rect 60752 57066 60780 57174
rect 60922 57151 60978 57160
rect 60660 57038 60780 57066
rect 60660 4146 60688 57038
rect 60648 4140 60700 4146
rect 60648 4082 60700 4088
rect 61304 3670 61332 60044
rect 61580 57390 61608 60044
rect 61568 57384 61620 57390
rect 61568 57326 61620 57332
rect 61856 3874 61884 60044
rect 62132 57769 62160 60044
rect 62118 57760 62174 57769
rect 62118 57695 62174 57704
rect 62500 57361 62528 60044
rect 62776 57633 62804 60044
rect 62762 57624 62818 57633
rect 62762 57559 62818 57568
rect 63052 57497 63080 60044
rect 63038 57488 63094 57497
rect 63038 57423 63094 57432
rect 62486 57352 62542 57361
rect 62028 57316 62080 57322
rect 62486 57287 62542 57296
rect 62028 57258 62080 57264
rect 61844 3868 61896 3874
rect 61844 3810 61896 3816
rect 61292 3664 61344 3670
rect 61292 3606 61344 3612
rect 60004 3528 60056 3534
rect 60004 3470 60056 3476
rect 60832 3460 60884 3466
rect 60832 3402 60884 3408
rect 60844 480 60872 3402
rect 62040 480 62068 57258
rect 63328 56681 63356 60044
rect 63696 56953 63724 60044
rect 63682 56944 63738 56953
rect 63682 56879 63738 56888
rect 63314 56672 63370 56681
rect 63314 56607 63370 56616
rect 63972 3738 64000 60044
rect 64248 57390 64276 60044
rect 64236 57384 64288 57390
rect 64236 57326 64288 57332
rect 63960 3732 64012 3738
rect 63960 3674 64012 3680
rect 64328 3596 64380 3602
rect 64328 3538 64380 3544
rect 63224 3528 63276 3534
rect 63224 3470 63276 3476
rect 63236 480 63264 3470
rect 64340 480 64368 3538
rect 64524 2990 64552 60044
rect 64788 57384 64840 57390
rect 64788 57326 64840 57332
rect 64800 3602 64828 57326
rect 64892 55214 64920 60044
rect 64892 55186 65012 55214
rect 64984 3942 65012 55186
rect 65168 4010 65196 60044
rect 65444 56817 65472 60044
rect 65430 56808 65486 56817
rect 65430 56743 65486 56752
rect 65720 4078 65748 60044
rect 66088 57526 66116 60044
rect 66076 57520 66128 57526
rect 66076 57462 66128 57468
rect 66168 57520 66220 57526
rect 66168 57462 66220 57468
rect 65708 4072 65760 4078
rect 65708 4014 65760 4020
rect 65156 4004 65208 4010
rect 65156 3946 65208 3952
rect 64972 3936 65024 3942
rect 64972 3878 65024 3884
rect 64788 3596 64840 3602
rect 64788 3538 64840 3544
rect 66180 3534 66208 57462
rect 66364 57458 66392 60044
rect 66640 57594 66668 60044
rect 66916 57662 66944 60044
rect 66904 57656 66956 57662
rect 66904 57598 66956 57604
rect 66628 57588 66680 57594
rect 66628 57530 66680 57536
rect 66352 57452 66404 57458
rect 66352 57394 66404 57400
rect 67284 3806 67312 60044
rect 67560 57798 67588 60044
rect 67548 57792 67600 57798
rect 67548 57734 67600 57740
rect 67548 57656 67600 57662
rect 67548 57598 67600 57604
rect 67272 3800 67324 3806
rect 67272 3742 67324 3748
rect 67560 3534 67588 57598
rect 65524 3528 65576 3534
rect 65524 3470 65576 3476
rect 66168 3528 66220 3534
rect 66168 3470 66220 3476
rect 66720 3528 66772 3534
rect 66720 3470 66772 3476
rect 67548 3528 67600 3534
rect 67548 3470 67600 3476
rect 64512 2984 64564 2990
rect 64512 2926 64564 2932
rect 65536 480 65564 3470
rect 66732 480 66760 3470
rect 67836 3398 67864 60044
rect 68112 57730 68140 60044
rect 68480 57866 68508 60044
rect 68468 57860 68520 57866
rect 68468 57802 68520 57808
rect 68100 57724 68152 57730
rect 68100 57666 68152 57672
rect 68756 57186 68784 60044
rect 68744 57180 68796 57186
rect 68744 57122 68796 57128
rect 68928 57180 68980 57186
rect 68928 57122 68980 57128
rect 68940 3534 68968 57122
rect 69032 55214 69060 60044
rect 69032 55186 69244 55214
rect 67916 3528 67968 3534
rect 67916 3470 67968 3476
rect 68928 3528 68980 3534
rect 68928 3470 68980 3476
rect 69112 3528 69164 3534
rect 69112 3470 69164 3476
rect 67824 3392 67876 3398
rect 67824 3334 67876 3340
rect 67928 480 67956 3470
rect 69124 480 69152 3470
rect 69216 3330 69244 55186
rect 69308 54534 69336 60044
rect 69296 54528 69348 54534
rect 69296 54470 69348 54476
rect 69204 3324 69256 3330
rect 69204 3266 69256 3272
rect 69676 3262 69704 60044
rect 69952 57934 69980 60044
rect 69940 57928 69992 57934
rect 69940 57870 69992 57876
rect 70228 57610 70256 60044
rect 70136 57582 70256 57610
rect 70308 57588 70360 57594
rect 70136 57118 70164 57582
rect 70308 57530 70360 57536
rect 70216 57452 70268 57458
rect 70216 57394 70268 57400
rect 70124 57112 70176 57118
rect 70124 57054 70176 57060
rect 70228 3534 70256 57394
rect 70216 3528 70268 3534
rect 70216 3470 70268 3476
rect 69664 3256 69716 3262
rect 69664 3198 69716 3204
rect 70320 480 70348 57530
rect 70504 57050 70532 60044
rect 70492 57044 70544 57050
rect 70492 56986 70544 56992
rect 70872 54602 70900 60044
rect 71148 54670 71176 60044
rect 71424 54738 71452 60044
rect 71700 56982 71728 60044
rect 71688 56976 71740 56982
rect 71688 56918 71740 56924
rect 72068 56914 72096 60044
rect 72056 56908 72108 56914
rect 72056 56850 72108 56856
rect 72148 56908 72200 56914
rect 72148 56850 72200 56856
rect 72160 56642 72188 56850
rect 72148 56636 72200 56642
rect 72148 56578 72200 56584
rect 72344 54806 72372 60044
rect 72424 56636 72476 56642
rect 72424 56578 72476 56584
rect 72332 54800 72384 54806
rect 72332 54742 72384 54748
rect 71412 54732 71464 54738
rect 71412 54674 71464 54680
rect 71136 54664 71188 54670
rect 71136 54606 71188 54612
rect 70860 54596 70912 54602
rect 70860 54538 70912 54544
rect 71504 4072 71556 4078
rect 71504 4014 71556 4020
rect 71516 480 71544 4014
rect 72436 3602 72464 56578
rect 72620 6914 72648 60044
rect 72528 6886 72648 6914
rect 72424 3596 72476 3602
rect 72424 3538 72476 3544
rect 72528 3194 72556 6886
rect 72608 3528 72660 3534
rect 72608 3470 72660 3476
rect 72516 3188 72568 3194
rect 72516 3130 72568 3136
rect 72620 480 72648 3470
rect 72988 3126 73016 60044
rect 73068 57724 73120 57730
rect 73068 57666 73120 57672
rect 73080 3534 73108 57666
rect 73264 54874 73292 60044
rect 73540 56846 73568 60044
rect 73528 56840 73580 56846
rect 73528 56782 73580 56788
rect 73816 56778 73844 60044
rect 74184 56914 74212 60044
rect 74172 56908 74224 56914
rect 74172 56850 74224 56856
rect 73804 56772 73856 56778
rect 73804 56714 73856 56720
rect 73252 54868 73304 54874
rect 73252 54810 73304 54816
rect 73068 3528 73120 3534
rect 73068 3470 73120 3476
rect 73804 3460 73856 3466
rect 73804 3402 73856 3408
rect 72976 3120 73028 3126
rect 72976 3062 73028 3068
rect 73816 480 73844 3402
rect 74460 3058 74488 60044
rect 74736 57050 74764 60044
rect 75012 57254 75040 60044
rect 75092 57860 75144 57866
rect 75092 57802 75144 57808
rect 75104 57458 75132 57802
rect 75092 57452 75144 57458
rect 75092 57394 75144 57400
rect 75184 57452 75236 57458
rect 75184 57394 75236 57400
rect 75000 57248 75052 57254
rect 75000 57190 75052 57196
rect 74724 57044 74776 57050
rect 74724 56986 74776 56992
rect 75000 3596 75052 3602
rect 75000 3538 75052 3544
rect 74448 3052 74500 3058
rect 74448 2994 74500 3000
rect 75012 480 75040 3538
rect 75196 3466 75224 57394
rect 75380 3534 75408 60044
rect 75656 57322 75684 60044
rect 75828 57588 75880 57594
rect 75828 57530 75880 57536
rect 75644 57316 75696 57322
rect 75644 57258 75696 57264
rect 75840 3602 75868 57530
rect 75932 56642 75960 60044
rect 76208 57390 76236 60044
rect 76576 57526 76604 60044
rect 76852 57934 76880 60044
rect 76840 57928 76892 57934
rect 76840 57870 76892 57876
rect 76564 57520 76616 57526
rect 76564 57462 76616 57468
rect 76196 57384 76248 57390
rect 76196 57326 76248 57332
rect 77128 57254 77156 60044
rect 77404 57866 77432 60044
rect 77392 57860 77444 57866
rect 77392 57802 77444 57808
rect 77772 57730 77800 60044
rect 77760 57724 77812 57730
rect 77760 57666 77812 57672
rect 77116 57248 77168 57254
rect 77116 57190 77168 57196
rect 78048 57186 78076 60044
rect 78324 57798 78352 60044
rect 78312 57792 78364 57798
rect 78312 57734 78364 57740
rect 78600 57458 78628 60044
rect 78968 57594 78996 60044
rect 78956 57588 79008 57594
rect 78956 57530 79008 57536
rect 78588 57452 78640 57458
rect 78588 57394 78640 57400
rect 76564 57180 76616 57186
rect 76564 57122 76616 57128
rect 78036 57180 78088 57186
rect 78036 57122 78088 57128
rect 75920 56636 75972 56642
rect 75920 56578 75972 56584
rect 76576 4078 76604 57122
rect 79244 57050 79272 60044
rect 77208 57044 77260 57050
rect 77208 56986 77260 56992
rect 79232 57044 79284 57050
rect 79232 56986 79284 56992
rect 76564 4072 76616 4078
rect 76564 4014 76616 4020
rect 75828 3596 75880 3602
rect 75828 3538 75880 3544
rect 77220 3534 77248 56986
rect 75368 3528 75420 3534
rect 75368 3470 75420 3476
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 75184 3460 75236 3466
rect 75184 3402 75236 3408
rect 76208 480 76236 3470
rect 78588 3392 78640 3398
rect 78588 3334 78640 3340
rect 77392 3188 77444 3194
rect 77392 3130 77444 3136
rect 77404 480 77432 3130
rect 78600 480 78628 3334
rect 79520 3194 79548 60044
rect 79692 3528 79744 3534
rect 79692 3470 79744 3476
rect 79508 3188 79560 3194
rect 79508 3130 79560 3136
rect 79704 480 79732 3470
rect 79796 3398 79824 60044
rect 80164 55214 80192 60044
rect 80164 55186 80376 55214
rect 80348 3534 80376 55186
rect 80440 3534 80468 60044
rect 80716 57662 80744 60044
rect 80704 57656 80756 57662
rect 80704 57598 80756 57604
rect 80992 56846 81020 60044
rect 81256 57656 81308 57662
rect 81256 57598 81308 57604
rect 80980 56840 81032 56846
rect 80980 56782 81032 56788
rect 81268 3534 81296 57598
rect 81360 3602 81388 60044
rect 81636 57458 81664 60044
rect 81912 57594 81940 60044
rect 82188 57662 82216 60044
rect 82176 57656 82228 57662
rect 82176 57598 82228 57604
rect 81900 57588 81952 57594
rect 81900 57530 81952 57536
rect 81624 57452 81676 57458
rect 81624 57394 81676 57400
rect 82452 57452 82504 57458
rect 82452 57394 82504 57400
rect 82464 4146 82492 57394
rect 82452 4140 82504 4146
rect 82452 4082 82504 4088
rect 82556 3670 82584 60044
rect 82636 57656 82688 57662
rect 82636 57598 82688 57604
rect 82648 3806 82676 57598
rect 82728 57588 82780 57594
rect 82728 57530 82780 57536
rect 82636 3800 82688 3806
rect 82636 3742 82688 3748
rect 82544 3664 82596 3670
rect 82544 3606 82596 3612
rect 81348 3596 81400 3602
rect 81348 3538 81400 3544
rect 80336 3528 80388 3534
rect 80336 3470 80388 3476
rect 80428 3528 80480 3534
rect 80428 3470 80480 3476
rect 80888 3528 80940 3534
rect 80888 3470 80940 3476
rect 81256 3528 81308 3534
rect 81256 3470 81308 3476
rect 82084 3528 82136 3534
rect 82084 3470 82136 3476
rect 79784 3392 79836 3398
rect 79784 3334 79836 3340
rect 80900 480 80928 3470
rect 82096 480 82124 3470
rect 82740 2854 82768 57530
rect 82832 57526 82860 60044
rect 83108 57662 83136 60044
rect 83096 57656 83148 57662
rect 83096 57598 83148 57604
rect 82820 57520 82872 57526
rect 82820 57462 82872 57468
rect 83384 57390 83412 60044
rect 83372 57384 83424 57390
rect 83372 57326 83424 57332
rect 83096 56840 83148 56846
rect 83096 56782 83148 56788
rect 83108 16574 83136 56782
rect 83752 55214 83780 60044
rect 84028 57610 84056 60044
rect 84304 57798 84332 60044
rect 84292 57792 84344 57798
rect 84292 57734 84344 57740
rect 84672 57730 84700 60044
rect 84660 57724 84712 57730
rect 84660 57666 84712 57672
rect 83936 57582 84056 57610
rect 84108 57656 84160 57662
rect 84108 57598 84160 57604
rect 83752 55186 83872 55214
rect 83108 16546 83320 16574
rect 82728 2848 82780 2854
rect 82728 2790 82780 2796
rect 83292 480 83320 16546
rect 83844 6186 83872 55186
rect 83832 6180 83884 6186
rect 83832 6122 83884 6128
rect 83936 3466 83964 57582
rect 84016 57520 84068 57526
rect 84016 57462 84068 57468
rect 84028 3738 84056 57462
rect 84016 3732 84068 3738
rect 84016 3674 84068 3680
rect 84120 3602 84148 57598
rect 84948 57050 84976 60044
rect 85224 57662 85252 60044
rect 85212 57656 85264 57662
rect 85212 57598 85264 57604
rect 84936 57044 84988 57050
rect 84936 56986 84988 56992
rect 85500 7614 85528 60044
rect 85868 57594 85896 60044
rect 85856 57588 85908 57594
rect 85856 57530 85908 57536
rect 86144 57322 86172 60044
rect 86316 57724 86368 57730
rect 86316 57666 86368 57672
rect 86224 57656 86276 57662
rect 86224 57598 86276 57604
rect 86132 57316 86184 57322
rect 86132 57258 86184 57264
rect 85488 7608 85540 7614
rect 85488 7550 85540 7556
rect 85672 4140 85724 4146
rect 85672 4082 85724 4088
rect 84108 3596 84160 3602
rect 84108 3538 84160 3544
rect 84476 3528 84528 3534
rect 84476 3470 84528 3476
rect 83924 3460 83976 3466
rect 83924 3402 83976 3408
rect 84488 480 84516 3470
rect 85684 480 85712 4082
rect 86236 3398 86264 57598
rect 86328 7682 86356 57666
rect 86420 57662 86448 60044
rect 86408 57656 86460 57662
rect 86408 57598 86460 57604
rect 86316 7676 86368 7682
rect 86316 7618 86368 7624
rect 86224 3392 86276 3398
rect 86224 3334 86276 3340
rect 86696 3126 86724 60044
rect 86868 57656 86920 57662
rect 86868 57598 86920 57604
rect 86776 57588 86828 57594
rect 86776 57530 86828 57536
rect 86684 3120 86736 3126
rect 86684 3062 86736 3068
rect 86788 2922 86816 57530
rect 86880 2990 86908 57598
rect 87064 57254 87092 60044
rect 87340 57526 87368 60044
rect 87328 57520 87380 57526
rect 87328 57462 87380 57468
rect 87616 57458 87644 60044
rect 87892 57934 87920 60044
rect 87880 57928 87932 57934
rect 87880 57870 87932 57876
rect 88260 57644 88288 60044
rect 88076 57616 88288 57644
rect 87604 57452 87656 57458
rect 87604 57394 87656 57400
rect 87052 57248 87104 57254
rect 87052 57190 87104 57196
rect 87604 57044 87656 57050
rect 87604 56986 87656 56992
rect 86868 2984 86920 2990
rect 86868 2926 86920 2932
rect 86776 2916 86828 2922
rect 86776 2858 86828 2864
rect 87616 2854 87644 56986
rect 88076 4010 88104 57616
rect 88536 57526 88564 60044
rect 88812 57730 88840 60044
rect 88984 57792 89036 57798
rect 88984 57734 89036 57740
rect 88800 57724 88852 57730
rect 88800 57666 88852 57672
rect 88156 57520 88208 57526
rect 88156 57462 88208 57468
rect 88524 57520 88576 57526
rect 88524 57462 88576 57468
rect 88064 4004 88116 4010
rect 88064 3946 88116 3952
rect 87972 3800 88024 3806
rect 87972 3742 88024 3748
rect 86868 2848 86920 2854
rect 86868 2790 86920 2796
rect 87604 2848 87656 2854
rect 87604 2790 87656 2796
rect 86880 480 86908 2790
rect 87984 480 88012 3742
rect 88168 3058 88196 57462
rect 88248 57452 88300 57458
rect 88248 57394 88300 57400
rect 88260 3194 88288 57394
rect 88996 3330 89024 57734
rect 89088 55214 89116 60044
rect 89456 57644 89484 60044
rect 89456 57616 89668 57644
rect 89536 57520 89588 57526
rect 89536 57462 89588 57468
rect 89088 55186 89484 55214
rect 89168 3664 89220 3670
rect 89168 3606 89220 3612
rect 88984 3324 89036 3330
rect 88984 3266 89036 3272
rect 88248 3188 88300 3194
rect 88248 3130 88300 3136
rect 88156 3052 88208 3058
rect 88156 2994 88208 3000
rect 89180 480 89208 3606
rect 89456 3398 89484 55186
rect 89444 3392 89496 3398
rect 89444 3334 89496 3340
rect 89548 3262 89576 57462
rect 89640 3942 89668 57616
rect 89732 57594 89760 60044
rect 90008 57662 90036 60044
rect 89996 57656 90048 57662
rect 89996 57598 90048 57604
rect 89720 57588 89772 57594
rect 89720 57530 89772 57536
rect 90284 55214 90312 60044
rect 90652 57526 90680 60044
rect 90732 57656 90784 57662
rect 90928 57644 90956 60044
rect 90732 57598 90784 57604
rect 90836 57616 90956 57644
rect 90640 57520 90692 57526
rect 90640 57462 90692 57468
rect 90284 55186 90680 55214
rect 89628 3936 89680 3942
rect 89628 3878 89680 3884
rect 90652 3874 90680 55186
rect 90744 4078 90772 57598
rect 90732 4072 90784 4078
rect 90732 4014 90784 4020
rect 90640 3868 90692 3874
rect 90640 3810 90692 3816
rect 90836 3738 90864 57616
rect 91008 57588 91060 57594
rect 91008 57530 91060 57536
rect 90916 57520 90968 57526
rect 90916 57462 90968 57468
rect 90928 3806 90956 57462
rect 91020 4146 91048 57530
rect 91204 57186 91232 60044
rect 91480 57662 91508 60044
rect 91848 57866 91876 60044
rect 91836 57860 91888 57866
rect 91836 57802 91888 57808
rect 91468 57656 91520 57662
rect 91468 57598 91520 57604
rect 91192 57180 91244 57186
rect 91192 57122 91244 57128
rect 92124 55214 92152 60044
rect 92400 57746 92428 60044
rect 92676 57798 92704 60044
rect 92308 57718 92428 57746
rect 92664 57792 92716 57798
rect 92664 57734 92716 57740
rect 92308 57050 92336 57718
rect 92388 57656 92440 57662
rect 92388 57598 92440 57604
rect 92296 57044 92348 57050
rect 92296 56986 92348 56992
rect 92124 55186 92336 55214
rect 92308 4282 92336 55186
rect 92296 4276 92348 4282
rect 92296 4218 92348 4224
rect 91008 4140 91060 4146
rect 91008 4082 91060 4088
rect 90916 3800 90968 3806
rect 90916 3742 90968 3748
rect 90364 3732 90416 3738
rect 90364 3674 90416 3680
rect 90824 3732 90876 3738
rect 90824 3674 90876 3680
rect 89536 3256 89588 3262
rect 89536 3198 89588 3204
rect 90376 480 90404 3674
rect 92400 3670 92428 57598
rect 93044 57526 93072 60044
rect 93320 57662 93348 60044
rect 93308 57656 93360 57662
rect 93596 57644 93624 60044
rect 93596 57616 93808 57644
rect 93308 57598 93360 57604
rect 93032 57520 93084 57526
rect 93032 57462 93084 57468
rect 93676 57520 93728 57526
rect 93676 57462 93728 57468
rect 92664 57384 92716 57390
rect 92664 57326 92716 57332
rect 92676 16574 92704 57326
rect 92676 16546 92796 16574
rect 92388 3664 92440 3670
rect 92388 3606 92440 3612
rect 91560 3596 91612 3602
rect 91560 3538 91612 3544
rect 91572 480 91600 3538
rect 92768 480 92796 16546
rect 93688 6322 93716 57462
rect 93676 6316 93728 6322
rect 93676 6258 93728 6264
rect 93780 4350 93808 57616
rect 93872 57526 93900 60044
rect 93860 57520 93912 57526
rect 93860 57462 93912 57468
rect 94240 56914 94268 60044
rect 94516 57594 94544 60044
rect 94504 57588 94556 57594
rect 94504 57530 94556 57536
rect 94228 56908 94280 56914
rect 94228 56850 94280 56856
rect 94792 55214 94820 60044
rect 95068 57610 95096 60044
rect 95436 57934 95464 60044
rect 95332 57928 95384 57934
rect 95332 57870 95384 57876
rect 95424 57928 95476 57934
rect 95424 57870 95476 57876
rect 94976 57582 95096 57610
rect 95148 57588 95200 57594
rect 94976 57118 95004 57582
rect 95148 57530 95200 57536
rect 95056 57520 95108 57526
rect 95056 57462 95108 57468
rect 94964 57112 95016 57118
rect 94964 57054 95016 57060
rect 94792 55186 95004 55214
rect 94976 7954 95004 55186
rect 94964 7948 95016 7954
rect 94964 7890 95016 7896
rect 95068 6254 95096 57462
rect 95056 6248 95108 6254
rect 95056 6190 95108 6196
rect 93952 6180 94004 6186
rect 93952 6122 94004 6128
rect 93768 4344 93820 4350
rect 93768 4286 93820 4292
rect 93964 480 93992 6122
rect 95160 4418 95188 57530
rect 95344 56982 95372 57870
rect 95712 57526 95740 60044
rect 95988 57594 96016 60044
rect 96356 57610 96384 60044
rect 95976 57588 96028 57594
rect 96356 57582 96476 57610
rect 95976 57530 96028 57536
rect 95700 57520 95752 57526
rect 95700 57462 95752 57468
rect 96344 57520 96396 57526
rect 96344 57462 96396 57468
rect 95332 56976 95384 56982
rect 95332 56918 95384 56924
rect 96356 7886 96384 57462
rect 96344 7880 96396 7886
rect 96344 7822 96396 7828
rect 96448 4486 96476 57582
rect 96528 57588 96580 57594
rect 96528 57530 96580 57536
rect 96436 4480 96488 4486
rect 96436 4422 96488 4428
rect 95148 4412 95200 4418
rect 95148 4354 95200 4360
rect 96540 3534 96568 57530
rect 96632 57526 96660 60044
rect 96620 57520 96672 57526
rect 96620 57462 96672 57468
rect 96908 57458 96936 60044
rect 97184 57594 97212 60044
rect 97172 57588 97224 57594
rect 97172 57530 97224 57536
rect 96896 57452 96948 57458
rect 96896 57394 96948 57400
rect 97552 57390 97580 60044
rect 97828 57610 97856 60044
rect 97724 57588 97776 57594
rect 97828 57582 97948 57610
rect 97724 57530 97776 57536
rect 97632 57520 97684 57526
rect 97632 57462 97684 57468
rect 97540 57384 97592 57390
rect 97540 57326 97592 57332
rect 97264 57180 97316 57186
rect 97264 57122 97316 57128
rect 97276 8498 97304 57122
rect 97264 8492 97316 8498
rect 97264 8434 97316 8440
rect 97644 7818 97672 57462
rect 97632 7812 97684 7818
rect 97632 7754 97684 7760
rect 97448 7676 97500 7682
rect 97448 7618 97500 7624
rect 95148 3528 95200 3534
rect 95148 3470 95200 3476
rect 96528 3528 96580 3534
rect 96528 3470 96580 3476
rect 95160 480 95188 3470
rect 96252 3324 96304 3330
rect 96252 3266 96304 3272
rect 96264 480 96292 3266
rect 97460 480 97488 7618
rect 97736 4554 97764 57530
rect 97816 57452 97868 57458
rect 97816 57394 97868 57400
rect 97724 4548 97776 4554
rect 97724 4490 97776 4496
rect 97828 3602 97856 57394
rect 97920 4049 97948 57582
rect 98104 57458 98132 60044
rect 98092 57452 98144 57458
rect 98092 57394 98144 57400
rect 98380 57186 98408 60044
rect 98368 57180 98420 57186
rect 98368 57122 98420 57128
rect 98748 56642 98776 60044
rect 99024 57610 99052 60044
rect 98920 57588 98972 57594
rect 99024 57582 99144 57610
rect 99300 57594 99328 60044
rect 98920 57530 98972 57536
rect 98736 56636 98788 56642
rect 98736 56578 98788 56584
rect 98932 7682 98960 57530
rect 99012 57180 99064 57186
rect 99012 57122 99064 57128
rect 99024 7750 99052 57122
rect 99012 7744 99064 7750
rect 99012 7686 99064 7692
rect 98920 7676 98972 7682
rect 98920 7618 98972 7624
rect 98828 7608 98880 7614
rect 98828 7550 98880 7556
rect 97906 4040 97962 4049
rect 97906 3975 97962 3984
rect 97816 3596 97868 3602
rect 97816 3538 97868 3544
rect 98840 3534 98868 7550
rect 99116 4622 99144 57582
rect 99288 57588 99340 57594
rect 99288 57530 99340 57536
rect 99288 57452 99340 57458
rect 99288 57394 99340 57400
rect 99196 56636 99248 56642
rect 99196 56578 99248 56584
rect 99104 4616 99156 4622
rect 99104 4558 99156 4564
rect 99208 3913 99236 56578
rect 99194 3904 99250 3913
rect 99194 3839 99250 3848
rect 98460 3528 98512 3534
rect 98460 3470 98512 3476
rect 98828 3528 98880 3534
rect 98828 3470 98880 3476
rect 98472 2786 98500 3470
rect 99196 3460 99248 3466
rect 99196 3402 99248 3408
rect 98644 2848 98696 2854
rect 98644 2790 98696 2796
rect 98460 2780 98512 2786
rect 98460 2722 98512 2728
rect 98656 480 98684 2790
rect 99208 1018 99236 3402
rect 99300 3233 99328 57394
rect 99576 56710 99604 60044
rect 99564 56704 99616 56710
rect 99564 56646 99616 56652
rect 99944 56642 99972 60044
rect 99932 56636 99984 56642
rect 99932 56578 99984 56584
rect 100220 51074 100248 60044
rect 100392 56636 100444 56642
rect 100392 56578 100444 56584
rect 100404 55026 100432 56578
rect 100496 55162 100524 60044
rect 100668 56704 100720 56710
rect 100668 56646 100720 56652
rect 100496 55134 100616 55162
rect 100404 54998 100524 55026
rect 100220 51046 100432 51074
rect 100404 7614 100432 51046
rect 100392 7608 100444 7614
rect 100392 7550 100444 7556
rect 100496 4690 100524 54998
rect 100484 4684 100536 4690
rect 100484 4626 100536 4632
rect 100588 3641 100616 55134
rect 100574 3632 100630 3641
rect 99392 3590 99604 3618
rect 99286 3224 99342 3233
rect 99286 3159 99342 3168
rect 99392 2854 99420 3590
rect 99576 3466 99604 3590
rect 100680 3602 100708 56646
rect 100772 55350 100800 60044
rect 101140 56710 101168 60044
rect 101312 57316 101364 57322
rect 101312 57258 101364 57264
rect 101128 56704 101180 56710
rect 101128 56646 101180 56652
rect 100760 55344 100812 55350
rect 100760 55286 100812 55292
rect 101324 51074 101352 57258
rect 101416 55570 101444 60044
rect 101692 56642 101720 60044
rect 101968 56794 101996 60044
rect 101784 56766 101996 56794
rect 101680 56636 101732 56642
rect 101680 56578 101732 56584
rect 101416 55542 101720 55570
rect 101324 51046 101444 51074
rect 101416 3602 101444 51046
rect 101692 9450 101720 55542
rect 101680 9444 101732 9450
rect 101680 9386 101732 9392
rect 101784 5506 101812 56766
rect 102336 56710 102364 60044
rect 102612 57322 102640 60044
rect 102600 57316 102652 57322
rect 102600 57258 102652 57264
rect 102784 56976 102836 56982
rect 102784 56918 102836 56924
rect 101864 56704 101916 56710
rect 101864 56646 101916 56652
rect 102324 56704 102376 56710
rect 102324 56646 102376 56652
rect 101772 5500 101824 5506
rect 101772 5442 101824 5448
rect 101876 4758 101904 56646
rect 102048 56636 102100 56642
rect 102048 56578 102100 56584
rect 102060 55434 102088 56578
rect 101968 55406 102088 55434
rect 101864 4752 101916 4758
rect 101864 4694 101916 4700
rect 100574 3567 100630 3576
rect 100668 3596 100720 3602
rect 100668 3538 100720 3544
rect 101404 3596 101456 3602
rect 101404 3538 101456 3544
rect 101220 3528 101272 3534
rect 100128 3466 100340 3482
rect 101496 3528 101548 3534
rect 101272 3476 101496 3482
rect 101968 3505 101996 55406
rect 102048 55344 102100 55350
rect 102048 55286 102100 55292
rect 102060 3777 102088 55286
rect 102796 5302 102824 56918
rect 102888 56642 102916 60044
rect 102968 57248 103020 57254
rect 102968 57190 103020 57196
rect 102876 56636 102928 56642
rect 102876 56578 102928 56584
rect 102980 51074 103008 57190
rect 103060 56704 103112 56710
rect 103060 56646 103112 56652
rect 102888 51046 103008 51074
rect 103072 51074 103100 56646
rect 103164 54482 103192 60044
rect 103532 57186 103560 60044
rect 103520 57180 103572 57186
rect 103520 57122 103572 57128
rect 103428 56636 103480 56642
rect 103428 56578 103480 56584
rect 103164 54454 103376 54482
rect 103072 51046 103284 51074
rect 102784 5296 102836 5302
rect 102784 5238 102836 5244
rect 102046 3768 102102 3777
rect 102046 3703 102102 3712
rect 101220 3470 101548 3476
rect 101954 3496 102010 3505
rect 99564 3460 99616 3466
rect 99564 3402 99616 3408
rect 100116 3460 100352 3466
rect 100168 3454 100300 3460
rect 100116 3402 100168 3408
rect 101232 3454 101536 3470
rect 102888 3466 102916 51046
rect 103256 9382 103284 51046
rect 103244 9376 103296 9382
rect 103244 9318 103296 9324
rect 103348 9314 103376 54454
rect 103336 9308 103388 9314
rect 103336 9250 103388 9256
rect 103440 5438 103468 56578
rect 103808 55486 103836 60044
rect 103980 57928 104032 57934
rect 103980 57870 104032 57876
rect 103888 57724 103940 57730
rect 103888 57666 103940 57672
rect 103796 55480 103848 55486
rect 103796 55422 103848 55428
rect 103900 51074 103928 57666
rect 103992 57458 104020 57870
rect 103980 57452 104032 57458
rect 103980 57394 104032 57400
rect 104084 56642 104112 60044
rect 104256 57588 104308 57594
rect 104256 57530 104308 57536
rect 104164 57520 104216 57526
rect 104164 57462 104216 57468
rect 104176 57118 104204 57462
rect 104164 57112 104216 57118
rect 104164 57054 104216 57060
rect 104268 56914 104296 57530
rect 104256 56908 104308 56914
rect 104256 56850 104308 56856
rect 104360 56710 104388 60044
rect 104348 56704 104400 56710
rect 104348 56646 104400 56652
rect 104072 56636 104124 56642
rect 104072 56578 104124 56584
rect 104532 56636 104584 56642
rect 104532 56578 104584 56584
rect 103900 51046 104204 51074
rect 103704 8492 103756 8498
rect 103704 8434 103756 8440
rect 103428 5432 103480 5438
rect 103428 5374 103480 5380
rect 103428 5296 103480 5302
rect 103428 5238 103480 5244
rect 103440 3602 103468 5238
rect 103336 3596 103388 3602
rect 103336 3538 103388 3544
rect 103428 3596 103480 3602
rect 103428 3538 103480 3544
rect 101954 3431 102010 3440
rect 102324 3460 102376 3466
rect 100300 3402 100352 3408
rect 102324 3402 102376 3408
rect 102876 3460 102928 3466
rect 102876 3402 102928 3408
rect 101036 3392 101088 3398
rect 101036 3334 101088 3340
rect 99380 2848 99432 2854
rect 99380 2790 99432 2796
rect 99196 1012 99248 1018
rect 99196 954 99248 960
rect 99840 1012 99892 1018
rect 99840 954 99892 960
rect 99852 480 99880 954
rect 101048 480 101076 3334
rect 102336 2922 102364 3402
rect 102232 2916 102284 2922
rect 102232 2858 102284 2864
rect 102324 2916 102376 2922
rect 102324 2858 102376 2864
rect 102244 480 102272 2858
rect 103348 480 103376 3538
rect 103716 2922 103744 8434
rect 104176 5114 104204 51046
rect 104544 9246 104572 56578
rect 104728 55570 104756 60044
rect 105004 56710 105032 60044
rect 105280 56778 105308 60044
rect 105268 56772 105320 56778
rect 105268 56714 105320 56720
rect 104808 56704 104860 56710
rect 104808 56646 104860 56652
rect 104992 56704 105044 56710
rect 104992 56646 105044 56652
rect 104636 55542 104756 55570
rect 104532 9240 104584 9246
rect 104532 9182 104584 9188
rect 104636 5302 104664 55542
rect 104716 55480 104768 55486
rect 104716 55422 104768 55428
rect 104728 5370 104756 55422
rect 104716 5364 104768 5370
rect 104716 5306 104768 5312
rect 104624 5296 104676 5302
rect 104624 5238 104676 5244
rect 104176 5086 104664 5114
rect 104636 2990 104664 5086
rect 104820 3369 104848 56646
rect 105556 56642 105584 60044
rect 105820 56704 105872 56710
rect 105820 56646 105872 56652
rect 105544 56636 105596 56642
rect 105544 56578 105596 56584
rect 105832 51074 105860 56646
rect 105924 55570 105952 60044
rect 106200 57118 106228 60044
rect 106188 57112 106240 57118
rect 106188 57054 106240 57060
rect 106188 56772 106240 56778
rect 106188 56714 106240 56720
rect 106096 56636 106148 56642
rect 106096 56578 106148 56584
rect 105924 55542 106044 55570
rect 105832 51046 105952 51074
rect 105924 9178 105952 51046
rect 105912 9172 105964 9178
rect 105912 9114 105964 9120
rect 106016 9110 106044 55542
rect 106004 9104 106056 9110
rect 106004 9046 106056 9052
rect 106108 5234 106136 56578
rect 106096 5228 106148 5234
rect 106096 5170 106148 5176
rect 104806 3360 104862 3369
rect 104806 3295 104862 3304
rect 106200 3126 106228 56714
rect 106476 56710 106504 60044
rect 106464 56704 106516 56710
rect 106464 56646 106516 56652
rect 106752 56642 106780 60044
rect 107120 57934 107148 60044
rect 107108 57928 107160 57934
rect 107108 57870 107160 57876
rect 106740 56636 106792 56642
rect 106740 56578 106792 56584
rect 107396 8974 107424 60044
rect 107568 56704 107620 56710
rect 107568 56646 107620 56652
rect 107476 56636 107528 56642
rect 107476 56578 107528 56584
rect 107488 9042 107516 56578
rect 107476 9036 107528 9042
rect 107476 8978 107528 8984
rect 107384 8968 107436 8974
rect 107384 8910 107436 8916
rect 107580 5166 107608 56646
rect 107672 56642 107700 60044
rect 107660 56636 107712 56642
rect 107660 56578 107712 56584
rect 108040 51882 108068 60044
rect 108028 51876 108080 51882
rect 108028 51818 108080 51824
rect 108316 51074 108344 60044
rect 108488 56636 108540 56642
rect 108488 56578 108540 56584
rect 108500 55434 108528 56578
rect 108592 55570 108620 60044
rect 108868 55570 108896 60044
rect 109236 56710 109264 60044
rect 109512 56846 109540 60044
rect 109500 56840 109552 56846
rect 109500 56782 109552 56788
rect 109788 56778 109816 60044
rect 109776 56772 109828 56778
rect 109776 56714 109828 56720
rect 109224 56704 109276 56710
rect 109224 56646 109276 56652
rect 109960 56704 110012 56710
rect 109960 56646 110012 56652
rect 108592 55542 108804 55570
rect 108868 55542 108988 55570
rect 108500 55406 108712 55434
rect 108316 51046 108620 51074
rect 108592 10878 108620 51046
rect 108684 10946 108712 55406
rect 108672 10940 108724 10946
rect 108672 10882 108724 10888
rect 108580 10872 108632 10878
rect 108580 10814 108632 10820
rect 108776 10810 108804 55542
rect 108856 51876 108908 51882
rect 108856 51818 108908 51824
rect 108764 10804 108816 10810
rect 108764 10746 108816 10752
rect 107568 5160 107620 5166
rect 107568 5102 107620 5108
rect 108868 5098 108896 51818
rect 108856 5092 108908 5098
rect 108856 5034 108908 5040
rect 108960 5030 108988 55542
rect 109972 51074 110000 56646
rect 110064 53666 110092 60044
rect 110236 56840 110288 56846
rect 110236 56782 110288 56788
rect 110064 53638 110184 53666
rect 109972 51046 110092 51074
rect 110064 10742 110092 51046
rect 110052 10736 110104 10742
rect 110052 10678 110104 10684
rect 110156 10606 110184 53638
rect 110248 10674 110276 56782
rect 110432 56778 110460 60044
rect 110708 56846 110736 60044
rect 110696 56840 110748 56846
rect 110696 56782 110748 56788
rect 110328 56772 110380 56778
rect 110328 56714 110380 56720
rect 110420 56772 110472 56778
rect 110420 56714 110472 56720
rect 110236 10668 110288 10674
rect 110236 10610 110288 10616
rect 110144 10600 110196 10606
rect 110144 10542 110196 10548
rect 108948 5024 109000 5030
rect 108948 4966 109000 4972
rect 110340 4962 110368 56714
rect 110984 56710 111012 60044
rect 110972 56704 111024 56710
rect 110972 56646 111024 56652
rect 111260 51074 111288 60044
rect 111432 56772 111484 56778
rect 111432 56714 111484 56720
rect 111260 51046 111380 51074
rect 111352 10402 111380 51046
rect 111444 10538 111472 56714
rect 111524 56704 111576 56710
rect 111524 56646 111576 56652
rect 111432 10532 111484 10538
rect 111432 10474 111484 10480
rect 111536 10470 111564 56646
rect 111524 10464 111576 10470
rect 111524 10406 111576 10412
rect 111340 10396 111392 10402
rect 111340 10338 111392 10344
rect 110328 4956 110380 4962
rect 110328 4898 110380 4904
rect 111628 4826 111656 60044
rect 111904 56846 111932 60044
rect 111708 56840 111760 56846
rect 111708 56782 111760 56788
rect 111892 56840 111944 56846
rect 111892 56782 111944 56788
rect 111720 4894 111748 56782
rect 112180 56778 112208 60044
rect 112168 56772 112220 56778
rect 112168 56714 112220 56720
rect 112456 55554 112484 60044
rect 112720 56704 112772 56710
rect 112720 56646 112772 56652
rect 112444 55548 112496 55554
rect 112444 55490 112496 55496
rect 112732 15366 112760 56646
rect 112720 15360 112772 15366
rect 112720 15302 112772 15308
rect 112824 9790 112852 60044
rect 112904 56840 112956 56846
rect 112904 56782 112956 56788
rect 112916 10334 112944 56782
rect 112996 56772 113048 56778
rect 112996 56714 113048 56720
rect 112904 10328 112956 10334
rect 112904 10270 112956 10276
rect 112812 9784 112864 9790
rect 112812 9726 112864 9732
rect 111708 4888 111760 4894
rect 111708 4830 111760 4836
rect 111616 4820 111668 4826
rect 111616 4762 111668 4768
rect 111616 4004 111668 4010
rect 111616 3946 111668 3952
rect 106844 3602 107148 3618
rect 106832 3596 107148 3602
rect 106884 3590 107148 3596
rect 106832 3538 106884 3544
rect 106924 3460 106976 3466
rect 106924 3402 106976 3408
rect 105728 3120 105780 3126
rect 105728 3062 105780 3068
rect 106188 3120 106240 3126
rect 106188 3062 106240 3068
rect 104532 2984 104584 2990
rect 104532 2926 104584 2932
rect 104624 2984 104676 2990
rect 104624 2926 104676 2932
rect 103612 2916 103664 2922
rect 103612 2858 103664 2864
rect 103704 2916 103756 2922
rect 103704 2858 103756 2864
rect 103624 2802 103652 2858
rect 103888 2848 103940 2854
rect 103624 2796 103888 2802
rect 103624 2790 103940 2796
rect 103624 2774 103928 2790
rect 104544 480 104572 2926
rect 105740 480 105768 3062
rect 106936 480 106964 3402
rect 107120 3398 107148 3590
rect 107476 3596 107528 3602
rect 107212 3556 107476 3584
rect 107016 3392 107068 3398
rect 107016 3334 107068 3340
rect 107108 3392 107160 3398
rect 107108 3334 107160 3340
rect 107028 3244 107056 3334
rect 107212 3244 107240 3556
rect 107476 3538 107528 3544
rect 110144 3460 110196 3466
rect 110144 3402 110196 3408
rect 107028 3216 107240 3244
rect 109316 3188 109368 3194
rect 109316 3130 109368 3136
rect 108120 3052 108172 3058
rect 108120 2994 108172 3000
rect 108132 480 108160 2994
rect 109328 480 109356 3130
rect 110156 2854 110184 3402
rect 110512 3392 110564 3398
rect 110512 3334 110564 3340
rect 110604 3392 110656 3398
rect 110604 3334 110656 3340
rect 110144 2848 110196 2854
rect 110144 2790 110196 2796
rect 110524 480 110552 3334
rect 110616 2922 110644 3334
rect 110604 2916 110656 2922
rect 110604 2858 110656 2864
rect 111628 480 111656 3946
rect 113008 3262 113036 56714
rect 113100 56710 113128 60044
rect 113376 56982 113404 60044
rect 113364 56976 113416 56982
rect 113364 56918 113416 56924
rect 113652 56710 113680 60044
rect 113732 57860 113784 57866
rect 113732 57802 113784 57808
rect 113744 56846 113772 57802
rect 113824 57724 113876 57730
rect 113824 57666 113876 57672
rect 113836 57118 113864 57666
rect 113824 57112 113876 57118
rect 113824 57054 113876 57060
rect 113732 56840 113784 56846
rect 113732 56782 113784 56788
rect 113088 56704 113140 56710
rect 113088 56646 113140 56652
rect 113640 56704 113692 56710
rect 113640 56646 113692 56652
rect 113088 55548 113140 55554
rect 113088 55490 113140 55496
rect 113100 4010 113128 55490
rect 114020 51074 114048 60044
rect 114296 57186 114324 60044
rect 114284 57180 114336 57186
rect 114284 57122 114336 57128
rect 114572 56778 114600 60044
rect 114560 56772 114612 56778
rect 114560 56714 114612 56720
rect 114848 56710 114876 60044
rect 114468 56704 114520 56710
rect 114468 56646 114520 56652
rect 114836 56704 114888 56710
rect 114836 56646 114888 56652
rect 114020 51046 114416 51074
rect 114388 15434 114416 51046
rect 114376 15428 114428 15434
rect 114376 15370 114428 15376
rect 114480 9858 114508 56646
rect 115216 55622 115244 60044
rect 115492 56914 115520 60044
rect 115480 56908 115532 56914
rect 115480 56850 115532 56856
rect 115480 56772 115532 56778
rect 115480 56714 115532 56720
rect 115204 55616 115256 55622
rect 115204 55558 115256 55564
rect 115492 9926 115520 56714
rect 115572 56704 115624 56710
rect 115572 56646 115624 56652
rect 115584 15502 115612 56646
rect 115768 55570 115796 60044
rect 115848 56908 115900 56914
rect 115848 56850 115900 56856
rect 115676 55542 115796 55570
rect 115676 15570 115704 55542
rect 115860 51074 115888 56850
rect 116044 55690 116072 60044
rect 116412 56710 116440 60044
rect 116688 56778 116716 60044
rect 116676 56772 116728 56778
rect 116676 56714 116728 56720
rect 116400 56704 116452 56710
rect 116400 56646 116452 56652
rect 116860 56704 116912 56710
rect 116860 56646 116912 56652
rect 116032 55684 116084 55690
rect 116032 55626 116084 55632
rect 115768 51046 115888 51074
rect 115664 15564 115716 15570
rect 115664 15506 115716 15512
rect 115572 15496 115624 15502
rect 115572 15438 115624 15444
rect 115768 9994 115796 51046
rect 116872 10062 116900 56646
rect 116964 17134 116992 60044
rect 117044 56772 117096 56778
rect 117044 56714 117096 56720
rect 116952 17128 117004 17134
rect 116952 17070 117004 17076
rect 117056 15638 117084 56714
rect 117240 45554 117268 60044
rect 117608 57118 117636 60044
rect 117596 57112 117648 57118
rect 117596 57054 117648 57060
rect 117884 56574 117912 60044
rect 118160 57866 118188 60044
rect 118148 57860 118200 57866
rect 118148 57802 118200 57808
rect 117872 56568 117924 56574
rect 117872 56510 117924 56516
rect 117148 45526 117268 45554
rect 117044 15632 117096 15638
rect 117044 15574 117096 15580
rect 117148 10130 117176 45526
rect 118436 15774 118464 60044
rect 118608 57860 118660 57866
rect 118608 57802 118660 57808
rect 118516 57112 118568 57118
rect 118516 57054 118568 57060
rect 118424 15768 118476 15774
rect 118424 15710 118476 15716
rect 118528 15706 118556 57054
rect 118516 15700 118568 15706
rect 118516 15642 118568 15648
rect 118620 10198 118648 57802
rect 118804 55758 118832 60044
rect 118792 55752 118844 55758
rect 118792 55694 118844 55700
rect 119080 52902 119108 60044
rect 119356 55486 119384 60044
rect 119344 55480 119396 55486
rect 119344 55422 119396 55428
rect 119068 52896 119120 52902
rect 119068 52838 119120 52844
rect 118608 10192 118660 10198
rect 118608 10134 118660 10140
rect 117136 10124 117188 10130
rect 117136 10066 117188 10072
rect 116860 10056 116912 10062
rect 116860 9998 116912 10004
rect 115756 9988 115808 9994
rect 115756 9930 115808 9936
rect 115480 9920 115532 9926
rect 115480 9862 115532 9868
rect 114468 9852 114520 9858
rect 114468 9794 114520 9800
rect 119724 5574 119752 60044
rect 120000 55570 120028 60044
rect 120276 56778 120304 60044
rect 120264 56772 120316 56778
rect 120264 56714 120316 56720
rect 120552 56642 120580 60044
rect 120920 57866 120948 60044
rect 120908 57860 120960 57866
rect 120908 57802 120960 57808
rect 120540 56636 120592 56642
rect 120540 56578 120592 56584
rect 119816 55542 120028 55570
rect 119816 18698 119844 55542
rect 119896 55480 119948 55486
rect 119896 55422 119948 55428
rect 119804 18692 119856 18698
rect 119804 18634 119856 18640
rect 119908 15842 119936 55422
rect 121196 16522 121224 60044
rect 121276 56772 121328 56778
rect 121276 56714 121328 56720
rect 121288 16590 121316 56714
rect 121472 56642 121500 60044
rect 121748 57050 121776 60044
rect 121736 57044 121788 57050
rect 121736 56986 121788 56992
rect 121368 56636 121420 56642
rect 121368 56578 121420 56584
rect 121460 56636 121512 56642
rect 121460 56578 121512 56584
rect 121276 16584 121328 16590
rect 121276 16526 121328 16532
rect 121184 16516 121236 16522
rect 121184 16458 121236 16464
rect 119896 15836 119948 15842
rect 119896 15778 119948 15784
rect 121380 5642 121408 56578
rect 122012 56500 122064 56506
rect 122012 56442 122064 56448
rect 122024 48314 122052 56442
rect 122116 55434 122144 60044
rect 122392 55570 122420 60044
rect 122668 56982 122696 60044
rect 122656 56976 122708 56982
rect 122656 56918 122708 56924
rect 122944 56642 122972 60044
rect 122748 56636 122800 56642
rect 122748 56578 122800 56584
rect 122932 56636 122984 56642
rect 122932 56578 122984 56584
rect 122392 55542 122696 55570
rect 122116 55406 122604 55434
rect 122024 48286 122144 48314
rect 121368 5636 121420 5642
rect 121368 5578 121420 5584
rect 119712 5568 119764 5574
rect 119712 5510 119764 5516
rect 117596 4140 117648 4146
rect 117596 4082 117648 4088
rect 113088 4004 113140 4010
rect 113088 3946 113140 3952
rect 116400 3936 116452 3942
rect 116400 3878 116452 3884
rect 115204 3324 115256 3330
rect 115204 3266 115256 3272
rect 112812 3256 112864 3262
rect 112812 3198 112864 3204
rect 112996 3256 113048 3262
rect 112996 3198 113048 3204
rect 112824 480 112852 3198
rect 114008 2984 114060 2990
rect 114008 2926 114060 2932
rect 114020 480 114048 2926
rect 115216 480 115244 3266
rect 116412 480 116440 3878
rect 117608 480 117636 4082
rect 118792 4072 118844 4078
rect 118792 4014 118844 4020
rect 118804 480 118832 4014
rect 119896 3868 119948 3874
rect 119896 3810 119948 3816
rect 119908 480 119936 3810
rect 122116 3806 122144 48286
rect 122576 16454 122604 55406
rect 122564 16448 122616 16454
rect 122564 16390 122616 16396
rect 122668 5778 122696 55542
rect 122656 5772 122708 5778
rect 122656 5714 122708 5720
rect 122760 5710 122788 56578
rect 123312 50386 123340 60044
rect 123588 56846 123616 60044
rect 123576 56840 123628 56846
rect 123576 56782 123628 56788
rect 123760 56636 123812 56642
rect 123760 56578 123812 56584
rect 123772 51074 123800 56578
rect 123864 55570 123892 60044
rect 123864 55542 123984 55570
rect 123772 51046 123892 51074
rect 123300 50380 123352 50386
rect 123300 50322 123352 50328
rect 123864 16386 123892 51046
rect 123852 16380 123904 16386
rect 123852 16322 123904 16328
rect 123956 16318 123984 55542
rect 124140 51074 124168 60044
rect 124508 52970 124536 60044
rect 124784 56642 124812 60044
rect 124864 56908 124916 56914
rect 124864 56850 124916 56856
rect 124772 56636 124824 56642
rect 124772 56578 124824 56584
rect 124496 52964 124548 52970
rect 124496 52906 124548 52912
rect 124048 51046 124168 51074
rect 123944 16312 123996 16318
rect 123944 16254 123996 16260
rect 124048 5914 124076 51046
rect 124128 50380 124180 50386
rect 124128 50322 124180 50328
rect 124036 5908 124088 5914
rect 124036 5850 124088 5856
rect 124140 5846 124168 50322
rect 124128 5840 124180 5846
rect 124128 5782 124180 5788
rect 122748 5704 122800 5710
rect 122748 5646 122800 5652
rect 121092 3800 121144 3806
rect 121092 3742 121144 3748
rect 122104 3800 122156 3806
rect 122104 3742 122156 3748
rect 121104 480 121132 3742
rect 122288 3732 122340 3738
rect 122288 3674 122340 3680
rect 122300 480 122328 3674
rect 124680 3664 124732 3670
rect 124680 3606 124732 3612
rect 123484 3392 123536 3398
rect 123484 3334 123536 3340
rect 123496 480 123524 3334
rect 124692 480 124720 3606
rect 124876 3398 124904 56850
rect 125060 51074 125088 60044
rect 125336 53038 125364 60044
rect 125704 56642 125732 60044
rect 125980 56778 126008 60044
rect 126256 58562 126284 60044
rect 126256 58534 126468 58562
rect 126440 57866 126468 58534
rect 126428 57860 126480 57866
rect 126428 57802 126480 57808
rect 126244 57792 126296 57798
rect 126244 57734 126296 57740
rect 125968 56772 126020 56778
rect 125968 56714 126020 56720
rect 125416 56636 125468 56642
rect 125416 56578 125468 56584
rect 125692 56636 125744 56642
rect 125692 56578 125744 56584
rect 125324 53032 125376 53038
rect 125324 52974 125376 52980
rect 125060 51046 125272 51074
rect 125244 5982 125272 51046
rect 125428 16250 125456 56578
rect 126256 51074 126284 57734
rect 126428 56636 126480 56642
rect 126428 56578 126480 56584
rect 126440 51074 126468 56578
rect 126532 55570 126560 60044
rect 126796 56772 126848 56778
rect 126796 56714 126848 56720
rect 126532 55542 126744 55570
rect 126256 51046 126376 51074
rect 126440 51046 126652 51074
rect 125416 16244 125468 16250
rect 125416 16186 125468 16192
rect 125232 5976 125284 5982
rect 125232 5918 125284 5924
rect 124864 3392 124916 3398
rect 124864 3334 124916 3340
rect 125876 3392 125928 3398
rect 125876 3334 125928 3340
rect 125888 480 125916 3334
rect 126348 3194 126376 51046
rect 126624 16182 126652 51046
rect 126612 16176 126664 16182
rect 126612 16118 126664 16124
rect 126716 16114 126744 55542
rect 126704 16108 126756 16114
rect 126704 16050 126756 16056
rect 126808 6050 126836 56714
rect 126900 6118 126928 60044
rect 127176 56642 127204 60044
rect 127452 56642 127480 60044
rect 127728 57746 127756 60044
rect 127728 57718 128032 57746
rect 128004 57662 128032 57718
rect 127900 57656 127952 57662
rect 127900 57598 127952 57604
rect 127992 57656 128044 57662
rect 127992 57598 128044 57604
rect 127806 57080 127862 57089
rect 127716 57044 127768 57050
rect 127806 57015 127862 57024
rect 127716 56986 127768 56992
rect 127728 56846 127756 56986
rect 127820 56982 127848 57015
rect 127808 56976 127860 56982
rect 127808 56918 127860 56924
rect 127716 56840 127768 56846
rect 127716 56782 127768 56788
rect 127164 56636 127216 56642
rect 127164 56578 127216 56584
rect 127440 56636 127492 56642
rect 127440 56578 127492 56584
rect 127912 56574 127940 57598
rect 127992 56636 128044 56642
rect 127992 56578 128044 56584
rect 127256 56568 127308 56574
rect 127256 56510 127308 56516
rect 127900 56568 127952 56574
rect 127900 56510 127952 56516
rect 127268 55554 127296 56510
rect 127256 55548 127308 55554
rect 127256 55490 127308 55496
rect 128004 16046 128032 56578
rect 127992 16040 128044 16046
rect 127992 15982 128044 15988
rect 128096 11218 128124 60044
rect 128176 57656 128228 57662
rect 128176 57598 128228 57604
rect 128188 56658 128216 57598
rect 128372 56914 128400 60044
rect 128452 57792 128504 57798
rect 128452 57734 128504 57740
rect 128464 57050 128492 57734
rect 128452 57044 128504 57050
rect 128452 56986 128504 56992
rect 128360 56908 128412 56914
rect 128360 56850 128412 56856
rect 128188 56630 128308 56658
rect 128176 56500 128228 56506
rect 128176 56442 128228 56448
rect 128084 11212 128136 11218
rect 128084 11154 128136 11160
rect 128188 11150 128216 56442
rect 128176 11144 128228 11150
rect 128176 11086 128228 11092
rect 128280 6866 128308 56630
rect 128648 53446 128676 60044
rect 128924 56642 128952 60044
rect 128912 56636 128964 56642
rect 128912 56578 128964 56584
rect 128636 53440 128688 53446
rect 128636 53382 128688 53388
rect 129292 17814 129320 60044
rect 129372 56908 129424 56914
rect 129372 56850 129424 56856
rect 129384 17882 129412 56850
rect 129464 56636 129516 56642
rect 129464 56578 129516 56584
rect 129372 17876 129424 17882
rect 129372 17818 129424 17824
rect 129280 17808 129332 17814
rect 129280 17750 129332 17756
rect 128268 6860 128320 6866
rect 128268 6802 128320 6808
rect 129476 6798 129504 56578
rect 129568 53530 129596 60044
rect 129844 56710 129872 60044
rect 129832 56704 129884 56710
rect 129832 56646 129884 56652
rect 130120 56642 130148 60044
rect 130108 56636 130160 56642
rect 130108 56578 130160 56584
rect 130488 55350 130516 60044
rect 130660 56636 130712 56642
rect 130660 56578 130712 56584
rect 130476 55344 130528 55350
rect 130476 55286 130528 55292
rect 129568 53502 129688 53530
rect 129556 53440 129608 53446
rect 129556 53382 129608 53388
rect 129464 6792 129516 6798
rect 129464 6734 129516 6740
rect 129568 6186 129596 53382
rect 129660 6730 129688 53502
rect 130672 17746 130700 56578
rect 130764 55570 130792 60044
rect 130936 56704 130988 56710
rect 130936 56646 130988 56652
rect 130764 55542 130884 55570
rect 130752 55480 130804 55486
rect 130752 55422 130804 55428
rect 130660 17740 130712 17746
rect 130660 17682 130712 17688
rect 130764 17678 130792 55422
rect 130752 17672 130804 17678
rect 130752 17614 130804 17620
rect 130856 11354 130884 55542
rect 130844 11348 130896 11354
rect 130844 11290 130896 11296
rect 130948 11286 130976 56646
rect 131040 55486 131068 60044
rect 131408 56710 131436 60044
rect 131396 56704 131448 56710
rect 131396 56646 131448 56652
rect 131684 56642 131712 60044
rect 131856 57588 131908 57594
rect 131856 57530 131908 57536
rect 131868 56914 131896 57530
rect 131856 56908 131908 56914
rect 131856 56850 131908 56856
rect 131120 56636 131172 56642
rect 131120 56578 131172 56584
rect 131672 56636 131724 56642
rect 131672 56578 131724 56584
rect 131028 55480 131080 55486
rect 131028 55422 131080 55428
rect 131028 55344 131080 55350
rect 131028 55286 131080 55292
rect 130936 11280 130988 11286
rect 130936 11222 130988 11228
rect 129648 6724 129700 6730
rect 129648 6666 129700 6672
rect 131040 6662 131068 55286
rect 131132 16574 131160 56578
rect 131960 51074 131988 60044
rect 132040 57588 132092 57594
rect 132040 57530 132092 57536
rect 132052 57458 132080 57530
rect 132040 57452 132092 57458
rect 132040 57394 132092 57400
rect 131960 51046 132172 51074
rect 132144 17610 132172 51046
rect 132132 17604 132184 17610
rect 132132 17546 132184 17552
rect 131132 16546 131804 16574
rect 131028 6656 131080 6662
rect 131028 6598 131080 6604
rect 130568 6316 130620 6322
rect 130568 6258 130620 6264
rect 129556 6180 129608 6186
rect 129556 6122 129608 6128
rect 126888 6112 126940 6118
rect 126888 6054 126940 6060
rect 126796 6044 126848 6050
rect 126796 5986 126848 5992
rect 126980 4276 127032 4282
rect 126980 4218 127032 4224
rect 126336 3188 126388 3194
rect 126336 3130 126388 3136
rect 126992 480 127020 4218
rect 128176 3800 128228 3806
rect 128176 3742 128228 3748
rect 128188 480 128216 3742
rect 129372 3188 129424 3194
rect 129372 3130 129424 3136
rect 129384 480 129412 3130
rect 130580 480 130608 6258
rect 131776 480 131804 16546
rect 132236 6526 132264 60044
rect 132604 56710 132632 60044
rect 132316 56704 132368 56710
rect 132316 56646 132368 56652
rect 132592 56704 132644 56710
rect 132592 56646 132644 56652
rect 132328 6594 132356 56646
rect 132880 56642 132908 60044
rect 132960 57520 133012 57526
rect 132960 57462 133012 57468
rect 132972 57089 133000 57462
rect 132958 57080 133014 57089
rect 132958 57015 133014 57024
rect 133156 56846 133184 60044
rect 133144 56840 133196 56846
rect 133144 56782 133196 56788
rect 133432 56794 133460 60044
rect 133800 57934 133828 60044
rect 133788 57928 133840 57934
rect 133788 57870 133840 57876
rect 134076 56846 134104 60044
rect 133788 56840 133840 56846
rect 133432 56766 133736 56794
rect 133788 56782 133840 56788
rect 134064 56840 134116 56846
rect 134064 56782 134116 56788
rect 133604 56704 133656 56710
rect 133604 56646 133656 56652
rect 132408 56636 132460 56642
rect 132408 56578 132460 56584
rect 132868 56636 132920 56642
rect 132868 56578 132920 56584
rect 133328 56636 133380 56642
rect 133328 56578 133380 56584
rect 132316 6588 132368 6594
rect 132316 6530 132368 6536
rect 132224 6520 132276 6526
rect 132224 6462 132276 6468
rect 132420 3194 132448 56578
rect 133340 51074 133368 56578
rect 133340 51046 133552 51074
rect 133524 17542 133552 51046
rect 133512 17536 133564 17542
rect 133512 17478 133564 17484
rect 133616 11422 133644 56646
rect 133708 11490 133736 56766
rect 133696 11484 133748 11490
rect 133696 11426 133748 11432
rect 133604 11416 133656 11422
rect 133604 11358 133656 11364
rect 133800 6458 133828 56782
rect 134352 56642 134380 60044
rect 134628 56710 134656 60044
rect 134616 56704 134668 56710
rect 134616 56646 134668 56652
rect 134340 56636 134392 56642
rect 134340 56578 134392 56584
rect 134892 56636 134944 56642
rect 134892 56578 134944 56584
rect 134904 11558 134932 56578
rect 134892 11552 134944 11558
rect 134892 11494 134944 11500
rect 133788 6452 133840 6458
rect 133788 6394 133840 6400
rect 134996 6322 135024 60044
rect 135076 56840 135128 56846
rect 135076 56782 135128 56788
rect 135088 6390 135116 56782
rect 135272 56710 135300 60044
rect 135548 57730 135576 60044
rect 135536 57724 135588 57730
rect 135536 57666 135588 57672
rect 135352 56908 135404 56914
rect 135352 56850 135404 56856
rect 135168 56704 135220 56710
rect 135168 56646 135220 56652
rect 135260 56704 135312 56710
rect 135260 56646 135312 56652
rect 135076 6384 135128 6390
rect 135076 6326 135128 6332
rect 134984 6316 135036 6322
rect 134984 6258 135036 6264
rect 134156 6248 134208 6254
rect 134156 6190 134208 6196
rect 132960 4344 133012 4350
rect 132960 4286 133012 4292
rect 132408 3188 132460 3194
rect 132408 3130 132460 3136
rect 132972 480 133000 4286
rect 134168 480 134196 6190
rect 135180 3330 135208 56646
rect 135364 45554 135392 56850
rect 135824 56642 135852 60044
rect 136088 56704 136140 56710
rect 136088 56646 136140 56652
rect 135812 56636 135864 56642
rect 135812 56578 135864 56584
rect 136100 54534 136128 56646
rect 136088 54528 136140 54534
rect 136088 54470 136140 54476
rect 136192 53582 136220 60044
rect 136272 57860 136324 57866
rect 136272 57802 136324 57808
rect 136284 56710 136312 57802
rect 136272 56704 136324 56710
rect 136272 56646 136324 56652
rect 136468 54618 136496 60044
rect 136640 57044 136692 57050
rect 136640 56986 136692 56992
rect 136548 56636 136600 56642
rect 136548 56578 136600 56584
rect 136284 54590 136496 54618
rect 136180 53576 136232 53582
rect 136180 53518 136232 53524
rect 135272 45526 135392 45554
rect 135168 3324 135220 3330
rect 135168 3266 135220 3272
rect 135272 480 135300 45526
rect 136284 17338 136312 54590
rect 136456 54528 136508 54534
rect 136456 54470 136508 54476
rect 136364 53576 136416 53582
rect 136364 53518 136416 53524
rect 136272 17332 136324 17338
rect 136272 17274 136324 17280
rect 136376 11694 136404 53518
rect 136364 11688 136416 11694
rect 136364 11630 136416 11636
rect 136468 11626 136496 54470
rect 136456 11620 136508 11626
rect 136456 11562 136508 11568
rect 136560 6254 136588 56578
rect 136652 52766 136680 56986
rect 136744 54262 136772 60044
rect 137020 56642 137048 60044
rect 137388 57866 137416 60044
rect 137376 57860 137428 57866
rect 137376 57802 137428 57808
rect 137192 57656 137244 57662
rect 137244 57604 137416 57610
rect 137192 57598 137416 57604
rect 137204 57582 137416 57598
rect 137388 57526 137416 57582
rect 137284 57520 137336 57526
rect 137284 57462 137336 57468
rect 137376 57520 137428 57526
rect 137376 57462 137428 57468
rect 137008 56636 137060 56642
rect 137008 56578 137060 56584
rect 136732 54256 136784 54262
rect 136732 54198 136784 54204
rect 136640 52760 136692 52766
rect 136640 52702 136692 52708
rect 137296 17202 137324 57462
rect 137284 17196 137336 17202
rect 137284 17138 137336 17144
rect 137664 11778 137692 60044
rect 137744 56636 137796 56642
rect 137744 56578 137796 56584
rect 137756 12442 137784 56578
rect 137940 51074 137968 60044
rect 138020 57452 138072 57458
rect 138020 57394 138072 57400
rect 137848 51046 137968 51074
rect 137744 12436 137796 12442
rect 137744 12378 137796 12384
rect 137848 12374 137876 51046
rect 138032 16574 138060 57394
rect 138216 56642 138244 60044
rect 138584 56846 138612 60044
rect 138664 57656 138716 57662
rect 138664 57598 138716 57604
rect 138572 56840 138624 56846
rect 138572 56782 138624 56788
rect 138204 56636 138256 56642
rect 138204 56578 138256 56584
rect 138032 16546 138612 16574
rect 137836 12368 137888 12374
rect 137836 12310 137888 12316
rect 137664 11750 137784 11778
rect 137652 7948 137704 7954
rect 137652 7890 137704 7896
rect 136548 6248 136600 6254
rect 136548 6190 136600 6196
rect 136456 4412 136508 4418
rect 136456 4354 136508 4360
rect 136468 480 136496 4354
rect 137664 480 137692 7890
rect 137756 3398 137784 11750
rect 138584 3482 138612 16546
rect 138676 3670 138704 57598
rect 138860 51074 138888 60044
rect 139136 56914 139164 60044
rect 139124 56908 139176 56914
rect 139124 56850 139176 56856
rect 139308 56636 139360 56642
rect 139308 56578 139360 56584
rect 138860 51046 139256 51074
rect 139228 12306 139256 51046
rect 139216 12300 139268 12306
rect 139216 12242 139268 12248
rect 139320 4146 139348 56578
rect 139412 55826 139440 60044
rect 139492 57928 139544 57934
rect 139492 57870 139544 57876
rect 139400 55820 139452 55826
rect 139400 55762 139452 55768
rect 139504 50318 139532 57870
rect 139780 56642 139808 60044
rect 140056 57050 140084 60044
rect 140044 57044 140096 57050
rect 140044 56986 140096 56992
rect 139768 56636 139820 56642
rect 139768 56578 139820 56584
rect 140332 54398 140360 60044
rect 140504 56636 140556 56642
rect 140504 56578 140556 56584
rect 140320 54392 140372 54398
rect 140320 54334 140372 54340
rect 139492 50312 139544 50318
rect 139492 50254 139544 50260
rect 140516 12238 140544 56578
rect 140504 12232 140556 12238
rect 140504 12174 140556 12180
rect 140608 12170 140636 60044
rect 140976 57594 141004 60044
rect 140964 57588 141016 57594
rect 140964 57530 141016 57536
rect 141252 54466 141280 60044
rect 141424 56704 141476 56710
rect 141424 56646 141476 56652
rect 141240 54460 141292 54466
rect 141240 54402 141292 54408
rect 140596 12164 140648 12170
rect 140596 12106 140648 12112
rect 141240 7880 141292 7886
rect 141240 7822 141292 7828
rect 139308 4140 139360 4146
rect 139308 4082 139360 4088
rect 138664 3664 138716 3670
rect 138664 3606 138716 3612
rect 140044 3664 140096 3670
rect 140044 3606 140096 3612
rect 138584 3454 138888 3482
rect 137744 3392 137796 3398
rect 137744 3334 137796 3340
rect 138860 480 138888 3454
rect 140056 480 140084 3606
rect 141252 480 141280 7822
rect 141436 4418 141464 56646
rect 141528 56642 141556 60044
rect 141804 57934 141832 60044
rect 141792 57928 141844 57934
rect 141792 57870 141844 57876
rect 141608 57520 141660 57526
rect 141608 57462 141660 57468
rect 141516 56636 141568 56642
rect 141516 56578 141568 56584
rect 141620 51074 141648 57462
rect 141884 56772 141936 56778
rect 141884 56714 141936 56720
rect 141896 52834 141924 56714
rect 142068 56636 142120 56642
rect 142068 56578 142120 56584
rect 141884 52828 141936 52834
rect 141884 52770 141936 52776
rect 141528 51046 141648 51074
rect 141528 14482 141556 51046
rect 141516 14476 141568 14482
rect 141516 14418 141568 14424
rect 142080 12102 142108 56578
rect 142172 55214 142200 60044
rect 142448 56642 142476 60044
rect 142528 57792 142580 57798
rect 142528 57734 142580 57740
rect 142540 57526 142568 57734
rect 142724 57662 142752 60044
rect 142712 57656 142764 57662
rect 142712 57598 142764 57604
rect 142528 57520 142580 57526
rect 142528 57462 142580 57468
rect 142436 56636 142488 56642
rect 142436 56578 142488 56584
rect 142160 55208 142212 55214
rect 142160 55150 142212 55156
rect 143092 55146 143120 60044
rect 143172 56636 143224 56642
rect 143172 56578 143224 56584
rect 143080 55140 143132 55146
rect 143080 55082 143132 55088
rect 142068 12096 142120 12102
rect 142068 12038 142120 12044
rect 143184 12034 143212 56578
rect 143172 12028 143224 12034
rect 143172 11970 143224 11976
rect 143368 11966 143396 60044
rect 143644 57458 143672 60044
rect 143632 57452 143684 57458
rect 143632 57394 143684 57400
rect 143540 57112 143592 57118
rect 143540 57054 143592 57060
rect 143552 55418 143580 57054
rect 143632 56840 143684 56846
rect 143632 56782 143684 56788
rect 143540 55412 143592 55418
rect 143540 55354 143592 55360
rect 143644 54330 143672 56782
rect 143920 55078 143948 60044
rect 144184 56976 144236 56982
rect 144184 56918 144236 56924
rect 143908 55072 143960 55078
rect 143908 55014 143960 55020
rect 143632 54324 143684 54330
rect 143632 54266 143684 54272
rect 144196 17066 144224 56918
rect 144288 56642 144316 60044
rect 144276 56636 144328 56642
rect 144276 56578 144328 56584
rect 144184 17060 144236 17066
rect 144184 17002 144236 17008
rect 143356 11960 143408 11966
rect 143356 11902 143408 11908
rect 143540 4480 143592 4486
rect 143540 4422 143592 4428
rect 141424 4412 141476 4418
rect 141424 4354 141476 4360
rect 142436 3596 142488 3602
rect 142436 3538 142488 3544
rect 142448 480 142476 3538
rect 143552 480 143580 4422
rect 144564 4078 144592 60044
rect 144644 56636 144696 56642
rect 144644 56578 144696 56584
rect 144656 11898 144684 56578
rect 144840 51074 144868 60044
rect 145116 56778 145144 60044
rect 145484 56846 145512 60044
rect 145472 56840 145524 56846
rect 145472 56782 145524 56788
rect 145104 56772 145156 56778
rect 145104 56714 145156 56720
rect 145760 56642 145788 60044
rect 145748 56636 145800 56642
rect 145748 56578 145800 56584
rect 146036 52358 146064 60044
rect 146312 57118 146340 60044
rect 146392 57180 146444 57186
rect 146392 57122 146444 57128
rect 146300 57112 146352 57118
rect 146300 57054 146352 57060
rect 146116 56908 146168 56914
rect 146116 56850 146168 56856
rect 146024 52352 146076 52358
rect 146024 52294 146076 52300
rect 144748 51046 144868 51074
rect 146128 51066 146156 56850
rect 146208 56636 146260 56642
rect 146208 56578 146260 56584
rect 146116 51060 146168 51066
rect 144748 16574 144776 51046
rect 146116 51002 146168 51008
rect 144748 16546 144868 16574
rect 144644 11892 144696 11898
rect 144644 11834 144696 11840
rect 144736 7812 144788 7818
rect 144736 7754 144788 7760
rect 144552 4072 144604 4078
rect 144552 4014 144604 4020
rect 144748 480 144776 7754
rect 144840 7070 144868 16546
rect 146220 7138 146248 56578
rect 146404 55486 146432 57122
rect 146680 56710 146708 60044
rect 146852 57520 146904 57526
rect 146852 57462 146904 57468
rect 146668 56704 146720 56710
rect 146668 56646 146720 56652
rect 146392 55480 146444 55486
rect 146392 55422 146444 55428
rect 146864 51074 146892 57462
rect 146956 52290 146984 60044
rect 147232 56642 147260 60044
rect 147404 56704 147456 56710
rect 147404 56646 147456 56652
rect 147220 56636 147272 56642
rect 147220 56578 147272 56584
rect 146944 52284 146996 52290
rect 146944 52226 146996 52232
rect 146864 51046 146984 51074
rect 146956 17950 146984 51046
rect 146944 17944 146996 17950
rect 146944 17886 146996 17892
rect 147416 7206 147444 56646
rect 147508 7274 147536 60044
rect 147772 57384 147824 57390
rect 147772 57326 147824 57332
rect 147680 56772 147732 56778
rect 147680 56714 147732 56720
rect 147588 56636 147640 56642
rect 147588 56578 147640 56584
rect 147496 7268 147548 7274
rect 147496 7210 147548 7216
rect 147404 7200 147456 7206
rect 147404 7142 147456 7148
rect 146208 7132 146260 7138
rect 146208 7074 146260 7080
rect 144828 7064 144880 7070
rect 144828 7006 144880 7012
rect 147128 4548 147180 4554
rect 147128 4490 147180 4496
rect 145932 3528 145984 3534
rect 145932 3470 145984 3476
rect 145944 480 145972 3470
rect 147140 480 147168 4490
rect 147600 3942 147628 56578
rect 147692 52426 147720 56714
rect 147680 52420 147732 52426
rect 147680 52362 147732 52368
rect 147784 16574 147812 57326
rect 147876 52222 147904 60044
rect 148152 57390 148180 60044
rect 148428 57594 148456 60044
rect 148704 57662 148732 60044
rect 148692 57656 148744 57662
rect 148692 57598 148744 57604
rect 148416 57588 148468 57594
rect 148416 57530 148468 57536
rect 148324 57520 148376 57526
rect 148324 57462 148376 57468
rect 148140 57384 148192 57390
rect 148140 57326 148192 57332
rect 147864 52216 147916 52222
rect 147864 52158 147916 52164
rect 148336 17270 148364 57462
rect 149072 56778 149100 60044
rect 149348 59004 149376 60044
rect 149164 58976 149376 59004
rect 149428 59016 149480 59022
rect 149164 56982 149192 58976
rect 149428 58958 149480 58964
rect 149440 57974 149468 58958
rect 149348 57946 149468 57974
rect 149152 56976 149204 56982
rect 149152 56918 149204 56924
rect 149060 56772 149112 56778
rect 149060 56714 149112 56720
rect 149348 56642 149376 57946
rect 149624 57526 149652 60044
rect 149612 57520 149664 57526
rect 149612 57462 149664 57468
rect 149900 56710 149928 60044
rect 150268 59022 150296 60044
rect 150256 59016 150308 59022
rect 150544 59004 150572 60044
rect 150624 59084 150676 59090
rect 150624 59026 150676 59032
rect 150256 58958 150308 58964
rect 150452 58976 150572 59004
rect 150164 56976 150216 56982
rect 150164 56918 150216 56924
rect 149888 56704 149940 56710
rect 149888 56646 149940 56652
rect 149336 56636 149388 56642
rect 149336 56578 149388 56584
rect 150072 56636 150124 56642
rect 150072 56578 150124 56584
rect 148324 17264 148376 17270
rect 148324 17206 148376 17212
rect 147784 16546 148364 16574
rect 147588 3936 147640 3942
rect 147588 3878 147640 3884
rect 148336 480 148364 16546
rect 150084 7410 150112 56578
rect 150072 7404 150124 7410
rect 150072 7346 150124 7352
rect 150176 7342 150204 56918
rect 150256 56772 150308 56778
rect 150256 56714 150308 56720
rect 150164 7336 150216 7342
rect 150164 7278 150216 7284
rect 149518 4040 149574 4049
rect 149518 3975 149574 3984
rect 149532 480 149560 3975
rect 150268 3874 150296 56714
rect 150348 56704 150400 56710
rect 150348 56646 150400 56652
rect 150256 3868 150308 3874
rect 150256 3810 150308 3816
rect 150360 3806 150388 56646
rect 150452 52154 150480 58976
rect 150636 57974 150664 59026
rect 150716 59016 150768 59022
rect 150716 58958 150768 58964
rect 150544 57946 150664 57974
rect 150440 52148 150492 52154
rect 150440 52090 150492 52096
rect 150544 52086 150572 57946
rect 150728 56710 150756 58958
rect 150820 56846 150848 60044
rect 150808 56840 150860 56846
rect 150808 56782 150860 56788
rect 150716 56704 150768 56710
rect 150716 56646 150768 56652
rect 151096 56642 151124 60044
rect 151464 59090 151492 60044
rect 151452 59084 151504 59090
rect 151452 59026 151504 59032
rect 151740 59022 151768 60044
rect 151728 59016 151780 59022
rect 151728 58958 151780 58964
rect 152016 57186 152044 60044
rect 152004 57180 152056 57186
rect 152004 57122 152056 57128
rect 151636 56840 151688 56846
rect 151636 56782 151688 56788
rect 151360 56704 151412 56710
rect 151360 56646 151412 56652
rect 151084 56636 151136 56642
rect 151084 56578 151136 56584
rect 150532 52080 150584 52086
rect 150532 52022 150584 52028
rect 151372 6769 151400 56646
rect 151544 56636 151596 56642
rect 151544 56578 151596 56584
rect 151556 7478 151584 56578
rect 151544 7472 151596 7478
rect 151544 7414 151596 7420
rect 151648 6905 151676 56782
rect 152292 52018 152320 60044
rect 152660 57390 152688 60044
rect 152556 57384 152608 57390
rect 152556 57326 152608 57332
rect 152648 57384 152700 57390
rect 152648 57326 152700 57332
rect 152568 57050 152596 57326
rect 152556 57044 152608 57050
rect 152556 56986 152608 56992
rect 152280 52012 152332 52018
rect 152280 51954 152332 51960
rect 152936 8294 152964 60044
rect 153108 57384 153160 57390
rect 153108 57326 153160 57332
rect 153016 57180 153068 57186
rect 153016 57122 153068 57128
rect 152924 8288 152976 8294
rect 152924 8230 152976 8236
rect 151820 7744 151872 7750
rect 151820 7686 151872 7692
rect 151634 6896 151690 6905
rect 151634 6831 151690 6840
rect 151358 6760 151414 6769
rect 151358 6695 151414 6704
rect 150348 3800 150400 3806
rect 150348 3742 150400 3748
rect 150622 3224 150678 3233
rect 150622 3159 150678 3168
rect 150636 480 150664 3159
rect 151832 480 151860 7686
rect 153028 7546 153056 57122
rect 153016 7540 153068 7546
rect 153016 7482 153068 7488
rect 153120 6633 153148 57326
rect 153212 53786 153240 60044
rect 153488 57186 153516 60044
rect 153856 57390 153884 60044
rect 153844 57384 153896 57390
rect 153844 57326 153896 57332
rect 153476 57180 153528 57186
rect 153476 57122 153528 57128
rect 154132 56778 154160 60044
rect 154304 57384 154356 57390
rect 154304 57326 154356 57332
rect 154212 57180 154264 57186
rect 154212 57122 154264 57128
rect 154120 56772 154172 56778
rect 154120 56714 154172 56720
rect 153200 53780 153252 53786
rect 153200 53722 153252 53728
rect 154224 6914 154252 57122
rect 154316 8226 154344 57326
rect 154304 8220 154356 8226
rect 154304 8162 154356 8168
rect 154224 6886 154344 6914
rect 153106 6624 153162 6633
rect 153106 6559 153162 6568
rect 154212 4616 154264 4622
rect 154212 4558 154264 4564
rect 153014 3904 153070 3913
rect 153014 3839 153070 3848
rect 153028 480 153056 3839
rect 154224 480 154252 4558
rect 154316 2174 154344 6886
rect 154304 2168 154356 2174
rect 154304 2110 154356 2116
rect 154408 2106 154436 60044
rect 154776 57186 154804 60044
rect 155052 57390 155080 60044
rect 155040 57384 155092 57390
rect 155040 57326 155092 57332
rect 154764 57180 154816 57186
rect 154764 57122 154816 57128
rect 155132 57112 155184 57118
rect 155132 57054 155184 57060
rect 155144 49026 155172 57054
rect 155328 56982 155356 60044
rect 155604 57610 155632 60044
rect 155604 57582 155816 57610
rect 155684 57384 155736 57390
rect 155684 57326 155736 57332
rect 155316 56976 155368 56982
rect 155316 56918 155368 56924
rect 155132 49020 155184 49026
rect 155132 48962 155184 48968
rect 155696 12578 155724 57326
rect 155684 12572 155736 12578
rect 155684 12514 155736 12520
rect 155788 8090 155816 57582
rect 155972 57186 156000 60044
rect 155868 57180 155920 57186
rect 155868 57122 155920 57128
rect 155960 57180 156012 57186
rect 155960 57122 156012 57128
rect 155880 8158 155908 57122
rect 156248 57118 156276 60044
rect 156524 57390 156552 60044
rect 156800 57610 156828 60044
rect 156800 57582 157012 57610
rect 156512 57384 156564 57390
rect 156512 57326 156564 57332
rect 156880 57180 156932 57186
rect 156880 57122 156932 57128
rect 156236 57112 156288 57118
rect 156236 57054 156288 57060
rect 156892 12646 156920 57122
rect 156984 12714 157012 57582
rect 157064 57384 157116 57390
rect 157064 57326 157116 57332
rect 156972 12708 157024 12714
rect 156972 12650 157024 12656
rect 156880 12640 156932 12646
rect 156880 12582 156932 12588
rect 155868 8152 155920 8158
rect 155868 8094 155920 8100
rect 155776 8084 155828 8090
rect 155776 8026 155828 8032
rect 157076 8022 157104 57326
rect 157064 8016 157116 8022
rect 157064 7958 157116 7964
rect 155408 7676 155460 7682
rect 155408 7618 155460 7624
rect 154396 2100 154448 2106
rect 154396 2042 154448 2048
rect 155420 480 155448 7618
rect 157168 6361 157196 60044
rect 157340 57180 157392 57186
rect 157340 57122 157392 57128
rect 157248 57112 157300 57118
rect 157248 57054 157300 57060
rect 157260 6497 157288 57054
rect 157352 56778 157380 57122
rect 157444 56778 157472 60044
rect 157340 56772 157392 56778
rect 157340 56714 157392 56720
rect 157432 56772 157484 56778
rect 157432 56714 157484 56720
rect 157720 56642 157748 60044
rect 157996 56710 158024 60044
rect 158364 56794 158392 60044
rect 158640 56930 158668 60044
rect 158640 56902 158760 56930
rect 158916 56914 158944 60044
rect 158364 56766 158668 56794
rect 157984 56704 158036 56710
rect 157984 56646 158036 56652
rect 158444 56704 158496 56710
rect 158444 56646 158496 56652
rect 158536 56704 158588 56710
rect 158536 56646 158588 56652
rect 157708 56636 157760 56642
rect 157708 56578 157760 56584
rect 158260 56636 158312 56642
rect 158260 56578 158312 56584
rect 158352 56636 158404 56642
rect 158352 56578 158404 56584
rect 158272 12782 158300 56578
rect 158364 12850 158392 56578
rect 158352 12844 158404 12850
rect 158352 12786 158404 12792
rect 158260 12776 158312 12782
rect 158260 12718 158312 12724
rect 158456 8362 158484 56646
rect 158444 8356 158496 8362
rect 158444 8298 158496 8304
rect 158548 7954 158576 56646
rect 158536 7948 158588 7954
rect 158536 7890 158588 7896
rect 158640 7886 158668 56766
rect 158732 56642 158760 56902
rect 158812 56908 158864 56914
rect 158812 56850 158864 56856
rect 158904 56908 158956 56914
rect 158904 56850 158956 56856
rect 158720 56636 158772 56642
rect 158720 56578 158772 56584
rect 158824 51074 158852 56850
rect 159192 56642 159220 60044
rect 159364 57044 159416 57050
rect 159364 56986 159416 56992
rect 159180 56636 159232 56642
rect 159180 56578 159232 56584
rect 158732 51046 158852 51074
rect 158732 49162 158760 51046
rect 158720 49156 158772 49162
rect 158720 49098 158772 49104
rect 159376 19990 159404 56986
rect 159560 51074 159588 60044
rect 159732 56636 159784 56642
rect 159732 56578 159784 56584
rect 159744 55434 159772 56578
rect 159836 55570 159864 60044
rect 159836 55542 160048 55570
rect 159744 55406 159956 55434
rect 159560 51046 159864 51074
rect 159364 19984 159416 19990
rect 159364 19926 159416 19932
rect 159836 12918 159864 51046
rect 159824 12912 159876 12918
rect 159824 12854 159876 12860
rect 158628 7880 158680 7886
rect 158628 7822 158680 7828
rect 159928 7818 159956 55406
rect 159916 7812 159968 7818
rect 159916 7754 159968 7760
rect 158904 7608 158956 7614
rect 158904 7550 158956 7556
rect 157246 6488 157302 6497
rect 157246 6423 157302 6432
rect 157154 6352 157210 6361
rect 157154 6287 157210 6296
rect 157800 4684 157852 4690
rect 157800 4626 157852 4632
rect 156604 3460 156656 3466
rect 156604 3402 156656 3408
rect 156616 480 156644 3402
rect 157812 480 157840 4626
rect 158916 480 158944 7550
rect 160020 3738 160048 55542
rect 160112 54534 160140 60044
rect 160388 56642 160416 60044
rect 160756 56710 160784 60044
rect 160744 56704 160796 56710
rect 160744 56646 160796 56652
rect 160376 56636 160428 56642
rect 160376 56578 160428 56584
rect 160928 56636 160980 56642
rect 160928 56578 160980 56584
rect 160940 55434 160968 56578
rect 161032 55570 161060 60044
rect 161032 55542 161244 55570
rect 160940 55406 161152 55434
rect 161020 54664 161072 54670
rect 161020 54606 161072 54612
rect 160100 54528 160152 54534
rect 160100 54470 160152 54476
rect 161032 13054 161060 54606
rect 161020 13048 161072 13054
rect 161020 12990 161072 12996
rect 161124 12986 161152 55406
rect 161112 12980 161164 12986
rect 161112 12922 161164 12928
rect 161216 7682 161244 55542
rect 161308 54670 161336 60044
rect 161388 56704 161440 56710
rect 161388 56646 161440 56652
rect 161296 54664 161348 54670
rect 161296 54606 161348 54612
rect 161296 54528 161348 54534
rect 161296 54470 161348 54476
rect 161308 7750 161336 54470
rect 161296 7744 161348 7750
rect 161296 7686 161348 7692
rect 161204 7676 161256 7682
rect 161204 7618 161256 7624
rect 161294 3768 161350 3777
rect 160008 3732 160060 3738
rect 161294 3703 161350 3712
rect 160008 3674 160060 3680
rect 160098 3632 160154 3641
rect 160098 3567 160154 3576
rect 160112 480 160140 3567
rect 161308 480 161336 3703
rect 161400 3670 161428 56646
rect 161584 56642 161612 60044
rect 161848 57724 161900 57730
rect 161848 57666 161900 57672
rect 161572 56636 161624 56642
rect 161572 56578 161624 56584
rect 161860 51074 161888 57666
rect 161952 55298 161980 60044
rect 162228 55434 162256 60044
rect 162504 55570 162532 60044
rect 162676 56636 162728 56642
rect 162676 56578 162728 56584
rect 162504 55542 162624 55570
rect 162228 55406 162532 55434
rect 161952 55270 162440 55298
rect 161860 51046 162164 51074
rect 162136 17406 162164 51046
rect 162124 17400 162176 17406
rect 162124 17342 162176 17348
rect 162412 7614 162440 55270
rect 162504 13802 162532 55406
rect 162492 13796 162544 13802
rect 162492 13738 162544 13744
rect 162596 8498 162624 55542
rect 162584 8492 162636 8498
rect 162584 8434 162636 8440
rect 162688 8430 162716 56578
rect 162780 55010 162808 60044
rect 163148 56642 163176 60044
rect 163424 56914 163452 60044
rect 163412 56908 163464 56914
rect 163412 56850 163464 56856
rect 163136 56636 163188 56642
rect 163136 56578 163188 56584
rect 163700 56574 163728 60044
rect 163872 56636 163924 56642
rect 163872 56578 163924 56584
rect 163688 56568 163740 56574
rect 163688 56510 163740 56516
rect 162768 55004 162820 55010
rect 162768 54946 162820 54952
rect 163884 51074 163912 56578
rect 163976 55570 164004 60044
rect 164344 56710 164372 60044
rect 164332 56704 164384 56710
rect 164332 56646 164384 56652
rect 163976 55542 164096 55570
rect 163884 51046 164004 51074
rect 163976 13734 164004 51046
rect 163964 13728 164016 13734
rect 163964 13670 164016 13676
rect 164068 13666 164096 55542
rect 164620 54942 164648 60044
rect 164896 56642 164924 60044
rect 165068 56704 165120 56710
rect 165068 56646 165120 56652
rect 164884 56636 164936 56642
rect 164884 56578 164936 56584
rect 164608 54936 164660 54942
rect 164608 54878 164660 54884
rect 165080 51074 165108 56646
rect 165172 55570 165200 60044
rect 165344 56636 165396 56642
rect 165344 56578 165396 56584
rect 165172 55542 165292 55570
rect 165080 51046 165200 51074
rect 164056 13660 164108 13666
rect 164056 13602 164108 13608
rect 163688 9444 163740 9450
rect 163688 9386 163740 9392
rect 162676 8424 162728 8430
rect 162676 8366 162728 8372
rect 162400 7608 162452 7614
rect 162400 7550 162452 7556
rect 162492 4752 162544 4758
rect 162492 4694 162544 4700
rect 161388 3664 161440 3670
rect 161388 3606 161440 3612
rect 162504 480 162532 4694
rect 163700 480 163728 9386
rect 165172 6225 165200 51046
rect 165158 6216 165214 6225
rect 165158 6151 165214 6160
rect 165264 3602 165292 55542
rect 165356 13598 165384 56578
rect 165540 54874 165568 60044
rect 165712 57452 165764 57458
rect 165712 57394 165764 57400
rect 165528 54868 165580 54874
rect 165528 54810 165580 54816
rect 165724 49094 165752 57394
rect 165816 56710 165844 60044
rect 165804 56704 165856 56710
rect 165804 56646 165856 56652
rect 166092 56642 166120 60044
rect 166080 56636 166132 56642
rect 166080 56578 166132 56584
rect 166460 54806 166488 60044
rect 166632 56636 166684 56642
rect 166632 56578 166684 56584
rect 166448 54800 166500 54806
rect 166448 54742 166500 54748
rect 165712 49088 165764 49094
rect 165712 49030 165764 49036
rect 165344 13592 165396 13598
rect 165344 13534 165396 13540
rect 166644 8566 166672 56578
rect 166736 13462 166764 60044
rect 167012 57322 167040 60044
rect 167184 57452 167236 57458
rect 167184 57394 167236 57400
rect 167000 57316 167052 57322
rect 167000 57258 167052 57264
rect 166816 56704 166868 56710
rect 166816 56646 166868 56652
rect 166828 13530 166856 56646
rect 167196 54738 167224 57394
rect 167288 56506 167316 60044
rect 167656 57730 167684 60044
rect 167644 57724 167696 57730
rect 167644 57666 167696 57672
rect 167276 56500 167328 56506
rect 167276 56442 167328 56448
rect 167932 55214 167960 60044
rect 168104 57724 168156 57730
rect 168104 57666 168156 57672
rect 167932 55186 168052 55214
rect 167184 54732 167236 54738
rect 167184 54674 167236 54680
rect 166816 13524 166868 13530
rect 166816 13466 166868 13472
rect 166724 13456 166776 13462
rect 166724 13398 166776 13404
rect 167184 9376 167236 9382
rect 167184 9318 167236 9324
rect 166632 8560 166684 8566
rect 166632 8502 166684 8508
rect 166080 5500 166132 5506
rect 166080 5442 166132 5448
rect 165252 3596 165304 3602
rect 165252 3538 165304 3544
rect 164882 3496 164938 3505
rect 164882 3431 164938 3440
rect 164896 480 164924 3431
rect 166092 480 166120 5442
rect 167196 480 167224 9318
rect 168024 3534 168052 55186
rect 168116 13394 168144 57666
rect 168208 57458 168236 60044
rect 168196 57452 168248 57458
rect 168196 57394 168248 57400
rect 168484 57390 168512 60044
rect 168852 57458 168880 60044
rect 168840 57452 168892 57458
rect 168840 57394 168892 57400
rect 168472 57384 168524 57390
rect 168472 57326 168524 57332
rect 168196 57316 168248 57322
rect 168196 57258 168248 57264
rect 168748 57316 168800 57322
rect 168748 57258 168800 57264
rect 168104 13388 168156 13394
rect 168104 13330 168156 13336
rect 168208 8634 168236 57258
rect 168196 8628 168248 8634
rect 168196 8570 168248 8576
rect 168760 6914 168788 57258
rect 169128 53718 169156 60044
rect 169300 57724 169352 57730
rect 169300 57666 169352 57672
rect 169116 53712 169168 53718
rect 169116 53654 169168 53660
rect 168392 6886 168788 6914
rect 168012 3528 168064 3534
rect 168012 3470 168064 3476
rect 168392 480 168420 6886
rect 169312 3233 169340 57666
rect 169404 13258 169432 60044
rect 169680 57730 169708 60044
rect 169668 57724 169720 57730
rect 169668 57666 169720 57672
rect 169576 57452 169628 57458
rect 169576 57394 169628 57400
rect 169484 57384 169536 57390
rect 169484 57326 169536 57332
rect 169496 13326 169524 57326
rect 169588 16574 169616 57394
rect 170048 53650 170076 60044
rect 170324 56982 170352 60044
rect 170312 56976 170364 56982
rect 170312 56918 170364 56924
rect 170600 55214 170628 60044
rect 170876 57168 170904 60044
rect 171244 57730 171272 60044
rect 171232 57724 171284 57730
rect 171232 57666 171284 57672
rect 170876 57140 170996 57168
rect 170864 56976 170916 56982
rect 170864 56918 170916 56924
rect 170600 55186 170812 55214
rect 170036 53644 170088 53650
rect 170036 53586 170088 53592
rect 169588 16546 169708 16574
rect 169484 13320 169536 13326
rect 169484 13262 169536 13268
rect 169392 13252 169444 13258
rect 169392 13194 169444 13200
rect 169576 5432 169628 5438
rect 169576 5374 169628 5380
rect 169298 3224 169354 3233
rect 169298 3159 169354 3168
rect 169588 480 169616 5374
rect 169680 3466 169708 16546
rect 170680 9308 170732 9314
rect 170680 9250 170732 9256
rect 169668 3460 169720 3466
rect 169668 3402 169720 3408
rect 170692 1714 170720 9250
rect 170784 4049 170812 55186
rect 170876 13190 170904 56918
rect 170864 13184 170916 13190
rect 170864 13126 170916 13132
rect 170968 8702 170996 57140
rect 171520 56778 171548 60044
rect 171600 57248 171652 57254
rect 171600 57190 171652 57196
rect 171508 56772 171560 56778
rect 171508 56714 171560 56720
rect 171612 16574 171640 57190
rect 171796 45554 171824 60044
rect 172072 54670 172100 60044
rect 172244 57724 172296 57730
rect 172244 57666 172296 57672
rect 172060 54664 172112 54670
rect 172060 54606 172112 54612
rect 171796 45526 172192 45554
rect 171612 16546 172008 16574
rect 170956 8696 171008 8702
rect 170956 8638 171008 8644
rect 170770 4040 170826 4049
rect 170770 3975 170826 3984
rect 170692 1686 170812 1714
rect 170784 480 170812 1686
rect 171980 480 172008 16546
rect 172164 8770 172192 45526
rect 172256 13122 172284 57666
rect 172440 45554 172468 60044
rect 172716 57730 172744 60044
rect 172704 57724 172756 57730
rect 172704 57666 172756 57672
rect 172992 51950 173020 60044
rect 173268 56642 173296 60044
rect 173256 56636 173308 56642
rect 173256 56578 173308 56584
rect 173636 55214 173664 60044
rect 173808 57724 173860 57730
rect 173808 57666 173860 57672
rect 173636 55186 173756 55214
rect 172980 51944 173032 51950
rect 172980 51886 173032 51892
rect 172348 45526 172468 45554
rect 172244 13116 172296 13122
rect 172244 13058 172296 13064
rect 172348 8906 172376 45526
rect 173728 9654 173756 55186
rect 173716 9648 173768 9654
rect 173716 9590 173768 9596
rect 172336 8900 172388 8906
rect 172336 8842 172388 8848
rect 173820 8838 173848 57666
rect 173912 51882 173940 60044
rect 174188 57458 174216 60044
rect 174464 57730 174492 60044
rect 174452 57724 174504 57730
rect 174452 57666 174504 57672
rect 174176 57452 174228 57458
rect 174176 57394 174228 57400
rect 173900 51876 173952 51882
rect 173900 51818 173952 51824
rect 174832 50998 174860 60044
rect 175108 57610 175136 60044
rect 175188 57724 175240 57730
rect 175188 57666 175240 57672
rect 175016 57582 175136 57610
rect 175016 56914 175044 57582
rect 175096 57452 175148 57458
rect 175096 57394 175148 57400
rect 175004 56908 175056 56914
rect 175004 56850 175056 56856
rect 174820 50992 174872 50998
rect 174820 50934 174872 50940
rect 175108 11830 175136 57394
rect 175096 11824 175148 11830
rect 175096 11766 175148 11772
rect 175200 9586 175228 57666
rect 175384 57458 175412 60044
rect 175556 57724 175608 57730
rect 175556 57666 175608 57672
rect 175372 57452 175424 57458
rect 175372 57394 175424 57400
rect 175568 51814 175596 57666
rect 175660 53514 175688 60044
rect 176028 55214 176056 60044
rect 176304 55214 176332 60044
rect 176580 57730 176608 60044
rect 176568 57724 176620 57730
rect 176568 57666 176620 57672
rect 176476 57452 176528 57458
rect 176476 57394 176528 57400
rect 176028 55186 176240 55214
rect 176304 55186 176424 55214
rect 175648 53508 175700 53514
rect 175648 53450 175700 53456
rect 175556 51808 175608 51814
rect 175556 51750 175608 51756
rect 175188 9580 175240 9586
rect 175188 9522 175240 9528
rect 174268 9240 174320 9246
rect 174268 9182 174320 9188
rect 173808 8832 173860 8838
rect 173808 8774 173860 8780
rect 172152 8764 172204 8770
rect 172152 8706 172204 8712
rect 173164 5364 173216 5370
rect 173164 5306 173216 5312
rect 173176 480 173204 5306
rect 174280 480 174308 9182
rect 176212 3913 176240 55186
rect 176396 9450 176424 55186
rect 176488 9518 176516 57394
rect 176856 57254 176884 60044
rect 177224 57730 177252 60044
rect 177212 57724 177264 57730
rect 177212 57666 177264 57672
rect 176844 57248 176896 57254
rect 176844 57190 176896 57196
rect 177304 56840 177356 56846
rect 177304 56782 177356 56788
rect 177316 17474 177344 56782
rect 177500 50930 177528 60044
rect 177776 55214 177804 60044
rect 177948 57724 178000 57730
rect 177948 57666 178000 57672
rect 178040 57724 178092 57730
rect 178040 57666 178092 57672
rect 177776 55186 177896 55214
rect 177488 50924 177540 50930
rect 177488 50866 177540 50872
rect 177304 17468 177356 17474
rect 177304 17410 177356 17416
rect 177868 11762 177896 55186
rect 177856 11756 177908 11762
rect 177856 11698 177908 11704
rect 176476 9512 176528 9518
rect 176476 9454 176528 9460
rect 176384 9444 176436 9450
rect 176384 9386 176436 9392
rect 177960 9382 177988 57666
rect 178052 50794 178080 57666
rect 178144 57458 178172 60044
rect 178132 57452 178184 57458
rect 178132 57394 178184 57400
rect 178420 50862 178448 60044
rect 178696 57390 178724 60044
rect 178972 57610 179000 60044
rect 179340 57730 179368 60044
rect 179328 57724 179380 57730
rect 179328 57666 179380 57672
rect 178972 57582 179368 57610
rect 179236 57452 179288 57458
rect 179236 57394 179288 57400
rect 178684 57384 178736 57390
rect 178684 57326 178736 57332
rect 178408 50856 178460 50862
rect 178408 50798 178460 50804
rect 178040 50788 178092 50794
rect 178040 50730 178092 50736
rect 177948 9376 178000 9382
rect 177948 9318 178000 9324
rect 179248 9314 179276 57394
rect 179236 9308 179288 9314
rect 179236 9250 179288 9256
rect 179340 9246 179368 57582
rect 179616 57322 179644 60044
rect 179604 57316 179656 57322
rect 179604 57258 179656 57264
rect 179892 56778 179920 60044
rect 179880 56772 179932 56778
rect 179880 56714 179932 56720
rect 180168 55214 180196 60044
rect 180536 57610 180564 60044
rect 180812 58154 180840 60044
rect 180812 58126 180932 58154
rect 180800 58064 180852 58070
rect 180800 58006 180852 58012
rect 180708 57996 180760 58002
rect 180812 57974 180840 58006
rect 180760 57946 180840 57974
rect 180708 57938 180760 57944
rect 180708 57724 180760 57730
rect 180708 57666 180760 57672
rect 180352 57582 180564 57610
rect 180352 57390 180380 57582
rect 180720 57474 180748 57666
rect 180444 57446 180748 57474
rect 180340 57384 180392 57390
rect 180340 57326 180392 57332
rect 180444 57254 180472 57446
rect 180708 57316 180760 57322
rect 180708 57258 180760 57264
rect 180800 57316 180852 57322
rect 180800 57258 180852 57264
rect 180432 57248 180484 57254
rect 180432 57190 180484 57196
rect 180522 57216 180578 57225
rect 180522 57151 180578 57160
rect 180536 56914 180564 57151
rect 180524 56908 180576 56914
rect 180524 56850 180576 56856
rect 180524 56772 180576 56778
rect 180524 56714 180576 56720
rect 180536 56658 180564 56714
rect 180536 56630 180656 56658
rect 180168 55186 180564 55214
rect 180536 13938 180564 55186
rect 180524 13932 180576 13938
rect 180524 13874 180576 13880
rect 179328 9240 179380 9246
rect 179328 9182 179380 9188
rect 180628 9178 180656 56630
rect 177856 9172 177908 9178
rect 177856 9114 177908 9120
rect 180616 9172 180668 9178
rect 180616 9114 180668 9120
rect 176660 5296 176712 5302
rect 176660 5238 176712 5244
rect 176198 3904 176254 3913
rect 176198 3839 176254 3848
rect 175462 3360 175518 3369
rect 175462 3295 175518 3304
rect 175476 480 175504 3295
rect 176672 480 176700 5238
rect 177868 480 177896 9114
rect 180248 5228 180300 5234
rect 180248 5170 180300 5176
rect 179052 3120 179104 3126
rect 179052 3062 179104 3068
rect 179064 480 179092 3062
rect 180260 480 180288 5170
rect 180720 3777 180748 57258
rect 180812 57225 180840 57258
rect 180798 57216 180854 57225
rect 180798 57151 180854 57160
rect 180904 56846 180932 58126
rect 181088 57730 181116 60044
rect 181168 58064 181220 58070
rect 181168 58006 181220 58012
rect 180984 57724 181036 57730
rect 180984 57666 181036 57672
rect 181076 57724 181128 57730
rect 181076 57666 181128 57672
rect 180892 56840 180944 56846
rect 180892 56782 180944 56788
rect 180996 56642 181024 57666
rect 181180 56710 181208 58006
rect 181364 57254 181392 60044
rect 181732 58002 181760 60044
rect 181720 57996 181772 58002
rect 181720 57938 181772 57944
rect 181720 57724 181772 57730
rect 181720 57666 181772 57672
rect 181352 57248 181404 57254
rect 181352 57190 181404 57196
rect 181168 56704 181220 56710
rect 181168 56646 181220 56652
rect 180984 56636 181036 56642
rect 180984 56578 181036 56584
rect 181732 14006 181760 57666
rect 182008 57610 182036 60044
rect 181824 57582 182036 57610
rect 181720 14000 181772 14006
rect 181720 13942 181772 13948
rect 181824 9489 181852 57582
rect 182284 57254 182312 60044
rect 182560 57730 182588 60044
rect 182548 57724 182600 57730
rect 182548 57666 182600 57672
rect 181996 57248 182048 57254
rect 181996 57190 182048 57196
rect 182272 57248 182324 57254
rect 182272 57190 182324 57196
rect 181904 56840 181956 56846
rect 181904 56782 181956 56788
rect 181810 9480 181866 9489
rect 181810 9415 181866 9424
rect 181916 9110 181944 56782
rect 181444 9104 181496 9110
rect 181444 9046 181496 9052
rect 181904 9104 181956 9110
rect 181904 9046 181956 9052
rect 180706 3768 180762 3777
rect 180706 3703 180762 3712
rect 181456 480 181484 9046
rect 182008 3641 182036 57190
rect 182928 56710 182956 60044
rect 183100 57724 183152 57730
rect 183100 57666 183152 57672
rect 182088 56704 182140 56710
rect 182088 56646 182140 56652
rect 182916 56704 182968 56710
rect 182916 56646 182968 56652
rect 181994 3632 182050 3641
rect 181994 3567 182050 3576
rect 182100 3505 182128 56646
rect 182548 14476 182600 14482
rect 182548 14418 182600 14424
rect 182086 3496 182142 3505
rect 182086 3431 182142 3440
rect 182560 480 182588 14418
rect 183112 3369 183140 57666
rect 183204 14142 183232 60044
rect 183284 57248 183336 57254
rect 183284 57190 183336 57196
rect 183192 14136 183244 14142
rect 183192 14078 183244 14084
rect 183296 14074 183324 57190
rect 183376 56704 183428 56710
rect 183376 56646 183428 56652
rect 183284 14068 183336 14074
rect 183284 14010 183336 14016
rect 183388 9353 183416 56646
rect 183480 56438 183508 60044
rect 183756 57730 183784 60044
rect 183744 57724 183796 57730
rect 183744 57666 183796 57672
rect 183560 57316 183612 57322
rect 183560 57258 183612 57264
rect 183572 56710 183600 57258
rect 184124 56846 184152 60044
rect 184112 56840 184164 56846
rect 184112 56782 184164 56788
rect 183560 56704 183612 56710
rect 183560 56646 183612 56652
rect 183468 56432 183520 56438
rect 183468 56374 183520 56380
rect 184400 56302 184428 60044
rect 184676 57304 184704 60044
rect 184756 57724 184808 57730
rect 184756 57666 184808 57672
rect 184584 57276 184704 57304
rect 184388 56296 184440 56302
rect 184388 56238 184440 56244
rect 183374 9344 183430 9353
rect 183374 9279 183430 9288
rect 184584 9081 184612 57276
rect 184664 56840 184716 56846
rect 184664 56782 184716 56788
rect 184676 14210 184704 56782
rect 184664 14204 184716 14210
rect 184664 14146 184716 14152
rect 184768 9217 184796 57666
rect 184952 56846 184980 60044
rect 184940 56840 184992 56846
rect 184940 56782 184992 56788
rect 185320 56370 185348 60044
rect 185308 56364 185360 56370
rect 185308 56306 185360 56312
rect 185596 55214 185624 60044
rect 185872 57610 185900 60044
rect 186148 58154 186176 60044
rect 186148 58126 186268 58154
rect 185872 57582 186176 57610
rect 186044 56840 186096 56846
rect 186044 56782 186096 56788
rect 185596 55186 185992 55214
rect 184754 9208 184810 9217
rect 184754 9143 184810 9152
rect 184570 9072 184626 9081
rect 185964 9042 185992 55186
rect 186056 14278 186084 56782
rect 186148 14346 186176 57582
rect 186240 56234 186268 58126
rect 186516 57458 186544 60044
rect 186792 57730 186820 60044
rect 186780 57724 186832 57730
rect 186780 57666 186832 57672
rect 186504 57452 186556 57458
rect 186504 57394 186556 57400
rect 186228 56228 186280 56234
rect 186228 56170 186280 56176
rect 187068 56030 187096 60044
rect 187056 56024 187108 56030
rect 187056 55966 187108 55972
rect 186136 14340 186188 14346
rect 186136 14282 186188 14288
rect 186044 14272 186096 14278
rect 186044 14214 186096 14220
rect 187344 12730 187372 60044
rect 187712 57730 187740 60044
rect 187424 57724 187476 57730
rect 187424 57666 187476 57672
rect 187700 57724 187752 57730
rect 187700 57666 187752 57672
rect 187436 14414 187464 57666
rect 187516 57452 187568 57458
rect 187516 57394 187568 57400
rect 187608 57452 187660 57458
rect 187608 57394 187660 57400
rect 187424 14408 187476 14414
rect 187424 14350 187476 14356
rect 187344 12702 187464 12730
rect 184570 9007 184626 9016
rect 184940 9036 184992 9042
rect 184940 8978 184992 8984
rect 185952 9036 186004 9042
rect 185952 8978 186004 8984
rect 183744 5160 183796 5166
rect 183744 5102 183796 5108
rect 183098 3360 183154 3369
rect 183098 3295 183154 3304
rect 183756 480 183784 5102
rect 184952 480 184980 8978
rect 187332 8968 187384 8974
rect 187436 8945 187464 12702
rect 187528 8974 187556 57394
rect 187620 56642 187648 57394
rect 187608 56636 187660 56642
rect 187608 56578 187660 56584
rect 187988 56166 188016 60044
rect 187976 56160 188028 56166
rect 187976 56102 188028 56108
rect 188264 53582 188292 60044
rect 188540 55214 188568 60044
rect 188908 57882 188936 60044
rect 188908 57854 189028 57882
rect 188896 57724 188948 57730
rect 188896 57666 188948 57672
rect 188540 55186 188752 55214
rect 188252 53576 188304 53582
rect 188252 53518 188304 53524
rect 188724 15094 188752 55186
rect 188908 15162 188936 57666
rect 189000 55962 189028 57854
rect 189080 57724 189132 57730
rect 189080 57666 189132 57672
rect 188988 55956 189040 55962
rect 188988 55898 189040 55904
rect 189092 54602 189120 57666
rect 189184 56098 189212 60044
rect 189460 56846 189488 60044
rect 189448 56840 189500 56846
rect 189448 56782 189500 56788
rect 189172 56092 189224 56098
rect 189172 56034 189224 56040
rect 189828 55214 189856 60044
rect 190104 57730 190132 60044
rect 190092 57724 190144 57730
rect 190092 57666 190144 57672
rect 190380 57610 190408 60044
rect 190656 57730 190684 60044
rect 190644 57724 190696 57730
rect 190644 57666 190696 57672
rect 190196 57582 190408 57610
rect 189828 55186 190132 55214
rect 189080 54596 189132 54602
rect 189080 54538 189132 54544
rect 188896 15156 188948 15162
rect 188896 15098 188948 15104
rect 188712 15088 188764 15094
rect 188712 15030 188764 15036
rect 188528 10940 188580 10946
rect 188528 10882 188580 10888
rect 187516 8968 187568 8974
rect 187332 8910 187384 8916
rect 187422 8936 187478 8945
rect 186136 4412 186188 4418
rect 186136 4354 186188 4360
rect 186148 480 186176 4354
rect 187344 480 187372 8910
rect 187516 8910 187568 8916
rect 187422 8871 187478 8880
rect 188540 480 188568 10882
rect 189724 5092 189776 5098
rect 189724 5034 189776 5040
rect 189736 480 189764 5034
rect 190104 4282 190132 55186
rect 190196 14958 190224 57582
rect 190368 57452 190420 57458
rect 190368 57394 190420 57400
rect 190276 56840 190328 56846
rect 190276 56782 190328 56788
rect 190288 15026 190316 56782
rect 190380 56710 190408 57394
rect 190368 56704 190420 56710
rect 190368 56646 190420 56652
rect 191024 53446 191052 60044
rect 191300 56846 191328 60044
rect 191576 57610 191604 60044
rect 191656 57724 191708 57730
rect 191656 57666 191708 57672
rect 191484 57582 191604 57610
rect 191288 56840 191340 56846
rect 191288 56782 191340 56788
rect 191012 53440 191064 53446
rect 191012 53382 191064 53388
rect 190276 15020 190328 15026
rect 190276 14962 190328 14968
rect 190184 14952 190236 14958
rect 190184 14894 190236 14900
rect 190828 10872 190880 10878
rect 190828 10814 190880 10820
rect 190092 4276 190144 4282
rect 190092 4218 190144 4224
rect 190840 480 190868 10814
rect 191484 4418 191512 57582
rect 191564 56840 191616 56846
rect 191564 56782 191616 56788
rect 191576 14890 191604 56782
rect 191564 14884 191616 14890
rect 191564 14826 191616 14832
rect 191472 4412 191524 4418
rect 191472 4354 191524 4360
rect 191668 4350 191696 57666
rect 191852 53174 191880 60044
rect 192024 57724 192076 57730
rect 192024 57666 192076 57672
rect 192036 53378 192064 57666
rect 192220 56846 192248 60044
rect 192208 56840 192260 56846
rect 192208 56782 192260 56788
rect 192496 55214 192524 60044
rect 192772 57730 192800 60044
rect 192760 57724 192812 57730
rect 192760 57666 192812 57672
rect 192944 56840 192996 56846
rect 192944 56782 192996 56788
rect 192496 55186 192800 55214
rect 192024 53372 192076 53378
rect 192024 53314 192076 53320
rect 191840 53168 191892 53174
rect 191840 53110 191892 53116
rect 192024 10804 192076 10810
rect 192024 10746 192076 10752
rect 191656 4344 191708 4350
rect 191656 4286 191708 4292
rect 192036 480 192064 10746
rect 192772 4486 192800 55186
rect 192956 14822 192984 56782
rect 192944 14816 192996 14822
rect 192944 14758 192996 14764
rect 193048 14754 193076 60044
rect 193416 56846 193444 60044
rect 193404 56840 193456 56846
rect 193404 56782 193456 56788
rect 193692 53310 193720 60044
rect 193968 57474 193996 60044
rect 194244 57610 194272 60044
rect 194244 57582 194456 57610
rect 193968 57446 194364 57474
rect 194232 56840 194284 56846
rect 194232 56782 194284 56788
rect 193680 53304 193732 53310
rect 193680 53246 193732 53252
rect 193036 14748 193088 14754
rect 193036 14690 193088 14696
rect 193220 10736 193272 10742
rect 193220 10678 193272 10684
rect 192760 4480 192812 4486
rect 192760 4422 192812 4428
rect 193232 3126 193260 10678
rect 194244 5030 194272 56782
rect 194336 14686 194364 57446
rect 194428 16574 194456 57582
rect 194612 53242 194640 60044
rect 194888 57730 194916 60044
rect 194876 57724 194928 57730
rect 194876 57666 194928 57672
rect 194600 53236 194652 53242
rect 194600 53178 194652 53184
rect 195164 45554 195192 60044
rect 195440 53106 195468 60044
rect 195704 57724 195756 57730
rect 195704 57666 195756 57672
rect 195428 53100 195480 53106
rect 195428 53042 195480 53048
rect 195164 45526 195560 45554
rect 194428 16546 194548 16574
rect 194324 14680 194376 14686
rect 194324 14622 194376 14628
rect 193312 5024 193364 5030
rect 193312 4966 193364 4972
rect 194232 5024 194284 5030
rect 194232 4966 194284 4972
rect 193220 3120 193272 3126
rect 193220 3062 193272 3068
rect 193324 2530 193352 4966
rect 194520 4554 194548 16546
rect 195428 10668 195480 10674
rect 195428 10610 195480 10616
rect 194508 4548 194560 4554
rect 194508 4490 194560 4496
rect 195440 3482 195468 10610
rect 195532 4622 195560 45526
rect 195716 14618 195744 57666
rect 195704 14612 195756 14618
rect 195704 14554 195756 14560
rect 195808 14550 195836 60044
rect 196084 56710 196112 60044
rect 196360 57730 196388 60044
rect 196348 57724 196400 57730
rect 196348 57666 196400 57672
rect 196072 56704 196124 56710
rect 196072 56646 196124 56652
rect 196636 55214 196664 60044
rect 197004 57882 197032 60044
rect 196912 57854 197032 57882
rect 196912 56846 196940 57854
rect 196992 57724 197044 57730
rect 196992 57666 197044 57672
rect 196900 56840 196952 56846
rect 196900 56782 196952 56788
rect 196636 55186 196940 55214
rect 195796 14544 195848 14550
rect 195796 14486 195848 14492
rect 196912 14482 196940 55186
rect 196900 14476 196952 14482
rect 196900 14418 196952 14424
rect 197004 10266 197032 57666
rect 197280 57610 197308 60044
rect 197096 57582 197308 57610
rect 197096 11014 197124 57582
rect 197268 56840 197320 56846
rect 197268 56782 197320 56788
rect 197176 56704 197228 56710
rect 197176 56646 197228 56652
rect 197084 11008 197136 11014
rect 197084 10950 197136 10956
rect 196992 10260 197044 10266
rect 196992 10202 197044 10208
rect 196808 4956 196860 4962
rect 196808 4898 196860 4904
rect 195520 4616 195572 4622
rect 195520 4558 195572 4564
rect 195440 3454 195652 3482
rect 194416 3120 194468 3126
rect 194416 3062 194468 3068
rect 193232 2502 193352 2530
rect 193232 480 193260 2502
rect 194428 480 194456 3062
rect 195624 480 195652 3454
rect 196820 480 196848 4898
rect 197188 4758 197216 56646
rect 197280 5506 197308 56782
rect 197556 50590 197584 60044
rect 197636 57724 197688 57730
rect 197636 57666 197688 57672
rect 197544 50584 197596 50590
rect 197544 50526 197596 50532
rect 197648 50454 197676 57666
rect 197832 56846 197860 60044
rect 197820 56840 197872 56846
rect 197820 56782 197872 56788
rect 198200 55214 198228 60044
rect 198476 57730 198504 60044
rect 198464 57724 198516 57730
rect 198464 57666 198516 57672
rect 198648 56840 198700 56846
rect 198648 56782 198700 56788
rect 198200 55186 198596 55214
rect 197636 50448 197688 50454
rect 197636 50390 197688 50396
rect 198568 10946 198596 55186
rect 198556 10940 198608 10946
rect 198556 10882 198608 10888
rect 197912 10600 197964 10606
rect 197912 10542 197964 10548
rect 197268 5500 197320 5506
rect 197268 5442 197320 5448
rect 197176 4752 197228 4758
rect 197176 4694 197228 4700
rect 197924 480 197952 10542
rect 198660 5438 198688 56782
rect 198752 56710 198780 60044
rect 199028 57730 199056 60044
rect 199016 57724 199068 57730
rect 199016 57666 199068 57672
rect 198740 56704 198792 56710
rect 198740 56646 198792 56652
rect 199396 51746 199424 60044
rect 199672 56846 199700 60044
rect 199752 57724 199804 57730
rect 199752 57666 199804 57672
rect 199660 56840 199712 56846
rect 199660 56782 199712 56788
rect 199660 56704 199712 56710
rect 199660 56646 199712 56652
rect 199384 51740 199436 51746
rect 199384 51682 199436 51688
rect 199108 10532 199160 10538
rect 199108 10474 199160 10480
rect 198648 5432 198700 5438
rect 198648 5374 198700 5380
rect 199120 480 199148 10474
rect 199672 5370 199700 56646
rect 199764 10878 199792 57666
rect 199948 57610 199976 60044
rect 199856 57582 199976 57610
rect 199752 10872 199804 10878
rect 199752 10814 199804 10820
rect 199856 10810 199884 57582
rect 199936 56840 199988 56846
rect 199936 56782 199988 56788
rect 199844 10804 199896 10810
rect 199844 10746 199896 10752
rect 199660 5364 199712 5370
rect 199660 5306 199712 5312
rect 199948 5302 199976 56782
rect 200224 50726 200252 60044
rect 200592 56914 200620 60044
rect 200868 57730 200896 60044
rect 200856 57724 200908 57730
rect 200856 57666 200908 57672
rect 200580 56908 200632 56914
rect 200580 56850 200632 56856
rect 200212 50720 200264 50726
rect 200212 50662 200264 50668
rect 201144 50658 201172 60044
rect 201316 57724 201368 57730
rect 201316 57666 201368 57672
rect 201132 50652 201184 50658
rect 201132 50594 201184 50600
rect 201328 10742 201356 57666
rect 201408 56908 201460 56914
rect 201408 56850 201460 56856
rect 201316 10736 201368 10742
rect 201316 10678 201368 10684
rect 199936 5296 199988 5302
rect 199936 5238 199988 5244
rect 201420 4894 201448 56850
rect 201512 56710 201540 60044
rect 201788 57730 201816 60044
rect 201776 57724 201828 57730
rect 201776 57666 201828 57672
rect 201500 56704 201552 56710
rect 201500 56646 201552 56652
rect 202064 50386 202092 60044
rect 202340 56914 202368 60044
rect 202512 57724 202564 57730
rect 202512 57666 202564 57672
rect 202328 56908 202380 56914
rect 202328 56850 202380 56856
rect 202420 56704 202472 56710
rect 202420 56646 202472 56652
rect 202052 50380 202104 50386
rect 202052 50322 202104 50328
rect 201592 10464 201644 10470
rect 201592 10406 201644 10412
rect 201500 10396 201552 10402
rect 201500 10338 201552 10344
rect 200304 4888 200356 4894
rect 200304 4830 200356 4836
rect 201408 4888 201460 4894
rect 201408 4830 201460 4836
rect 200316 480 200344 4830
rect 201512 4010 201540 10338
rect 201408 4004 201460 4010
rect 201408 3946 201460 3952
rect 201500 4004 201552 4010
rect 201500 3946 201552 3952
rect 201420 3126 201448 3946
rect 201604 3482 201632 10406
rect 202432 5234 202460 56646
rect 202524 10674 202552 57666
rect 202708 57610 202736 60044
rect 202616 57582 202736 57610
rect 202512 10668 202564 10674
rect 202512 10610 202564 10616
rect 202616 10606 202644 57582
rect 202696 56908 202748 56914
rect 202696 56850 202748 56856
rect 202604 10600 202656 10606
rect 202604 10542 202656 10548
rect 202420 5228 202472 5234
rect 202420 5170 202472 5176
rect 202708 5166 202736 56850
rect 202984 55894 203012 60044
rect 203260 56914 203288 60044
rect 203536 57730 203564 60044
rect 203524 57724 203576 57730
rect 203524 57666 203576 57672
rect 203904 57066 203932 60044
rect 203984 57724 204036 57730
rect 203984 57666 204036 57672
rect 203812 57038 203932 57066
rect 203248 56908 203300 56914
rect 203248 56850 203300 56856
rect 203812 56846 203840 57038
rect 203892 56908 203944 56914
rect 203892 56850 203944 56856
rect 203156 56840 203208 56846
rect 203156 56782 203208 56788
rect 203800 56840 203852 56846
rect 203800 56782 203852 56788
rect 202972 55888 203024 55894
rect 202972 55830 203024 55836
rect 203168 54534 203196 56782
rect 203156 54528 203208 54534
rect 203156 54470 203208 54476
rect 202696 5160 202748 5166
rect 202696 5102 202748 5108
rect 203904 5098 203932 56850
rect 203996 10538 204024 57666
rect 204180 45554 204208 60044
rect 204456 56914 204484 60044
rect 204444 56908 204496 56914
rect 204444 56850 204496 56856
rect 204732 50522 204760 60044
rect 205100 57730 205128 60044
rect 205088 57724 205140 57730
rect 205088 57666 205140 57672
rect 205376 57610 205404 60044
rect 205548 57724 205600 57730
rect 205548 57666 205600 57672
rect 205376 57582 205496 57610
rect 205364 56908 205416 56914
rect 205364 56850 205416 56856
rect 204720 50516 204772 50522
rect 204720 50458 204772 50464
rect 204088 45526 204208 45554
rect 203984 10532 204036 10538
rect 203984 10474 204036 10480
rect 203892 5092 203944 5098
rect 203892 5034 203944 5040
rect 204088 4962 204116 45526
rect 205376 10470 205404 56850
rect 205364 10464 205416 10470
rect 205364 10406 205416 10412
rect 205468 10402 205496 57582
rect 205456 10396 205508 10402
rect 205456 10338 205508 10344
rect 205088 10328 205140 10334
rect 205088 10270 205140 10276
rect 204996 5024 205048 5030
rect 204996 4966 205048 4972
rect 204076 4956 204128 4962
rect 204076 4898 204128 4904
rect 203892 4820 203944 4826
rect 203892 4762 203944 4768
rect 202696 4004 202748 4010
rect 202696 3946 202748 3952
rect 201512 3454 201632 3482
rect 201408 3120 201460 3126
rect 201408 3062 201460 3068
rect 201512 480 201540 3454
rect 202708 480 202736 3946
rect 203904 480 203932 4762
rect 205008 4554 205036 4966
rect 204996 4548 205048 4554
rect 204996 4490 205048 4496
rect 205100 480 205128 10270
rect 205560 4894 205588 57666
rect 205652 56914 205680 60044
rect 205640 56908 205692 56914
rect 205640 56850 205692 56856
rect 205928 56846 205956 60044
rect 206296 57730 206324 60044
rect 206284 57724 206336 57730
rect 206284 57666 206336 57672
rect 206572 57610 206600 60044
rect 206848 57882 206876 60044
rect 206848 57854 206968 57882
rect 206836 57724 206888 57730
rect 206836 57666 206888 57672
rect 206572 57582 206784 57610
rect 206652 56908 206704 56914
rect 206652 56850 206704 56856
rect 205916 56840 205968 56846
rect 205916 56782 205968 56788
rect 206664 15978 206692 56850
rect 206652 15972 206704 15978
rect 206652 15914 206704 15920
rect 206756 15910 206784 57582
rect 206744 15904 206796 15910
rect 206744 15846 206796 15852
rect 206848 10334 206876 57666
rect 206940 57225 206968 57854
rect 207124 57730 207152 60044
rect 207112 57724 207164 57730
rect 207112 57666 207164 57672
rect 206926 57216 206982 57225
rect 206926 57151 206982 57160
rect 207492 56914 207520 60044
rect 207768 58002 207796 60044
rect 207756 57996 207808 58002
rect 207756 57938 207808 57944
rect 208044 57633 208072 60044
rect 208320 58698 208348 60044
rect 208136 58670 208348 58698
rect 208030 57624 208086 57633
rect 208030 57559 208086 57568
rect 207480 56908 207532 56914
rect 207480 56850 207532 56856
rect 208136 56846 208164 58670
rect 208688 58070 208716 60044
rect 208964 58546 208992 60044
rect 209240 58818 209268 60044
rect 209228 58812 209280 58818
rect 209228 58754 209280 58760
rect 208952 58540 209004 58546
rect 208952 58482 209004 58488
rect 209516 58410 209544 60044
rect 209884 59158 209912 60044
rect 209872 59152 209924 59158
rect 209872 59094 209924 59100
rect 210160 58993 210188 60044
rect 210146 58984 210202 58993
rect 210146 58919 210202 58928
rect 209504 58404 209556 58410
rect 209504 58346 209556 58352
rect 208676 58064 208728 58070
rect 208676 58006 208728 58012
rect 208308 57996 208360 58002
rect 208308 57938 208360 57944
rect 208320 57730 208348 57938
rect 208216 57724 208268 57730
rect 208216 57666 208268 57672
rect 208308 57724 208360 57730
rect 208308 57666 208360 57672
rect 206928 56840 206980 56846
rect 206928 56782 206980 56788
rect 208124 56840 208176 56846
rect 208124 56782 208176 56788
rect 206836 10328 206888 10334
rect 206836 10270 206888 10276
rect 205824 5228 205876 5234
rect 205824 5170 205876 5176
rect 205548 4888 205600 4894
rect 205548 4830 205600 4836
rect 205836 4826 205864 5170
rect 206940 4826 206968 56782
rect 208228 11801 208256 57666
rect 210436 56914 210464 60044
rect 210712 58614 210740 60044
rect 210700 58608 210752 58614
rect 210700 58550 210752 58556
rect 211080 57769 211108 60044
rect 211356 58886 211384 60044
rect 211344 58880 211396 58886
rect 211344 58822 211396 58828
rect 211066 57760 211122 57769
rect 211066 57695 211122 57704
rect 211632 56953 211660 60044
rect 211618 56944 211674 56953
rect 208308 56908 208360 56914
rect 208308 56850 208360 56856
rect 210424 56908 210476 56914
rect 211618 56879 211674 56888
rect 210424 56850 210476 56856
rect 208214 11792 208270 11801
rect 208214 11727 208270 11736
rect 208320 11665 208348 56850
rect 211908 56817 211936 60044
rect 212276 58682 212304 60044
rect 212552 59129 212580 60044
rect 212538 59120 212594 59129
rect 212538 59055 212594 59064
rect 212264 58676 212316 58682
rect 212264 58618 212316 58624
rect 212828 57905 212856 60044
rect 212814 57896 212870 57905
rect 212814 57831 212870 57840
rect 213196 57089 213224 60044
rect 213182 57080 213238 57089
rect 213182 57015 213238 57024
rect 211894 56808 211950 56817
rect 211894 56743 211950 56752
rect 209044 56704 209096 56710
rect 209044 56646 209096 56652
rect 209056 18630 209084 56646
rect 213472 56642 213500 60044
rect 213748 57361 213776 60044
rect 213734 57352 213790 57361
rect 213734 57287 213790 57296
rect 214024 56710 214052 60044
rect 214392 58750 214420 60044
rect 214380 58744 214432 58750
rect 214380 58686 214432 58692
rect 214668 57497 214696 60044
rect 214944 58478 214972 60044
rect 214932 58472 214984 58478
rect 214932 58414 214984 58420
rect 215220 57769 215248 60044
rect 215588 58138 215616 60044
rect 215864 59022 215892 60044
rect 216140 59809 216168 60044
rect 216126 59800 216182 59809
rect 216126 59735 216182 59744
rect 215852 59016 215904 59022
rect 215852 58958 215904 58964
rect 216416 58342 216444 60044
rect 216784 59090 216812 60044
rect 217060 59362 217088 60044
rect 217048 59356 217100 59362
rect 217048 59298 217100 59304
rect 216772 59084 216824 59090
rect 216772 59026 216824 59032
rect 216404 58336 216456 58342
rect 216404 58278 216456 58284
rect 215576 58132 215628 58138
rect 215576 58074 215628 58080
rect 216588 57996 216640 58002
rect 216588 57938 216640 57944
rect 216600 57798 216628 57938
rect 216588 57792 216640 57798
rect 215206 57760 215262 57769
rect 216588 57734 216640 57740
rect 216680 57792 216732 57798
rect 216680 57734 216732 57740
rect 215206 57695 215262 57704
rect 214654 57488 214710 57497
rect 214654 57423 214710 57432
rect 216692 57186 216720 57734
rect 216864 57724 216916 57730
rect 216864 57666 216916 57672
rect 216680 57180 216732 57186
rect 216680 57122 216732 57128
rect 216876 57118 216904 57666
rect 217336 57202 217364 60044
rect 217612 59537 217640 60044
rect 217598 59528 217654 59537
rect 217598 59463 217654 59472
rect 217980 59362 218008 60044
rect 218256 59945 218284 60044
rect 218242 59936 218298 59945
rect 218242 59871 218298 59880
rect 217968 59356 218020 59362
rect 217968 59298 218020 59304
rect 218532 58274 218560 60044
rect 218520 58268 218572 58274
rect 218520 58210 218572 58216
rect 218244 57792 218296 57798
rect 218428 57792 218480 57798
rect 218296 57740 218428 57746
rect 218244 57734 218480 57740
rect 218256 57718 218468 57734
rect 217336 57174 217548 57202
rect 216864 57112 216916 57118
rect 216864 57054 216916 57060
rect 217416 57044 217468 57050
rect 217416 56986 217468 56992
rect 217140 56976 217192 56982
rect 217428 56930 217456 56986
rect 217192 56924 217456 56930
rect 217140 56918 217456 56924
rect 217152 56902 217456 56918
rect 214012 56704 214064 56710
rect 217520 56681 217548 57174
rect 218704 57180 218756 57186
rect 218704 57122 218756 57128
rect 218612 56976 218664 56982
rect 218612 56918 218664 56924
rect 214012 56646 214064 56652
rect 217506 56672 217562 56681
rect 213460 56636 213512 56642
rect 217506 56607 217562 56616
rect 213460 56578 213512 56584
rect 218624 55622 218652 56918
rect 218060 55616 218112 55622
rect 218060 55558 218112 55564
rect 218612 55616 218664 55622
rect 218612 55558 218664 55564
rect 213920 55480 213972 55486
rect 213920 55422 213972 55428
rect 209780 55412 209832 55418
rect 209780 55354 209832 55360
rect 209044 18624 209096 18630
rect 209044 18566 209096 18572
rect 208306 11656 208362 11665
rect 208306 11591 208362 11600
rect 209792 11082 209820 55354
rect 213932 16574 213960 55422
rect 213932 16546 214512 16574
rect 213368 15428 213420 15434
rect 213368 15370 213420 15376
rect 209872 15360 209924 15366
rect 209872 15302 209924 15308
rect 209780 11076 209832 11082
rect 209780 11018 209832 11024
rect 208584 9784 208636 9790
rect 208584 9726 208636 9732
rect 205824 4820 205876 4826
rect 205824 4762 205876 4768
rect 206928 4820 206980 4826
rect 206928 4762 206980 4768
rect 206192 3256 206244 3262
rect 206192 3198 206244 3204
rect 206204 480 206232 3198
rect 207388 3120 207440 3126
rect 207388 3062 207440 3068
rect 207400 480 207428 3062
rect 208596 480 208624 9726
rect 209884 3482 209912 15302
rect 210976 11076 211028 11082
rect 210976 11018 211028 11024
rect 209792 3454 209912 3482
rect 209792 480 209820 3454
rect 210988 480 211016 11018
rect 212172 9852 212224 9858
rect 212172 9794 212224 9800
rect 212184 480 212212 9794
rect 213380 480 213408 15370
rect 214484 480 214512 16546
rect 216864 15496 216916 15502
rect 216864 15438 216916 15444
rect 215668 9920 215720 9926
rect 215668 9862 215720 9868
rect 215680 480 215708 9862
rect 216876 480 216904 15438
rect 218072 480 218100 55558
rect 218612 9988 218664 9994
rect 218612 9930 218664 9936
rect 218624 3074 218652 9930
rect 218716 3262 218744 57122
rect 218808 56982 218836 60044
rect 219176 58954 219204 60044
rect 219164 58948 219216 58954
rect 219164 58890 219216 58896
rect 218888 57928 218940 57934
rect 218888 57870 218940 57876
rect 218980 57928 219032 57934
rect 218980 57870 219032 57876
rect 218796 56976 218848 56982
rect 218796 56918 218848 56924
rect 218900 3890 218928 57870
rect 218992 57186 219020 57870
rect 219452 57866 219480 60044
rect 219728 58857 219756 60044
rect 220004 59265 220032 60044
rect 219990 59256 220046 59265
rect 219990 59191 220046 59200
rect 219714 58848 219770 58857
rect 219714 58783 219770 58792
rect 220372 57934 220400 60044
rect 220648 58206 220676 60044
rect 220924 59294 220952 60044
rect 221200 59673 221228 60044
rect 221186 59664 221242 59673
rect 221186 59599 221242 59608
rect 220912 59288 220964 59294
rect 220912 59230 220964 59236
rect 221568 59226 221596 60044
rect 221556 59220 221608 59226
rect 221556 59162 221608 59168
rect 220636 58200 220688 58206
rect 220636 58142 220688 58148
rect 220360 57928 220412 57934
rect 220360 57870 220412 57876
rect 219440 57860 219492 57866
rect 219440 57802 219492 57808
rect 221648 57792 221700 57798
rect 221648 57734 221700 57740
rect 221464 57724 221516 57730
rect 221464 57666 221516 57672
rect 218980 57180 219032 57186
rect 218980 57122 219032 57128
rect 218980 57044 219032 57050
rect 218980 56986 219032 56992
rect 218992 4010 219020 56986
rect 220820 55684 220872 55690
rect 220820 55626 220872 55632
rect 219072 55616 219124 55622
rect 219072 55558 219124 55564
rect 219084 6089 219112 55558
rect 220832 16574 220860 55626
rect 220832 16546 221412 16574
rect 220452 15564 220504 15570
rect 220452 15506 220504 15512
rect 219070 6080 219126 6089
rect 219070 6015 219126 6024
rect 218980 4004 219032 4010
rect 218980 3946 219032 3952
rect 218900 3862 219388 3890
rect 218704 3256 218756 3262
rect 218704 3198 218756 3204
rect 218624 3046 219296 3074
rect 219360 3058 219388 3862
rect 219268 480 219296 3046
rect 219348 3052 219400 3058
rect 219348 2994 219400 3000
rect 220464 480 220492 15506
rect 221384 2802 221412 16546
rect 221476 2990 221504 57666
rect 221556 57180 221608 57186
rect 221556 57122 221608 57128
rect 221464 2984 221516 2990
rect 221464 2926 221516 2932
rect 221568 2922 221596 57122
rect 221660 3126 221688 57734
rect 221844 57730 221872 60044
rect 222120 59906 222148 60044
rect 222396 59945 222424 60044
rect 222382 59936 222438 59945
rect 222108 59900 222160 59906
rect 222382 59871 222438 59880
rect 222108 59842 222160 59848
rect 222568 59832 222620 59838
rect 222566 59800 222568 59809
rect 222764 59809 222792 60044
rect 222620 59800 222622 59809
rect 222566 59735 222622 59744
rect 222750 59800 222806 59809
rect 222750 59735 222806 59744
rect 223040 59401 223068 60044
rect 223026 59392 223082 59401
rect 223026 59327 223082 59336
rect 223316 57798 223344 60044
rect 223592 59498 223620 60044
rect 223960 59945 223988 60044
rect 223946 59936 224002 59945
rect 223946 59871 224002 59880
rect 224130 59936 224186 59945
rect 224130 59871 224186 59880
rect 224144 59838 224172 59871
rect 224132 59832 224184 59838
rect 224132 59774 224184 59780
rect 224236 59770 224264 60044
rect 224316 59832 224368 59838
rect 224316 59774 224368 59780
rect 224224 59764 224276 59770
rect 224224 59706 224276 59712
rect 223580 59492 223632 59498
rect 223580 59434 223632 59440
rect 223304 57792 223356 57798
rect 223304 57734 223356 57740
rect 221832 57724 221884 57730
rect 221832 57666 221884 57672
rect 224328 57361 224356 59774
rect 224512 59430 224540 60044
rect 224788 59770 224816 261122
rect 224880 223145 224908 395490
rect 224866 223136 224922 223145
rect 224866 223071 224922 223080
rect 224776 59764 224828 59770
rect 224776 59706 224828 59712
rect 224500 59424 224552 59430
rect 224500 59366 224552 59372
rect 224972 58070 225000 398686
rect 225236 398608 225288 398614
rect 225236 398550 225288 398556
rect 225144 398268 225196 398274
rect 225144 398210 225196 398216
rect 225052 398200 225104 398206
rect 225052 398142 225104 398148
rect 225064 58857 225092 398142
rect 225156 193769 225184 398210
rect 225248 198665 225276 398550
rect 225880 266144 225932 266150
rect 225880 266086 225932 266092
rect 225604 266076 225656 266082
rect 225604 266018 225656 266024
rect 225512 262812 225564 262818
rect 225512 262754 225564 262760
rect 225326 249112 225382 249121
rect 225326 249047 225382 249056
rect 225234 198656 225290 198665
rect 225234 198591 225290 198600
rect 225142 193760 225198 193769
rect 225142 193695 225198 193704
rect 225050 58848 225106 58857
rect 225050 58783 225106 58792
rect 224960 58064 225012 58070
rect 224960 58006 225012 58012
rect 225340 57934 225368 249047
rect 225418 238096 225474 238105
rect 225418 238031 225474 238040
rect 225328 57928 225380 57934
rect 225328 57870 225380 57876
rect 225432 57866 225460 238031
rect 225524 220697 225552 262754
rect 225510 220688 225566 220697
rect 225510 220623 225566 220632
rect 225616 93129 225644 266018
rect 225694 228712 225750 228721
rect 225694 228647 225750 228656
rect 225602 93120 225658 93129
rect 225602 93055 225658 93064
rect 225420 57860 225472 57866
rect 225420 57802 225472 57808
rect 224314 57352 224370 57361
rect 224314 57287 224370 57296
rect 225708 57118 225736 228647
rect 225786 228576 225842 228585
rect 225786 228511 225842 228520
rect 225696 57112 225748 57118
rect 225696 57054 225748 57060
rect 225800 56642 225828 228511
rect 225892 134881 225920 266086
rect 225970 247616 226026 247625
rect 225970 247551 226026 247560
rect 225984 152017 226012 247551
rect 226062 235376 226118 235385
rect 226062 235311 226118 235320
rect 226076 164257 226104 235311
rect 226246 234016 226302 234025
rect 226246 233951 226302 233960
rect 226154 232520 226210 232529
rect 226154 232455 226210 232464
rect 226168 213353 226196 232455
rect 226154 213344 226210 213353
rect 226154 213279 226210 213288
rect 226062 164248 226118 164257
rect 226062 164183 226118 164192
rect 225970 152008 226026 152017
rect 225970 151943 226026 151952
rect 225878 134872 225934 134881
rect 225878 134807 225934 134816
rect 226260 56817 226288 233951
rect 226352 88233 226380 399978
rect 226524 399968 226576 399974
rect 226524 399910 226576 399916
rect 226432 399424 226484 399430
rect 226432 399366 226484 399372
rect 226444 120193 226472 399366
rect 226536 159361 226564 399910
rect 226616 398540 226668 398546
rect 226616 398482 226668 398488
rect 226628 176633 226656 398482
rect 226720 183977 226748 399978
rect 231860 399900 231912 399906
rect 231860 399842 231912 399848
rect 230756 399696 230808 399702
rect 230756 399638 230808 399644
rect 230572 397316 230624 397322
rect 230572 397258 230624 397264
rect 229284 397112 229336 397118
rect 229284 397054 229336 397060
rect 229100 396500 229152 396506
rect 229100 396442 229152 396448
rect 227720 396432 227772 396438
rect 227720 396374 227772 396380
rect 226892 260568 226944 260574
rect 226892 260510 226944 260516
rect 226798 227216 226854 227225
rect 226798 227151 226854 227160
rect 226706 183968 226762 183977
rect 226706 183903 226762 183912
rect 226614 176624 226670 176633
rect 226614 176559 226670 176568
rect 226614 175264 226670 175273
rect 226614 175199 226670 175208
rect 226628 174185 226656 175199
rect 226614 174176 226670 174185
rect 226614 174111 226670 174120
rect 226522 159352 226578 159361
rect 226522 159287 226578 159296
rect 226522 150376 226578 150385
rect 226522 150311 226578 150320
rect 226536 149569 226564 150311
rect 226522 149560 226578 149569
rect 226522 149495 226578 149504
rect 226522 140720 226578 140729
rect 226522 140655 226578 140664
rect 226536 139777 226564 140655
rect 226522 139768 226578 139777
rect 226522 139703 226578 139712
rect 226430 120184 226486 120193
rect 226430 120119 226486 120128
rect 226338 88224 226394 88233
rect 226338 88159 226394 88168
rect 226522 84144 226578 84153
rect 226522 84079 226578 84088
rect 226536 83337 226564 84079
rect 226522 83328 226578 83337
rect 226522 83263 226578 83272
rect 226522 77208 226578 77217
rect 226522 77143 226578 77152
rect 226536 75993 226564 77143
rect 226522 75984 226578 75993
rect 226522 75919 226578 75928
rect 226812 71097 226840 227151
rect 226904 154465 226932 260510
rect 227166 250472 227222 250481
rect 227166 250407 227222 250416
rect 226982 231296 227038 231305
rect 226982 231231 227038 231240
rect 226890 154456 226946 154465
rect 226890 154391 226946 154400
rect 226996 144673 227024 231231
rect 227074 225992 227130 226001
rect 227074 225927 227130 225936
rect 226982 144664 227038 144673
rect 226982 144599 227038 144608
rect 227088 142225 227116 225927
rect 227180 171601 227208 250407
rect 227350 239456 227406 239465
rect 227350 239391 227406 239400
rect 227258 227352 227314 227361
rect 227258 227287 227314 227296
rect 227166 171592 227222 171601
rect 227166 171527 227222 171536
rect 227272 166705 227300 227287
rect 227364 188873 227392 239391
rect 227534 234288 227590 234297
rect 227534 234223 227590 234232
rect 227442 229800 227498 229809
rect 227442 229735 227498 229744
rect 227350 188864 227406 188873
rect 227350 188799 227406 188808
rect 227456 181529 227484 229735
rect 227548 196217 227576 234223
rect 227626 231432 227682 231441
rect 227626 231367 227682 231376
rect 227640 215801 227668 231367
rect 227626 215792 227682 215801
rect 227626 215727 227682 215736
rect 227626 209672 227682 209681
rect 227626 209607 227682 209616
rect 227640 208457 227668 209607
rect 227626 208448 227682 208457
rect 227626 208383 227682 208392
rect 227534 196208 227590 196217
rect 227534 196143 227590 196152
rect 227442 181520 227498 181529
rect 227442 181455 227498 181464
rect 227258 166696 227314 166705
rect 227258 166631 227314 166640
rect 227074 142216 227130 142225
rect 227074 142151 227130 142160
rect 226798 71088 226854 71097
rect 226798 71023 226854 71032
rect 226522 64832 226578 64841
rect 226522 64767 226578 64776
rect 226536 63753 226564 64767
rect 226522 63744 226578 63753
rect 226522 63679 226578 63688
rect 227732 58750 227760 396374
rect 227996 395820 228048 395826
rect 227996 395762 228048 395768
rect 227812 395616 227864 395622
rect 227812 395558 227864 395564
rect 227824 179081 227852 395558
rect 227904 264512 227956 264518
rect 227904 264454 227956 264460
rect 227810 179072 227866 179081
rect 227810 179007 227866 179016
rect 227916 68649 227944 264454
rect 228008 210905 228036 395762
rect 228548 264716 228600 264722
rect 228548 264658 228600 264664
rect 228364 263560 228416 263566
rect 228364 263502 228416 263508
rect 228086 240952 228142 240961
rect 228086 240887 228142 240896
rect 227994 210896 228050 210905
rect 227994 210831 228050 210840
rect 227902 68640 227958 68649
rect 227902 68575 227958 68584
rect 227720 58744 227772 58750
rect 227720 58686 227772 58692
rect 226984 57928 227036 57934
rect 226984 57870 227036 57876
rect 226996 57730 227024 57870
rect 228100 57769 228128 240887
rect 228178 234152 228234 234161
rect 228178 234087 228234 234096
rect 228086 57760 228142 57769
rect 226984 57724 227036 57730
rect 228086 57695 228142 57704
rect 226984 57666 227036 57672
rect 228192 57633 228220 234087
rect 228270 232656 228326 232665
rect 228270 232591 228326 232600
rect 228178 57624 228234 57633
rect 228178 57559 228234 57568
rect 226246 56808 226302 56817
rect 226246 56743 226302 56752
rect 228284 56710 228312 232591
rect 228376 105369 228404 263502
rect 228456 260500 228508 260506
rect 228456 260442 228508 260448
rect 228468 112713 228496 260442
rect 228560 169153 228588 264658
rect 228640 261316 228692 261322
rect 228640 261258 228692 261264
rect 228652 186425 228680 261258
rect 228638 186416 228694 186425
rect 228638 186351 228694 186360
rect 228546 169144 228602 169153
rect 228546 169079 228602 169088
rect 228454 112704 228510 112713
rect 228454 112639 228510 112648
rect 228362 105360 228418 105369
rect 228362 105295 228418 105304
rect 229112 59362 229140 396442
rect 229192 396364 229244 396370
rect 229192 396306 229244 396312
rect 229100 59356 229152 59362
rect 229100 59298 229152 59304
rect 229204 59022 229232 396306
rect 229296 59090 229324 397054
rect 230480 396636 230532 396642
rect 230480 396578 230532 396584
rect 229376 396568 229428 396574
rect 229376 396510 229428 396516
rect 229388 59294 229416 396510
rect 229468 264648 229520 264654
rect 229468 264590 229520 264596
rect 229376 59288 229428 59294
rect 229376 59230 229428 59236
rect 229284 59084 229336 59090
rect 229284 59026 229336 59032
rect 229192 59016 229244 59022
rect 229192 58958 229244 58964
rect 228272 56704 228324 56710
rect 229480 56681 229508 264590
rect 229652 262132 229704 262138
rect 229652 262074 229704 262080
rect 229560 260840 229612 260846
rect 229560 260782 229612 260788
rect 229572 56914 229600 260782
rect 229664 147121 229692 262074
rect 229834 239592 229890 239601
rect 229834 239527 229890 239536
rect 229742 231160 229798 231169
rect 229742 231095 229798 231104
rect 229650 147112 229706 147121
rect 229650 147047 229706 147056
rect 229756 117745 229784 231095
rect 229848 203561 229876 239527
rect 229926 236872 229982 236881
rect 229926 236807 229982 236816
rect 229940 218249 229968 236807
rect 229926 218240 229982 218249
rect 229926 218175 229982 218184
rect 229834 203552 229890 203561
rect 229834 203487 229890 203496
rect 229742 117736 229798 117745
rect 229742 117671 229798 117680
rect 230492 59226 230520 396578
rect 230480 59220 230532 59226
rect 230480 59162 230532 59168
rect 230584 58614 230612 397258
rect 230664 397180 230716 397186
rect 230664 397122 230716 397128
rect 230676 59158 230704 397122
rect 230768 61305 230796 399638
rect 230848 396772 230900 396778
rect 230848 396714 230900 396720
rect 230754 61296 230810 61305
rect 230754 61231 230810 61240
rect 230860 59401 230888 396714
rect 230940 396704 230992 396710
rect 230940 396646 230992 396652
rect 230952 60217 230980 396646
rect 231032 396296 231084 396302
rect 231032 396238 231084 396244
rect 230938 60208 230994 60217
rect 230938 60143 230994 60152
rect 231044 59673 231072 396238
rect 231124 266008 231176 266014
rect 231124 265950 231176 265956
rect 231136 78441 231164 265950
rect 231308 264580 231360 264586
rect 231308 264522 231360 264528
rect 231214 238232 231270 238241
rect 231214 238167 231270 238176
rect 231122 78432 231178 78441
rect 231122 78367 231178 78376
rect 231030 59664 231086 59673
rect 231030 59599 231086 59608
rect 230846 59392 230902 59401
rect 230846 59327 230902 59336
rect 230664 59152 230716 59158
rect 230664 59094 230716 59100
rect 230572 58608 230624 58614
rect 230572 58550 230624 58556
rect 231228 57497 231256 238167
rect 231320 161809 231348 264522
rect 231400 263560 231452 263566
rect 231400 263502 231452 263508
rect 231412 206009 231440 263502
rect 231398 206000 231454 206009
rect 231398 205935 231454 205944
rect 231306 161800 231362 161809
rect 231306 161735 231362 161744
rect 231872 85785 231900 399842
rect 232136 399832 232188 399838
rect 232136 399774 232188 399780
rect 232044 399628 232096 399634
rect 232044 399570 232096 399576
rect 231952 399560 232004 399566
rect 231952 399502 232004 399508
rect 231964 98025 231992 399502
rect 232056 122641 232084 399570
rect 232148 127537 232176 399774
rect 233240 399764 233292 399770
rect 233240 399706 233292 399712
rect 232228 399492 232280 399498
rect 232228 399434 232280 399440
rect 232240 129985 232268 399434
rect 232320 398132 232372 398138
rect 232320 398074 232372 398080
rect 232332 137329 232360 398074
rect 232504 261316 232556 261322
rect 232504 261258 232556 261264
rect 232410 242312 232466 242321
rect 232410 242247 232466 242256
rect 232318 137320 232374 137329
rect 232318 137255 232374 137264
rect 232226 129976 232282 129985
rect 232226 129911 232282 129920
rect 232134 127528 232190 127537
rect 232134 127463 232190 127472
rect 232042 122632 232098 122641
rect 232042 122567 232098 122576
rect 231950 98016 232006 98025
rect 231950 97951 232006 97960
rect 231858 85776 231914 85785
rect 231858 85711 231914 85720
rect 232424 66201 232452 242247
rect 232516 140729 232544 261258
rect 232502 140720 232558 140729
rect 232502 140655 232558 140664
rect 233252 95577 233280 399706
rect 244924 399560 244976 399566
rect 244924 399502 244976 399508
rect 242256 399492 242308 399498
rect 242256 399434 242308 399440
rect 235998 398168 236054 398177
rect 235998 398103 236054 398112
rect 235264 396364 235316 396370
rect 235264 396306 235316 396312
rect 233976 396296 234028 396302
rect 233976 396238 234028 396244
rect 233884 395548 233936 395554
rect 233884 395490 233936 395496
rect 233238 95568 233294 95577
rect 233238 95503 233294 95512
rect 232410 66192 232466 66201
rect 232410 66127 232466 66136
rect 231214 57488 231270 57497
rect 231214 57423 231270 57432
rect 229560 56908 229612 56914
rect 229560 56850 229612 56856
rect 233896 56846 233924 395490
rect 233988 110265 234016 396238
rect 234252 262812 234304 262818
rect 234252 262754 234304 262760
rect 234160 260500 234212 260506
rect 234160 260442 234212 260448
rect 234066 226808 234122 226817
rect 234066 226743 234122 226752
rect 233974 110256 234030 110265
rect 233974 110191 234030 110200
rect 233884 56840 233936 56846
rect 233884 56782 233936 56788
rect 228272 56646 228324 56652
rect 229466 56672 229522 56681
rect 225788 56636 225840 56642
rect 229466 56607 229522 56616
rect 225788 56578 225840 56584
rect 231860 55752 231912 55758
rect 231860 55694 231912 55700
rect 227720 55548 227772 55554
rect 227720 55490 227772 55496
rect 224960 17128 225012 17134
rect 224960 17070 225012 17076
rect 224972 16574 225000 17070
rect 227732 16574 227760 55490
rect 231872 16574 231900 55694
rect 233240 52896 233292 52902
rect 233240 52838 233292 52844
rect 233252 16574 233280 52838
rect 234080 20670 234108 226743
rect 234172 175273 234200 260442
rect 234264 191321 234292 262754
rect 234434 228440 234490 228449
rect 234434 228375 234490 228384
rect 234342 227080 234398 227089
rect 234342 227015 234398 227024
rect 234356 205737 234384 227015
rect 234448 218113 234476 228375
rect 234434 218104 234490 218113
rect 234434 218039 234490 218048
rect 235276 209681 235304 396306
rect 235448 262132 235500 262138
rect 235448 262074 235500 262080
rect 235354 230752 235410 230761
rect 235354 230687 235410 230696
rect 235262 209672 235318 209681
rect 235262 209607 235318 209616
rect 234342 205728 234398 205737
rect 234342 205663 234398 205672
rect 234250 191312 234306 191321
rect 234250 191247 234306 191256
rect 234158 175264 234214 175273
rect 234158 175199 234214 175208
rect 235262 120728 235318 120737
rect 235262 120663 235318 120672
rect 235276 100473 235304 120663
rect 235262 100464 235318 100473
rect 235262 100399 235318 100408
rect 235368 85649 235396 230687
rect 235460 150385 235488 262074
rect 235538 226944 235594 226953
rect 235538 226879 235594 226888
rect 235552 151881 235580 226879
rect 235538 151872 235594 151881
rect 235538 151807 235594 151816
rect 235446 150376 235502 150385
rect 235446 150311 235502 150320
rect 235354 85640 235410 85649
rect 235354 85575 235410 85584
rect 236012 58546 236040 398103
rect 236182 397352 236238 397361
rect 236182 397287 236238 397296
rect 239218 397352 239274 397361
rect 239218 397287 239274 397296
rect 236196 396914 236224 397287
rect 239232 397254 239260 397287
rect 239220 397248 239272 397254
rect 239220 397190 239272 397196
rect 236184 396908 236236 396914
rect 236184 396850 236236 396856
rect 237378 396808 237434 396817
rect 237378 396743 237434 396752
rect 240138 396808 240194 396817
rect 240138 396743 240194 396752
rect 241518 396808 241574 396817
rect 241518 396743 241574 396752
rect 236642 230888 236698 230897
rect 236642 230823 236698 230832
rect 236656 125633 236684 230823
rect 236734 228168 236790 228177
rect 236734 228103 236790 228112
rect 236748 178129 236776 228103
rect 236734 178120 236790 178129
rect 236734 178055 236790 178064
rect 236642 125624 236698 125633
rect 236642 125559 236698 125568
rect 237392 58818 237420 396743
rect 237472 396160 237524 396166
rect 237472 396102 237524 396108
rect 237484 393990 237512 396102
rect 238024 394052 238076 394058
rect 238024 393994 238076 394000
rect 237472 393984 237524 393990
rect 237472 393926 237524 393932
rect 238036 125089 238064 393994
rect 238208 261248 238260 261254
rect 238208 261190 238260 261196
rect 238114 226536 238170 226545
rect 238114 226471 238170 226480
rect 238022 125080 238078 125089
rect 238022 125015 238078 125024
rect 237380 58812 237432 58818
rect 237380 58754 237432 58760
rect 236000 58540 236052 58546
rect 236000 58482 236052 58488
rect 238128 33114 238156 226471
rect 238220 102921 238248 261190
rect 238300 260568 238352 260574
rect 238300 260510 238352 260516
rect 238312 201113 238340 260510
rect 239402 228032 239458 228041
rect 239402 227967 239458 227976
rect 238298 201104 238354 201113
rect 238298 201039 238354 201048
rect 239416 138145 239444 227967
rect 239402 138136 239458 138145
rect 239402 138071 239458 138080
rect 238206 102912 238262 102921
rect 238206 102847 238262 102856
rect 240152 58886 240180 396743
rect 240784 392692 240836 392698
rect 240784 392634 240836 392640
rect 240796 157321 240824 392634
rect 240874 227896 240930 227905
rect 240874 227831 240930 227840
rect 240782 157312 240838 157321
rect 240782 157247 240838 157256
rect 240888 59906 240916 227831
rect 241532 120737 241560 396743
rect 242164 396704 242216 396710
rect 242164 396646 242216 396652
rect 241518 120728 241574 120737
rect 241518 120663 241574 120672
rect 242176 84153 242204 396646
rect 242268 91089 242296 399434
rect 242898 396808 242954 396817
rect 242898 396743 242954 396752
rect 244370 396808 244426 396817
rect 244370 396743 244426 396752
rect 244554 396808 244610 396817
rect 244554 396743 244610 396752
rect 242912 242185 242940 396743
rect 242898 242176 242954 242185
rect 242898 242111 242954 242120
rect 242254 91080 242310 91089
rect 242254 91015 242310 91024
rect 242162 84144 242218 84153
rect 242162 84079 242218 84088
rect 240876 59900 240928 59906
rect 240876 59842 240928 59848
rect 240140 58880 240192 58886
rect 240140 58822 240192 58828
rect 244384 58410 244412 396743
rect 244568 396710 244596 396743
rect 244556 396704 244608 396710
rect 244556 396646 244608 396652
rect 244936 64841 244964 399502
rect 265070 398168 265126 398177
rect 265070 398103 265126 398112
rect 300122 398168 300178 398177
rect 300122 398103 300178 398112
rect 315762 398168 315818 398177
rect 315762 398103 315818 398112
rect 325882 398168 325938 398177
rect 325882 398103 325938 398112
rect 247682 397352 247738 397361
rect 247682 397287 247738 397296
rect 247958 397352 248014 397361
rect 247958 397287 248014 397296
rect 248602 397352 248658 397361
rect 248602 397287 248658 397296
rect 250074 397352 250130 397361
rect 250074 397287 250130 397296
rect 250350 397352 250406 397361
rect 250350 397287 250406 397296
rect 252742 397352 252798 397361
rect 252742 397287 252798 397296
rect 259458 397352 259514 397361
rect 259458 397287 259514 397296
rect 260930 397352 260986 397361
rect 260930 397287 260986 397296
rect 261942 397352 261998 397361
rect 261942 397287 261998 397296
rect 262310 397352 262366 397361
rect 262310 397287 262366 397296
rect 263598 397352 263654 397361
rect 263598 397287 263654 397296
rect 245658 396808 245714 396817
rect 245658 396743 245714 396752
rect 244922 64832 244978 64841
rect 244922 64767 244978 64776
rect 245672 58682 245700 396743
rect 246304 396500 246356 396506
rect 246304 396442 246356 396448
rect 246316 264042 246344 396442
rect 247696 396302 247724 397287
rect 247684 396296 247736 396302
rect 247684 396238 247736 396244
rect 247972 395554 248000 397287
rect 248616 396166 248644 397287
rect 250088 396982 250116 397287
rect 250076 396976 250128 396982
rect 250076 396918 250128 396924
rect 249064 396704 249116 396710
rect 249064 396646 249116 396652
rect 248604 396160 248656 396166
rect 248604 396102 248656 396108
rect 247960 395548 248012 395554
rect 247960 395490 248012 395496
rect 246304 264036 246356 264042
rect 246304 263978 246356 263984
rect 246302 226672 246358 226681
rect 246302 226607 246358 226616
rect 246316 165753 246344 226607
rect 246302 165744 246358 165753
rect 246302 165679 246358 165688
rect 249076 132433 249104 396646
rect 250364 395758 250392 397287
rect 251178 397080 251234 397089
rect 251178 397015 251234 397024
rect 250444 396772 250496 396778
rect 250444 396714 250496 396720
rect 250352 395752 250404 395758
rect 250352 395694 250404 395700
rect 249062 132424 249118 132433
rect 249062 132359 249118 132368
rect 250456 58954 250484 396714
rect 251192 394058 251220 397015
rect 252756 396846 252784 397287
rect 259472 397186 259500 397287
rect 253296 397180 253348 397186
rect 253296 397122 253348 397128
rect 259460 397180 259512 397186
rect 259460 397122 259512 397128
rect 252744 396840 252796 396846
rect 251362 396808 251418 396817
rect 251362 396743 251418 396752
rect 252558 396808 252614 396817
rect 252744 396782 252796 396788
rect 252558 396743 252614 396752
rect 251376 396710 251404 396743
rect 251364 396704 251416 396710
rect 251364 396646 251416 396652
rect 251916 396704 251968 396710
rect 251916 396646 251968 396652
rect 251824 396024 251876 396030
rect 251824 395966 251876 395972
rect 251180 394052 251232 394058
rect 251180 393994 251232 394000
rect 250444 58948 250496 58954
rect 250444 58890 250496 58896
rect 245660 58676 245712 58682
rect 245660 58618 245712 58624
rect 244372 58404 244424 58410
rect 244372 58346 244424 58352
rect 251836 56953 251864 395966
rect 251928 265538 251956 396646
rect 251916 265532 251968 265538
rect 251916 265474 251968 265480
rect 252572 264858 252600 396743
rect 253204 396296 253256 396302
rect 253204 396238 253256 396244
rect 252560 264852 252612 264858
rect 252560 264794 252612 264800
rect 251914 257952 251970 257961
rect 251914 257887 251970 257896
rect 251928 237969 251956 257887
rect 251914 237960 251970 237969
rect 251914 237895 251970 237904
rect 253216 58206 253244 396238
rect 253308 392630 253336 397122
rect 258078 396944 258134 396953
rect 258078 396879 258134 396888
rect 254122 396808 254178 396817
rect 254122 396743 254178 396752
rect 255410 396808 255466 396817
rect 255410 396743 255466 396752
rect 256146 396808 256202 396817
rect 256146 396743 256202 396752
rect 256882 396808 256938 396817
rect 256882 396743 256884 396752
rect 254136 396710 254164 396743
rect 254124 396704 254176 396710
rect 254124 396646 254176 396652
rect 253296 392624 253348 392630
rect 253296 392566 253348 392572
rect 253294 234696 253350 234705
rect 253294 234631 253350 234640
rect 253308 111897 253336 234631
rect 253294 111888 253350 111897
rect 253294 111823 253350 111832
rect 255424 58274 255452 396743
rect 255964 396160 256016 396166
rect 255964 396102 256016 396108
rect 255412 58268 255464 58274
rect 255412 58210 255464 58216
rect 253204 58200 253256 58206
rect 253204 58142 253256 58148
rect 255976 57089 256004 396102
rect 256160 396030 256188 396743
rect 256936 396743 256938 396752
rect 256884 396714 256936 396720
rect 256148 396024 256200 396030
rect 256148 395966 256200 395972
rect 258092 261254 258120 396879
rect 258170 396808 258226 396817
rect 258170 396743 258226 396752
rect 259550 396808 259606 396817
rect 259550 396743 259606 396752
rect 258184 392698 258212 396743
rect 258172 392692 258224 392698
rect 258172 392634 258224 392640
rect 258724 392624 258776 392630
rect 258724 392566 258776 392572
rect 258080 261248 258132 261254
rect 258080 261190 258132 261196
rect 255962 57080 256018 57089
rect 255962 57015 256018 57024
rect 258736 56982 258764 392566
rect 259564 265878 259592 396743
rect 260104 396432 260156 396438
rect 260104 396374 260156 396380
rect 259552 265872 259604 265878
rect 259552 265814 259604 265820
rect 260116 264178 260144 396374
rect 260944 396166 260972 397287
rect 261956 396302 261984 397287
rect 261944 396296 261996 396302
rect 261944 396238 261996 396244
rect 260932 396160 260984 396166
rect 260932 396102 260984 396108
rect 262324 395894 262352 397287
rect 262864 396772 262916 396778
rect 262864 396714 262916 396720
rect 262312 395888 262364 395894
rect 262312 395830 262364 395836
rect 260104 264172 260156 264178
rect 260104 264114 260156 264120
rect 260746 245712 260802 245721
rect 260746 245647 260802 245656
rect 260760 245614 260788 245647
rect 260748 245608 260800 245614
rect 260748 245550 260800 245556
rect 262876 58478 262904 396714
rect 263612 396506 263640 397287
rect 263690 396808 263746 396817
rect 263690 396743 263746 396752
rect 263600 396500 263652 396506
rect 263600 396442 263652 396448
rect 263704 59838 263732 396743
rect 265084 262070 265112 398103
rect 275284 397384 275336 397390
rect 268290 397352 268346 397361
rect 268290 397287 268346 397296
rect 268658 397352 268714 397361
rect 268658 397287 268714 397296
rect 272338 397352 272394 397361
rect 272338 397287 272394 397296
rect 275282 397352 275284 397361
rect 275336 397352 275338 397361
rect 275282 397287 275338 397296
rect 277674 397352 277730 397361
rect 277674 397287 277730 397296
rect 278870 397352 278926 397361
rect 278870 397287 278926 397296
rect 290186 397352 290242 397361
rect 290186 397287 290242 397296
rect 298466 397352 298522 397361
rect 298466 397287 298522 397296
rect 265162 396808 265218 396817
rect 265162 396743 265164 396752
rect 265216 396743 265218 396752
rect 266358 396808 266414 396817
rect 266358 396743 266414 396752
rect 265164 396714 265216 396720
rect 265072 262064 265124 262070
rect 265072 262006 265124 262012
rect 263692 59832 263744 59838
rect 263692 59774 263744 59780
rect 266372 59401 266400 396743
rect 266450 396672 266506 396681
rect 266450 396607 266506 396616
rect 266464 262818 266492 396607
rect 268304 395690 268332 397287
rect 268672 397050 268700 397287
rect 268660 397044 268712 397050
rect 268660 396986 268712 396992
rect 269394 396808 269450 396817
rect 268476 396772 268528 396778
rect 269394 396743 269396 396752
rect 268476 396714 268528 396720
rect 269448 396743 269450 396752
rect 270498 396808 270554 396817
rect 270498 396743 270554 396752
rect 269396 396714 269448 396720
rect 268384 396704 268436 396710
rect 268384 396646 268436 396652
rect 268292 395684 268344 395690
rect 268292 395626 268344 395632
rect 266452 262812 266504 262818
rect 266452 262754 266504 262760
rect 268396 59498 268424 396646
rect 268488 264926 268516 396714
rect 269764 396296 269816 396302
rect 269764 396238 269816 396244
rect 268476 264920 268528 264926
rect 268476 264862 268528 264868
rect 268384 59492 268436 59498
rect 268384 59434 268436 59440
rect 266358 59392 266414 59401
rect 266358 59327 266414 59336
rect 262864 58472 262916 58478
rect 262864 58414 262916 58420
rect 269776 57866 269804 396238
rect 270512 240825 270540 396743
rect 270590 396672 270646 396681
rect 270590 396607 270646 396616
rect 270604 260574 270632 396607
rect 272352 396370 272380 397287
rect 273350 396808 273406 396817
rect 273350 396743 273406 396752
rect 273626 396808 273682 396817
rect 273626 396743 273682 396752
rect 276110 396808 276166 396817
rect 276110 396743 276166 396752
rect 277490 396808 277546 396817
rect 277490 396743 277546 396752
rect 272340 396364 272392 396370
rect 272340 396306 272392 396312
rect 273364 264450 273392 396743
rect 273640 396710 273668 396743
rect 273628 396704 273680 396710
rect 273442 396672 273498 396681
rect 273628 396646 273680 396652
rect 276018 396672 276074 396681
rect 273442 396607 273498 396616
rect 276018 396607 276074 396616
rect 273352 264444 273404 264450
rect 273352 264386 273404 264392
rect 273456 261322 273484 396607
rect 273444 261316 273496 261322
rect 273444 261258 273496 261264
rect 270592 260568 270644 260574
rect 270592 260510 270644 260516
rect 270498 240816 270554 240825
rect 270498 240751 270554 240760
rect 271142 227760 271198 227769
rect 271142 227695 271198 227704
rect 271156 193186 271184 227695
rect 271144 193180 271196 193186
rect 271144 193122 271196 193128
rect 276032 59430 276060 396607
rect 276124 264382 276152 396743
rect 277504 392630 277532 396743
rect 277688 396234 277716 397287
rect 277676 396228 277728 396234
rect 277676 396170 277728 396176
rect 278884 395486 278912 397287
rect 280158 396808 280214 396817
rect 283746 396808 283802 396817
rect 280158 396743 280214 396752
rect 282184 396772 282236 396778
rect 278872 395480 278924 395486
rect 278872 395422 278924 395428
rect 277492 392624 277544 392630
rect 277492 392566 277544 392572
rect 276112 264376 276164 264382
rect 276112 264318 276164 264324
rect 280172 262138 280200 396743
rect 283746 396743 283748 396752
rect 282184 396714 282236 396720
rect 283800 396743 283802 396752
rect 285954 396808 286010 396817
rect 285954 396743 286010 396752
rect 287058 396808 287114 396817
rect 287058 396743 287114 396752
rect 283748 396714 283800 396720
rect 280160 262132 280212 262138
rect 280160 262074 280212 262080
rect 282196 261390 282224 396714
rect 285968 396710 285996 396743
rect 284944 396704 284996 396710
rect 284944 396646 284996 396652
rect 285956 396704 286008 396710
rect 285956 396646 286008 396652
rect 284956 261458 284984 396646
rect 287072 373318 287100 396743
rect 290200 395418 290228 397287
rect 292670 396808 292726 396817
rect 291844 396772 291896 396778
rect 292670 396743 292672 396752
rect 291844 396714 291896 396720
rect 292724 396743 292726 396752
rect 295338 396808 295394 396817
rect 295338 396743 295394 396752
rect 292672 396714 292724 396720
rect 290188 395412 290240 395418
rect 290188 395354 290240 395360
rect 287060 373312 287112 373318
rect 287060 373254 287112 373260
rect 291856 262750 291884 396714
rect 291844 262744 291896 262750
rect 291844 262686 291896 262692
rect 284944 261452 284996 261458
rect 284944 261394 284996 261400
rect 282184 261384 282236 261390
rect 282184 261326 282236 261332
rect 295352 260506 295380 396743
rect 298480 395350 298508 397287
rect 298468 395344 298520 395350
rect 298468 395286 298520 395292
rect 295340 260500 295392 260506
rect 295340 260442 295392 260448
rect 276020 59424 276072 59430
rect 276020 59366 276072 59372
rect 300136 57934 300164 398103
rect 308586 397352 308642 397361
rect 304264 397316 304316 397322
rect 308586 397287 308588 397296
rect 304264 397258 304316 397264
rect 308640 397287 308642 397296
rect 308588 397258 308640 397264
rect 302238 396808 302294 396817
rect 302238 396743 302294 396752
rect 302252 59906 302280 396743
rect 304276 262206 304304 397258
rect 304998 396808 305054 396817
rect 304998 396743 305054 396752
rect 310518 396808 310574 396817
rect 310518 396743 310574 396752
rect 313278 396808 313334 396817
rect 313278 396743 313334 396752
rect 304264 262200 304316 262206
rect 304264 262142 304316 262148
rect 305012 260642 305040 396743
rect 310532 263566 310560 396743
rect 313292 265810 313320 396743
rect 315776 396302 315804 398103
rect 317418 396808 317474 396817
rect 317418 396743 317474 396752
rect 320178 396808 320234 396817
rect 320178 396743 320234 396752
rect 322938 396808 322994 396817
rect 322938 396743 322994 396752
rect 315764 396296 315816 396302
rect 315764 396238 315816 396244
rect 316684 396160 316736 396166
rect 316684 396102 316736 396108
rect 313280 265804 313332 265810
rect 313280 265746 313332 265752
rect 310520 263560 310572 263566
rect 310520 263502 310572 263508
rect 305000 260636 305052 260642
rect 305000 260578 305052 260584
rect 302240 59900 302292 59906
rect 302240 59842 302292 59848
rect 316696 58138 316724 396102
rect 317432 265742 317460 396743
rect 317420 265736 317472 265742
rect 317420 265678 317472 265684
rect 320192 236609 320220 396743
rect 320178 236600 320234 236609
rect 320178 236535 320234 236544
rect 322952 235249 322980 396743
rect 325896 396438 325924 398103
rect 342626 397352 342682 397361
rect 342626 397287 342682 397296
rect 342350 396808 342406 396817
rect 342350 396743 342406 396752
rect 325884 396432 325936 396438
rect 325884 396374 325936 396380
rect 322938 235240 322994 235249
rect 322938 235175 322994 235184
rect 342364 58342 342392 396743
rect 342640 396166 342668 397287
rect 342628 396160 342680 396166
rect 342628 396102 342680 396108
rect 356532 77217 356560 484463
rect 357438 418840 357494 418849
rect 357438 418775 357494 418784
rect 356518 77208 356574 77217
rect 356518 77143 356574 77152
rect 357452 58993 357480 418775
rect 357530 414352 357586 414361
rect 357530 414287 357586 414296
rect 357544 243545 357572 414287
rect 358096 260370 358124 563042
rect 359002 478952 359058 478961
rect 359002 478887 359058 478896
rect 358818 415848 358874 415857
rect 358818 415783 358874 415792
rect 358084 260364 358136 260370
rect 358084 260306 358136 260312
rect 357530 243536 357586 243545
rect 357530 243471 357586 243480
rect 358832 59129 358860 415783
rect 358910 413128 358966 413137
rect 358910 413063 358966 413072
rect 358924 265946 358952 413063
rect 359016 399566 359044 478887
rect 359094 417208 359150 417217
rect 359094 417143 359150 417152
rect 359004 399560 359056 399566
rect 359004 399502 359056 399508
rect 359108 399498 359136 417143
rect 359096 399492 359148 399498
rect 359096 399434 359148 399440
rect 358912 265940 358964 265946
rect 358912 265882 358964 265888
rect 360856 260302 360884 616830
rect 363616 260438 363644 670686
rect 367756 262002 367784 700266
rect 367744 261996 367796 262002
rect 367744 261938 367796 261944
rect 370516 261934 370544 700402
rect 381544 700392 381596 700398
rect 381544 700334 381596 700340
rect 378784 696992 378836 696998
rect 378784 696934 378836 696940
rect 377404 643136 377456 643142
rect 377404 643078 377456 643084
rect 376024 536852 376076 536858
rect 376024 536794 376076 536800
rect 374644 484424 374696 484430
rect 374644 484366 374696 484372
rect 371884 404388 371936 404394
rect 371884 404330 371936 404336
rect 370504 261928 370556 261934
rect 370504 261870 370556 261876
rect 363604 260432 363656 260438
rect 363604 260374 363656 260380
rect 360844 260296 360896 260302
rect 360844 260238 360896 260244
rect 371896 260234 371924 404330
rect 374656 261730 374684 484366
rect 376036 261798 376064 536794
rect 377416 263294 377444 643078
rect 377404 263288 377456 263294
rect 377404 263230 377456 263236
rect 378796 261866 378824 696934
rect 381556 263362 381584 700334
rect 382936 263430 382964 700470
rect 385696 263498 385724 700538
rect 396724 683188 396776 683194
rect 396724 683130 396776 683136
rect 395344 630692 395396 630698
rect 395344 630634 395396 630640
rect 393964 576904 394016 576910
rect 393964 576846 394016 576852
rect 392584 524476 392636 524482
rect 392584 524418 392636 524424
rect 389824 470620 389876 470626
rect 389824 470562 389876 470568
rect 388444 430636 388496 430642
rect 388444 430578 388496 430584
rect 385684 263492 385736 263498
rect 385684 263434 385736 263440
rect 382924 263424 382976 263430
rect 382924 263366 382976 263372
rect 381544 263356 381596 263362
rect 381544 263298 381596 263304
rect 388456 262954 388484 430578
rect 389836 263090 389864 470562
rect 389824 263084 389876 263090
rect 389824 263026 389876 263032
rect 392596 263022 392624 524418
rect 392584 263016 392636 263022
rect 392584 262958 392636 262964
rect 388444 262948 388496 262954
rect 388444 262890 388496 262896
rect 378784 261860 378836 261866
rect 378784 261802 378836 261808
rect 376024 261792 376076 261798
rect 376024 261734 376076 261740
rect 374644 261724 374696 261730
rect 374644 261666 374696 261672
rect 393976 261662 394004 576846
rect 395356 263158 395384 630634
rect 396736 263226 396764 683130
rect 399496 264314 399524 700538
rect 399484 264308 399536 264314
rect 399484 264250 399536 264256
rect 396724 263220 396776 263226
rect 396724 263162 396776 263168
rect 395344 263152 395396 263158
rect 395344 263094 395396 263100
rect 412652 262886 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 425704 456816 425756 456822
rect 425704 456758 425756 456764
rect 412640 262880 412692 262886
rect 412640 262822 412692 262828
rect 393964 261656 394016 261662
rect 393964 261598 394016 261604
rect 371884 260228 371936 260234
rect 371884 260170 371936 260176
rect 425716 260166 425744 456758
rect 429212 261594 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700534 462360 703520
rect 478524 700602 478552 703520
rect 478512 700596 478564 700602
rect 478512 700538 478564 700544
rect 462320 700528 462372 700534
rect 462320 700470 462372 700476
rect 494808 700466 494836 703520
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 527192 700398 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 542372 264246 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 558184 590708 558236 590714
rect 558184 590650 558236 590656
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 542360 264240 542412 264246
rect 542360 264182 542412 264188
rect 429200 261588 429252 261594
rect 429200 261530 429252 261536
rect 558196 261526 558224 590650
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580262 418296 580318 418305
rect 580262 418231 580318 418240
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579618 365120 579674 365129
rect 579618 365055 579674 365064
rect 579632 364410 579660 365055
rect 579620 364404 579672 364410
rect 579620 364346 579672 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 580276 265674 580304 418231
rect 580264 265668 580316 265674
rect 580264 265610 580316 265616
rect 558184 261520 558236 261526
rect 558184 261462 558236 261468
rect 425704 260160 425756 260166
rect 425704 260102 425756 260108
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 580262 230616 580318 230625
rect 580262 230551 580318 230560
rect 410522 226400 410578 226409
rect 410522 226335 410578 226344
rect 410536 100706 410564 226335
rect 580172 193180 580224 193186
rect 580172 193122 580224 193128
rect 580184 192545 580212 193122
rect 580170 192536 580226 192545
rect 580170 192471 580226 192480
rect 410524 100700 410576 100706
rect 410524 100642 410576 100648
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 59968 580224 59974
rect 580172 59910 580224 59916
rect 580184 59673 580212 59910
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 358818 59120 358874 59129
rect 358818 59055 358874 59064
rect 357438 58984 357494 58993
rect 357438 58919 357494 58928
rect 342352 58336 342404 58342
rect 342352 58278 342404 58284
rect 316684 58132 316736 58138
rect 316684 58074 316736 58080
rect 300124 57928 300176 57934
rect 300124 57870 300176 57876
rect 269764 57860 269816 57866
rect 269764 57802 269816 57808
rect 347136 57656 347188 57662
rect 347136 57598 347188 57604
rect 347044 57588 347096 57594
rect 347044 57530 347096 57536
rect 258724 56976 258776 56982
rect 251822 56944 251878 56953
rect 258724 56918 258776 56924
rect 251822 56879 251878 56888
rect 271144 56772 271196 56778
rect 271144 56714 271196 56720
rect 258080 53032 258132 53038
rect 258080 52974 258132 52980
rect 253940 52964 253992 52970
rect 253940 52906 253992 52912
rect 251180 52828 251232 52834
rect 251180 52770 251232 52776
rect 240140 52760 240192 52766
rect 240140 52702 240192 52708
rect 238116 33108 238168 33114
rect 238116 33050 238168 33056
rect 234068 20664 234120 20670
rect 234068 20606 234120 20612
rect 236000 18692 236052 18698
rect 236000 18634 236052 18640
rect 236012 16574 236040 18634
rect 238116 16584 238168 16590
rect 224972 16546 225184 16574
rect 227732 16546 228772 16574
rect 231872 16546 232268 16574
rect 233252 16546 233464 16574
rect 236012 16546 237052 16574
rect 223948 15632 224000 15638
rect 223948 15574 224000 15580
rect 222752 10056 222804 10062
rect 222752 9998 222804 10004
rect 221648 3120 221700 3126
rect 221648 3062 221700 3068
rect 221556 2916 221608 2922
rect 221556 2858 221608 2864
rect 221384 2774 221596 2802
rect 221568 480 221596 2774
rect 222764 480 222792 9998
rect 223960 480 223988 15574
rect 225156 480 225184 16546
rect 227536 15700 227588 15706
rect 227536 15642 227588 15648
rect 226432 10124 226484 10130
rect 226432 10066 226484 10072
rect 226444 3482 226472 10066
rect 226352 3454 226472 3482
rect 226352 480 226380 3454
rect 227548 480 227576 15642
rect 228744 480 228772 16546
rect 231032 15768 231084 15774
rect 231032 15710 231084 15716
rect 229836 10192 229888 10198
rect 229836 10134 229888 10140
rect 229848 480 229876 10134
rect 231044 480 231072 15710
rect 232240 480 232268 16546
rect 233436 480 233464 16546
rect 234620 15836 234672 15842
rect 234620 15778 234672 15784
rect 234632 480 234660 15778
rect 235816 5568 235868 5574
rect 235816 5510 235868 5516
rect 235828 480 235856 5510
rect 237024 480 237052 16546
rect 240152 16574 240180 52702
rect 247040 17196 247092 17202
rect 247040 17138 247092 17144
rect 242900 17060 242952 17066
rect 242900 17002 242952 17008
rect 240152 16546 240548 16574
rect 238116 16526 238168 16532
rect 238128 480 238156 16526
rect 239312 5636 239364 5642
rect 239312 5578 239364 5584
rect 239324 480 239352 5578
rect 240520 480 240548 16546
rect 241704 16516 241756 16522
rect 241704 16458 241756 16464
rect 241716 480 241744 16458
rect 242912 2854 242940 17002
rect 247052 16574 247080 17138
rect 247052 16546 247632 16574
rect 245200 16448 245252 16454
rect 245200 16390 245252 16396
rect 242992 5704 243044 5710
rect 242992 5646 243044 5652
rect 242900 2848 242952 2854
rect 242900 2790 242952 2796
rect 243004 2666 243032 5646
rect 244096 2848 244148 2854
rect 244096 2790 244148 2796
rect 242912 2638 243032 2666
rect 242912 480 242940 2638
rect 244108 480 244136 2790
rect 245212 480 245240 16390
rect 246396 5772 246448 5778
rect 246396 5714 246448 5720
rect 246408 480 246436 5714
rect 247604 480 247632 16546
rect 248788 16380 248840 16386
rect 248788 16322 248840 16328
rect 248800 480 248828 16322
rect 249984 5840 250036 5846
rect 249984 5782 250036 5788
rect 249996 480 250024 5782
rect 251192 480 251220 52770
rect 253952 16574 253980 52906
rect 258092 16574 258120 52974
rect 260840 17944 260892 17950
rect 260840 17886 260892 17892
rect 260852 16574 260880 17886
rect 269120 17876 269172 17882
rect 269120 17818 269172 17824
rect 269132 16574 269160 17818
rect 253952 16546 254716 16574
rect 258092 16546 258304 16574
rect 260852 16546 261800 16574
rect 269132 16546 270080 16574
rect 252376 16312 252428 16318
rect 252376 16254 252428 16260
rect 252388 480 252416 16254
rect 253480 5908 253532 5914
rect 253480 5850 253532 5856
rect 253492 480 253520 5850
rect 254688 480 254716 16546
rect 255872 16244 255924 16250
rect 255872 16186 255924 16192
rect 255884 480 255912 16186
rect 257068 5976 257120 5982
rect 257068 5918 257120 5924
rect 257080 480 257108 5918
rect 258276 480 258304 16546
rect 259460 16176 259512 16182
rect 259460 16118 259512 16124
rect 259472 480 259500 16118
rect 260656 6044 260708 6050
rect 260656 5986 260708 5992
rect 260668 480 260696 5986
rect 261772 480 261800 16546
rect 262956 16108 263008 16114
rect 262956 16050 263008 16056
rect 262968 480 262996 16050
rect 266544 16040 266596 16046
rect 266544 15982 266596 15988
rect 265348 11144 265400 11150
rect 265348 11086 265400 11092
rect 264152 6112 264204 6118
rect 264152 6054 264204 6060
rect 264164 480 264192 6054
rect 265360 480 265388 11086
rect 266556 480 266584 15982
rect 268844 11212 268896 11218
rect 268844 11154 268896 11160
rect 267740 6860 267792 6866
rect 267740 6802 267792 6808
rect 267752 480 267780 6802
rect 268856 480 268884 11154
rect 270052 480 270080 16546
rect 270408 6792 270460 6798
rect 270408 6734 270460 6740
rect 270420 2854 270448 6734
rect 271156 6118 271184 56714
rect 313280 55820 313332 55826
rect 313280 55762 313332 55768
rect 309140 54324 309192 54330
rect 309140 54266 309192 54272
rect 302240 54256 302292 54262
rect 302240 54198 302292 54204
rect 291200 50312 291252 50318
rect 291200 50254 291252 50260
rect 273260 17808 273312 17814
rect 273260 17750 273312 17756
rect 273272 16574 273300 17750
rect 276020 17740 276072 17746
rect 276020 17682 276072 17688
rect 273272 16546 273668 16574
rect 271236 6180 271288 6186
rect 271236 6122 271288 6128
rect 271144 6112 271196 6118
rect 271144 6054 271196 6060
rect 270408 2848 270460 2854
rect 270408 2790 270460 2796
rect 271248 480 271276 6122
rect 272432 2848 272484 2854
rect 272432 2790 272484 2796
rect 272444 480 272472 2790
rect 273640 480 273668 16546
rect 274824 6724 274876 6730
rect 274824 6666 274876 6672
rect 274836 480 274864 6666
rect 276032 4214 276060 17682
rect 280160 17672 280212 17678
rect 280160 17614 280212 17620
rect 280172 16574 280200 17614
rect 284300 17604 284352 17610
rect 284300 17546 284352 17552
rect 280172 16546 280752 16574
rect 279516 11348 279568 11354
rect 279516 11290 279568 11296
rect 276112 11280 276164 11286
rect 276112 11222 276164 11228
rect 276020 4208 276072 4214
rect 276020 4150 276072 4156
rect 276124 3482 276152 11222
rect 278320 6656 278372 6662
rect 278320 6598 278372 6604
rect 277124 4208 277176 4214
rect 277124 4150 277176 4156
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 277136 480 277164 4150
rect 278332 480 278360 6598
rect 279528 480 279556 11290
rect 280724 480 280752 16546
rect 281908 6588 281960 6594
rect 281908 6530 281960 6536
rect 281920 480 281948 6530
rect 283104 3188 283156 3194
rect 283104 3130 283156 3136
rect 283116 480 283144 3130
rect 284312 480 284340 17546
rect 287060 17536 287112 17542
rect 287060 17478 287112 17484
rect 287072 16574 287100 17478
rect 291212 16574 291240 50254
rect 300860 17332 300912 17338
rect 300860 17274 300912 17280
rect 300872 16574 300900 17274
rect 302252 16574 302280 54198
rect 309152 16574 309180 54266
rect 311900 51060 311952 51066
rect 311900 51002 311952 51008
rect 311912 16574 311940 51002
rect 313292 16574 313320 55762
rect 324320 55208 324372 55214
rect 324320 55150 324372 55156
rect 320180 54460 320232 54466
rect 320180 54402 320232 54408
rect 316040 54392 316092 54398
rect 316040 54334 316092 54340
rect 287072 16546 287836 16574
rect 291212 16546 291424 16574
rect 300872 16546 302004 16574
rect 302252 16546 303200 16574
rect 309152 16546 310284 16574
rect 311912 16546 312676 16574
rect 313292 16546 313872 16574
rect 286600 11416 286652 11422
rect 286600 11358 286652 11364
rect 285404 6520 285456 6526
rect 285404 6462 285456 6468
rect 285416 480 285444 6462
rect 286612 480 286640 11358
rect 287808 480 287836 16546
rect 290188 11484 290240 11490
rect 290188 11426 290240 11432
rect 288992 6452 289044 6458
rect 288992 6394 289044 6400
rect 289004 480 289032 6394
rect 290200 480 290228 11426
rect 291396 480 291424 16546
rect 299480 11688 299532 11694
rect 299480 11630 299532 11636
rect 297272 11620 297324 11626
rect 297272 11562 297324 11568
rect 293684 11552 293736 11558
rect 293684 11494 293736 11500
rect 292580 6384 292632 6390
rect 292580 6326 292632 6332
rect 292592 480 292620 6326
rect 293696 480 293724 11494
rect 296076 6316 296128 6322
rect 296076 6258 296128 6264
rect 294880 3324 294932 3330
rect 294880 3266 294932 3272
rect 294892 480 294920 3266
rect 296088 480 296116 6258
rect 297284 480 297312 11562
rect 299492 3330 299520 11630
rect 299664 6248 299716 6254
rect 299664 6190 299716 6196
rect 299480 3324 299532 3330
rect 299480 3266 299532 3272
rect 298468 2916 298520 2922
rect 298468 2858 298520 2864
rect 298480 480 298508 2858
rect 299676 480 299704 6190
rect 300768 3324 300820 3330
rect 300768 3266 300820 3272
rect 300780 480 300808 3266
rect 301976 480 302004 16546
rect 303172 480 303200 16546
rect 304356 12436 304408 12442
rect 304356 12378 304408 12384
rect 304368 480 304396 12378
rect 307944 12368 307996 12374
rect 307944 12310 307996 12316
rect 306748 3392 306800 3398
rect 306748 3334 306800 3340
rect 305552 2984 305604 2990
rect 305552 2926 305604 2932
rect 305564 480 305592 2926
rect 306760 480 306788 3334
rect 307956 480 307984 12310
rect 309048 4140 309100 4146
rect 309048 4082 309100 4088
rect 309060 480 309088 4082
rect 310256 480 310284 16546
rect 311440 12300 311492 12306
rect 311440 12242 311492 12248
rect 311452 480 311480 12242
rect 312648 480 312676 16546
rect 313844 480 313872 16546
rect 315028 12232 315080 12238
rect 315028 12174 315080 12180
rect 315040 480 315068 12174
rect 316052 3398 316080 54334
rect 316132 49156 316184 49162
rect 316132 49098 316184 49104
rect 316144 16574 316172 49098
rect 318800 17264 318852 17270
rect 318800 17206 318852 17212
rect 318812 16574 318840 17206
rect 320192 16574 320220 54402
rect 324332 16574 324360 55150
rect 327080 55140 327132 55146
rect 327080 55082 327132 55088
rect 325700 17400 325752 17406
rect 325700 17342 325752 17348
rect 325712 16574 325740 17342
rect 327092 16574 327120 55082
rect 331220 55072 331272 55078
rect 331220 55014 331272 55020
rect 329840 49088 329892 49094
rect 329840 49030 329892 49036
rect 329852 16574 329880 49030
rect 331232 16574 331260 55014
rect 335360 52420 335412 52426
rect 335360 52362 335412 52368
rect 335372 16574 335400 52362
rect 339500 52352 339552 52358
rect 339500 52294 339552 52300
rect 336740 17468 336792 17474
rect 336740 17410 336792 17416
rect 336752 16574 336780 17410
rect 339512 16574 339540 52294
rect 342260 52284 342312 52290
rect 342260 52226 342312 52232
rect 340880 49020 340932 49026
rect 340880 48962 340932 48968
rect 340892 16574 340920 48962
rect 342272 16574 342300 52226
rect 346400 52216 346452 52222
rect 346400 52158 346452 52164
rect 346412 16574 346440 52158
rect 316144 16546 316264 16574
rect 318812 16546 319760 16574
rect 320192 16546 320956 16574
rect 324332 16546 324452 16574
rect 325712 16546 326844 16574
rect 327092 16546 328040 16574
rect 329852 16546 330432 16574
rect 331232 16546 331628 16574
rect 335372 16546 336320 16574
rect 336752 16546 337516 16574
rect 339512 16546 339908 16574
rect 340892 16546 341012 16574
rect 342272 16546 343404 16574
rect 346412 16546 346992 16574
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 316236 480 316264 16546
rect 318524 12164 318576 12170
rect 318524 12106 318576 12112
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 318536 480 318564 12106
rect 319732 480 319760 16546
rect 320928 480 320956 16546
rect 322112 12096 322164 12102
rect 322112 12038 322164 12044
rect 322124 480 322152 12038
rect 323308 3052 323360 3058
rect 323308 2994 323360 3000
rect 323320 480 323348 2994
rect 324424 480 324452 16546
rect 325608 12028 325660 12034
rect 325608 11970 325660 11976
rect 325620 480 325648 11970
rect 326816 480 326844 16546
rect 328012 480 328040 16546
rect 329196 11960 329248 11966
rect 329196 11902 329248 11908
rect 329208 480 329236 11902
rect 330404 480 330432 16546
rect 331600 480 331628 16546
rect 332692 11892 332744 11898
rect 332692 11834 332744 11840
rect 332704 480 332732 11834
rect 335084 7064 335136 7070
rect 335084 7006 335136 7012
rect 333888 4072 333940 4078
rect 333888 4014 333940 4020
rect 333900 480 333928 4014
rect 335096 480 335124 7006
rect 336292 480 336320 16546
rect 337488 480 337516 16546
rect 338672 7132 338724 7138
rect 338672 7074 338724 7080
rect 338684 480 338712 7074
rect 339880 480 339908 16546
rect 340984 480 341012 16546
rect 342168 7200 342220 7206
rect 342168 7142 342220 7148
rect 342180 480 342208 7142
rect 343376 480 343404 16546
rect 345756 7268 345808 7274
rect 345756 7210 345808 7216
rect 344560 3936 344612 3942
rect 344560 3878 344612 3884
rect 344572 480 344600 3878
rect 345768 480 345796 7210
rect 346964 480 346992 16546
rect 347056 3398 347084 57530
rect 347044 3392 347096 3398
rect 347044 3334 347096 3340
rect 347148 3330 347176 57598
rect 353300 57520 353352 57526
rect 353300 57462 353352 57468
rect 347780 19984 347832 19990
rect 347780 19926 347832 19932
rect 347792 16574 347820 19926
rect 353312 16574 353340 57462
rect 411904 57452 411956 57458
rect 411904 57394 411956 57400
rect 407764 56568 407816 56574
rect 407764 56510 407816 56516
rect 405740 55004 405792 55010
rect 405740 54946 405792 54952
rect 367100 53780 367152 53786
rect 367100 53722 367152 53728
rect 357440 52148 357492 52154
rect 357440 52090 357492 52096
rect 357452 16574 357480 52090
rect 360200 52080 360252 52086
rect 360200 52022 360252 52028
rect 360212 16574 360240 52022
rect 364340 52012 364392 52018
rect 364340 51954 364392 51960
rect 364352 16574 364380 51954
rect 367112 16574 367140 53722
rect 405752 16574 405780 54946
rect 347792 16546 348096 16574
rect 353312 16546 354076 16574
rect 357452 16546 357572 16574
rect 360212 16546 361160 16574
rect 364352 16546 364656 16574
rect 367112 16546 368244 16574
rect 405752 16546 406056 16574
rect 347136 3324 347188 3330
rect 347136 3266 347188 3272
rect 348068 480 348096 16546
rect 352840 7336 352892 7342
rect 352840 7278 352892 7284
rect 351644 3868 351696 3874
rect 351644 3810 351696 3816
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 349264 480 349292 3334
rect 350448 3324 350500 3330
rect 350448 3266 350500 3272
rect 350460 480 350488 3266
rect 351656 480 351684 3810
rect 352852 480 352880 7278
rect 354048 480 354076 16546
rect 356336 7404 356388 7410
rect 356336 7346 356388 7352
rect 355232 3800 355284 3806
rect 355232 3742 355284 3748
rect 355244 480 355272 3742
rect 356348 480 356376 7346
rect 357544 480 357572 16546
rect 359924 7472 359976 7478
rect 359924 7414 359976 7420
rect 358726 6896 358782 6905
rect 358726 6831 358782 6840
rect 358740 480 358768 6831
rect 359936 480 359964 7414
rect 361132 480 361160 16546
rect 363512 7540 363564 7546
rect 363512 7482 363564 7488
rect 362314 6760 362370 6769
rect 362314 6695 362370 6704
rect 362328 480 362356 6695
rect 363524 480 363552 7482
rect 364628 480 364656 16546
rect 367008 8288 367060 8294
rect 367008 8230 367060 8236
rect 365810 6624 365866 6633
rect 365810 6559 365866 6568
rect 365824 480 365852 6559
rect 367020 480 367048 8230
rect 368216 480 368244 16546
rect 403624 13796 403676 13802
rect 403624 13738 403676 13744
rect 398840 13048 398892 13054
rect 398840 12990 398892 12996
rect 396540 12980 396592 12986
rect 396540 12922 396592 12928
rect 393044 12912 393096 12918
rect 393044 12854 393096 12860
rect 389456 12844 389508 12850
rect 389456 12786 389508 12792
rect 385960 12776 386012 12782
rect 385960 12718 386012 12724
rect 382372 12708 382424 12714
rect 382372 12650 382424 12656
rect 378876 12640 378928 12646
rect 378876 12582 378928 12588
rect 374000 12572 374052 12578
rect 374000 12514 374052 12520
rect 370596 8220 370648 8226
rect 370596 8162 370648 8168
rect 369400 2168 369452 2174
rect 369400 2110 369452 2116
rect 369412 480 369440 2110
rect 370608 480 370636 8162
rect 374012 3398 374040 12514
rect 374092 8152 374144 8158
rect 374092 8094 374144 8100
rect 374000 3392 374052 3398
rect 374000 3334 374052 3340
rect 371700 3120 371752 3126
rect 371700 3062 371752 3068
rect 371712 480 371740 3062
rect 372896 2100 372948 2106
rect 372896 2042 372948 2048
rect 372908 480 372936 2042
rect 374104 480 374132 8094
rect 377680 8084 377732 8090
rect 377680 8026 377732 8032
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 375300 480 375328 3334
rect 376484 3256 376536 3262
rect 376484 3198 376536 3204
rect 376496 480 376524 3198
rect 377692 480 377720 8026
rect 378888 480 378916 12582
rect 381176 8016 381228 8022
rect 381176 7958 381228 7964
rect 379978 6488 380034 6497
rect 379978 6423 380034 6432
rect 379992 480 380020 6423
rect 381188 480 381216 7958
rect 382384 480 382412 12650
rect 384764 7948 384816 7954
rect 384764 7890 384816 7896
rect 383566 6352 383622 6361
rect 383566 6287 383622 6296
rect 383580 480 383608 6287
rect 384776 480 384804 7890
rect 385972 480 386000 12718
rect 387156 8356 387208 8362
rect 387156 8298 387208 8304
rect 387168 480 387196 8298
rect 388260 7880 388312 7886
rect 388260 7822 388312 7828
rect 388272 480 388300 7822
rect 389468 480 389496 12786
rect 391848 7812 391900 7818
rect 391848 7754 391900 7760
rect 390650 6080 390706 6089
rect 390650 6015 390706 6024
rect 390664 480 390692 6015
rect 391860 480 391888 7754
rect 393056 480 393084 12854
rect 395344 7744 395396 7750
rect 395344 7686 395396 7692
rect 394240 3732 394292 3738
rect 394240 3674 394292 3680
rect 394252 480 394280 3674
rect 395356 480 395384 7686
rect 396552 480 396580 12922
rect 397736 3664 397788 3670
rect 397736 3606 397788 3612
rect 397748 480 397776 3606
rect 398852 3398 398880 12990
rect 401324 8424 401376 8430
rect 401324 8366 401376 8372
rect 398932 7676 398984 7682
rect 398932 7618 398984 7624
rect 398840 3392 398892 3398
rect 398840 3334 398892 3340
rect 398944 480 398972 7618
rect 400128 3392 400180 3398
rect 400128 3334 400180 3340
rect 400140 480 400168 3334
rect 401336 480 401364 8366
rect 402520 7608 402572 7614
rect 402520 7550 402572 7556
rect 402532 480 402560 7550
rect 403636 480 403664 13738
rect 404820 8492 404872 8498
rect 404820 8434 404872 8440
rect 404832 480 404860 8434
rect 406028 480 406056 16546
rect 407212 13728 407264 13734
rect 407212 13670 407264 13676
rect 407224 480 407252 13670
rect 407776 3398 407804 56510
rect 411916 16574 411944 57394
rect 418804 57384 418856 57390
rect 418804 57326 418856 57332
rect 412640 54936 412692 54942
rect 412640 54878 412692 54884
rect 412652 16574 412680 54878
rect 414664 54868 414716 54874
rect 414664 54810 414716 54816
rect 411916 16546 412036 16574
rect 412652 16546 413140 16574
rect 410800 13660 410852 13666
rect 410800 13602 410852 13608
rect 408408 4004 408460 4010
rect 408408 3946 408460 3952
rect 407764 3392 407816 3398
rect 407764 3334 407816 3340
rect 408420 480 408448 3946
rect 409604 3392 409656 3398
rect 409604 3334 409656 3340
rect 409616 480 409644 3334
rect 410812 480 410840 13602
rect 411902 6216 411958 6225
rect 411902 6151 411958 6160
rect 411916 480 411944 6151
rect 412008 3738 412036 16546
rect 411996 3732 412048 3738
rect 411996 3674 412048 3680
rect 413112 480 413140 16546
rect 414296 13592 414348 13598
rect 414296 13534 414348 13540
rect 414308 480 414336 13534
rect 414676 3466 414704 54810
rect 417424 54800 417476 54806
rect 417424 54742 417476 54748
rect 417436 16574 417464 54742
rect 417436 16546 417556 16574
rect 417424 13524 417476 13530
rect 417424 13466 417476 13472
rect 415492 3596 415544 3602
rect 415492 3538 415544 3544
rect 414664 3460 414716 3466
rect 414664 3402 414716 3408
rect 415504 480 415532 3538
rect 416688 3460 416740 3466
rect 416688 3402 416740 3408
rect 416700 480 416728 3402
rect 417436 2938 417464 13466
rect 417528 3058 417556 16546
rect 418816 3806 418844 57326
rect 425704 57316 425756 57322
rect 425704 57258 425756 57264
rect 421564 56500 421616 56506
rect 421564 56442 421616 56448
rect 421380 13456 421432 13462
rect 421380 13398 421432 13404
rect 418988 8560 419040 8566
rect 418988 8502 419040 8508
rect 418804 3800 418856 3806
rect 418804 3742 418856 3748
rect 417516 3052 417568 3058
rect 417516 2994 417568 3000
rect 417436 2910 417924 2938
rect 417896 480 417924 2910
rect 419000 480 419028 8502
rect 420184 3052 420236 3058
rect 420184 2994 420236 3000
rect 420196 480 420224 2994
rect 421392 480 421420 13398
rect 421576 4146 421604 56442
rect 423772 13388 423824 13394
rect 423772 13330 423824 13336
rect 422576 8628 422628 8634
rect 422576 8570 422628 8576
rect 421564 4140 421616 4146
rect 421564 4082 421616 4088
rect 422588 480 422616 8570
rect 423680 4140 423732 4146
rect 423680 4082 423732 4088
rect 423692 2122 423720 4082
rect 423784 3534 423812 13330
rect 425716 3874 425744 57258
rect 429844 57248 429896 57254
rect 429844 57190 429896 57196
rect 436742 57216 436798 57225
rect 425796 54732 425848 54738
rect 425796 54674 425848 54680
rect 425704 3868 425756 3874
rect 425704 3810 425756 3816
rect 425808 3534 425836 54674
rect 428464 13320 428516 13326
rect 428464 13262 428516 13268
rect 423772 3528 423824 3534
rect 423772 3470 423824 3476
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 425796 3528 425848 3534
rect 425796 3470 425848 3476
rect 427268 3528 427320 3534
rect 427268 3470 427320 3476
rect 423692 2094 423812 2122
rect 423784 480 423812 2094
rect 424980 480 425008 3470
rect 426164 3460 426216 3466
rect 426164 3402 426216 3408
rect 426176 480 426204 3402
rect 427280 480 427308 3470
rect 428476 480 428504 13262
rect 429856 3602 429884 57190
rect 436742 57151 436798 57160
rect 430580 53712 430632 53718
rect 430580 53654 430632 53660
rect 430592 16574 430620 53654
rect 432604 53644 432656 53650
rect 432604 53586 432656 53592
rect 430592 16546 430896 16574
rect 429844 3596 429896 3602
rect 429844 3538 429896 3544
rect 429660 3392 429712 3398
rect 429660 3334 429712 3340
rect 429672 480 429700 3334
rect 430868 480 430896 16546
rect 432052 13252 432104 13258
rect 432052 13194 432104 13200
rect 432064 480 432092 13194
rect 432616 3466 432644 53586
rect 436756 16574 436784 57151
rect 443644 56432 443696 56438
rect 443644 56374 443696 56380
rect 439504 54664 439556 54670
rect 439504 54606 439556 54612
rect 436756 16546 436876 16574
rect 435548 13184 435600 13190
rect 435548 13126 435600 13132
rect 432604 3460 432656 3466
rect 432604 3402 432656 3408
rect 434444 3460 434496 3466
rect 434444 3402 434496 3408
rect 433246 3224 433302 3233
rect 433246 3159 433302 3168
rect 433260 480 433288 3159
rect 434456 480 434484 3402
rect 435560 480 435588 13126
rect 436742 4040 436798 4049
rect 436742 3975 436798 3984
rect 436756 480 436784 3975
rect 436848 3466 436876 16546
rect 439136 13116 439188 13122
rect 439136 13058 439188 13064
rect 437940 8696 437992 8702
rect 437940 8638 437992 8644
rect 436836 3460 436888 3466
rect 436836 3402 436888 3408
rect 437952 480 437980 8638
rect 439148 480 439176 13058
rect 439516 4146 439544 54606
rect 440240 18624 440292 18630
rect 440240 18566 440292 18572
rect 440252 16574 440280 18566
rect 440252 16546 440372 16574
rect 439504 4140 439556 4146
rect 439504 4082 439556 4088
rect 440344 480 440372 16546
rect 441528 8764 441580 8770
rect 441528 8706 441580 8712
rect 441540 480 441568 8706
rect 442632 4140 442684 4146
rect 442632 4082 442684 4088
rect 442644 480 442672 4082
rect 443656 3670 443684 56374
rect 450544 56364 450596 56370
rect 450544 56306 450596 56312
rect 447784 56296 447836 56302
rect 447784 56238 447836 56244
rect 445760 51944 445812 51950
rect 445760 51886 445812 51892
rect 445772 16574 445800 51886
rect 445772 16546 446260 16574
rect 443828 8900 443880 8906
rect 443828 8842 443880 8848
rect 443644 3664 443696 3670
rect 443644 3606 443696 3612
rect 443840 480 443868 8842
rect 445024 8832 445076 8838
rect 445024 8774 445076 8780
rect 445036 480 445064 8774
rect 446232 480 446260 16546
rect 447416 6180 447468 6186
rect 447416 6122 447468 6128
rect 447428 480 447456 6122
rect 447796 3942 447824 56238
rect 448520 51876 448572 51882
rect 448520 51818 448572 51824
rect 447784 3936 447836 3942
rect 447784 3878 447836 3884
rect 448532 3602 448560 51818
rect 450452 11824 450504 11830
rect 450452 11766 450504 11772
rect 448612 9648 448664 9654
rect 448612 9590 448664 9596
rect 448520 3596 448572 3602
rect 448520 3538 448572 3544
rect 448624 480 448652 9590
rect 449808 3596 449860 3602
rect 449808 3538 449860 3544
rect 449820 480 449848 3538
rect 450464 3482 450492 11766
rect 450556 3670 450584 56306
rect 454684 56228 454736 56234
rect 454684 56170 454736 56176
rect 452660 50992 452712 50998
rect 452660 50934 452712 50940
rect 452672 16574 452700 50934
rect 452672 16546 453344 16574
rect 452108 9580 452160 9586
rect 452108 9522 452160 9528
rect 450544 3664 450596 3670
rect 450544 3606 450596 3612
rect 450464 3454 450952 3482
rect 450924 480 450952 3454
rect 452120 480 452148 9522
rect 453316 480 453344 16546
rect 454696 3738 454724 56170
rect 461584 56160 461636 56166
rect 461584 56102 461636 56108
rect 456800 53508 456852 53514
rect 456800 53450 456852 53456
rect 456812 16574 456840 53450
rect 459560 51808 459612 51814
rect 459560 51750 459612 51756
rect 459572 16574 459600 51750
rect 461596 16574 461624 56102
rect 472624 56092 472676 56098
rect 472624 56034 472676 56040
rect 468484 53576 468536 53582
rect 468484 53518 468536 53524
rect 463700 50924 463752 50930
rect 463700 50866 463752 50872
rect 463712 16574 463740 50866
rect 466460 50856 466512 50862
rect 466460 50798 466512 50804
rect 466472 16574 466500 50798
rect 456812 16546 456932 16574
rect 459572 16546 460428 16574
rect 461596 16546 461716 16574
rect 463712 16546 464016 16574
rect 466472 16546 467512 16574
rect 455696 9512 455748 9518
rect 455696 9454 455748 9460
rect 454500 3732 454552 3738
rect 454500 3674 454552 3680
rect 454684 3732 454736 3738
rect 454684 3674 454736 3680
rect 454512 480 454540 3674
rect 455708 480 455736 9454
rect 456904 480 456932 16546
rect 459192 9444 459244 9450
rect 459192 9386 459244 9392
rect 458086 3904 458142 3913
rect 458086 3839 458142 3848
rect 458100 480 458128 3839
rect 459204 480 459232 9386
rect 460400 480 460428 16546
rect 461688 3806 461716 16546
rect 462780 9376 462832 9382
rect 462780 9318 462832 9324
rect 461584 3800 461636 3806
rect 461584 3742 461636 3748
rect 461676 3800 461728 3806
rect 461676 3742 461728 3748
rect 461596 480 461624 3742
rect 462792 480 462820 9318
rect 463988 480 464016 16546
rect 465172 11756 465224 11762
rect 465172 11698 465224 11704
rect 465184 480 465212 11698
rect 466276 9308 466328 9314
rect 466276 9250 466328 9256
rect 466288 480 466316 9250
rect 467484 480 467512 16546
rect 468496 4010 468524 53518
rect 470600 50788 470652 50794
rect 470600 50730 470652 50736
rect 470612 16574 470640 50730
rect 470612 16546 471100 16574
rect 469864 9240 469916 9246
rect 469864 9182 469916 9188
rect 468484 4004 468536 4010
rect 468484 3946 468536 3952
rect 468668 3868 468720 3874
rect 468668 3810 468720 3816
rect 468680 480 468708 3810
rect 469876 480 469904 9182
rect 471072 480 471100 16546
rect 472636 4146 472664 56034
rect 500960 56024 501012 56030
rect 500960 55966 501012 55972
rect 475384 54596 475436 54602
rect 475384 54538 475436 54544
rect 473360 13932 473412 13938
rect 473360 13874 473412 13880
rect 472624 4140 472676 4146
rect 472624 4082 472676 4088
rect 472254 3768 472310 3777
rect 472254 3703 472310 3712
rect 472268 480 472296 3703
rect 473372 3534 473400 13874
rect 473452 9172 473504 9178
rect 473452 9114 473504 9120
rect 473360 3528 473412 3534
rect 473360 3470 473412 3476
rect 473464 480 473492 9114
rect 475396 3874 475424 54538
rect 479524 53440 479576 53446
rect 479524 53382 479576 53388
rect 478144 14000 478196 14006
rect 478144 13942 478196 13948
rect 476948 9104 477000 9110
rect 476948 9046 477000 9052
rect 475384 3868 475436 3874
rect 475384 3810 475436 3816
rect 474556 3528 474608 3534
rect 474556 3470 474608 3476
rect 474568 480 474596 3470
rect 475752 3392 475804 3398
rect 475752 3334 475804 3340
rect 475764 480 475792 3334
rect 476960 480 476988 9046
rect 478156 480 478184 13942
rect 479536 4078 479564 53382
rect 483664 53372 483716 53378
rect 483664 53314 483716 53320
rect 481640 14068 481692 14074
rect 481640 14010 481692 14016
rect 479524 4072 479576 4078
rect 479524 4014 479576 4020
rect 479338 3632 479394 3641
rect 479338 3567 479394 3576
rect 479352 480 479380 3567
rect 481652 3534 481680 14010
rect 481730 9480 481786 9489
rect 481730 9415 481786 9424
rect 481640 3528 481692 3534
rect 480534 3496 480590 3505
rect 481640 3470 481692 3476
rect 480534 3431 480590 3440
rect 480548 480 480576 3431
rect 481744 480 481772 9415
rect 483676 3534 483704 53314
rect 500972 16574 501000 55966
rect 507860 55956 507912 55962
rect 507860 55898 507912 55904
rect 507872 16574 507900 55898
rect 564440 55888 564492 55894
rect 564440 55830 564492 55836
rect 544384 54528 544436 54534
rect 544384 54470 544436 54476
rect 512644 53304 512696 53310
rect 512644 53246 512696 53252
rect 500972 16546 501828 16574
rect 507872 16546 508912 16574
rect 500592 14408 500644 14414
rect 500592 14350 500644 14356
rect 497096 14340 497148 14346
rect 497096 14282 497148 14288
rect 493508 14272 493560 14278
rect 493508 14214 493560 14220
rect 489920 14204 489972 14210
rect 489920 14146 489972 14152
rect 486424 14136 486476 14142
rect 486424 14078 486476 14084
rect 485226 9344 485282 9353
rect 485226 9279 485282 9288
rect 482836 3528 482888 3534
rect 482836 3470 482888 3476
rect 483664 3528 483716 3534
rect 483664 3470 483716 3476
rect 482848 480 482876 3470
rect 484030 3360 484086 3369
rect 484030 3295 484086 3304
rect 484044 480 484072 3295
rect 485240 480 485268 9279
rect 486436 480 486464 14078
rect 488814 9208 488870 9217
rect 488814 9143 488870 9152
rect 487620 3596 487672 3602
rect 487620 3538 487672 3544
rect 487632 480 487660 3538
rect 488828 480 488856 9143
rect 489932 480 489960 14146
rect 492310 9072 492366 9081
rect 492310 9007 492366 9016
rect 491116 3936 491168 3942
rect 491116 3878 491168 3884
rect 491128 480 491156 3878
rect 492324 480 492352 9007
rect 493520 480 493548 14214
rect 495900 9036 495952 9042
rect 495900 8978 495952 8984
rect 494704 3664 494756 3670
rect 494704 3606 494756 3612
rect 494716 480 494744 3606
rect 495912 480 495940 8978
rect 497108 480 497136 14282
rect 499396 8968 499448 8974
rect 499396 8910 499448 8916
rect 498200 3732 498252 3738
rect 498200 3674 498252 3680
rect 498212 480 498240 3674
rect 499408 480 499436 8910
rect 500604 480 500632 14350
rect 501800 480 501828 16546
rect 504180 15156 504232 15162
rect 504180 15098 504232 15104
rect 502982 8936 503038 8945
rect 502982 8871 503038 8880
rect 502996 480 503024 8871
rect 504192 480 504220 15098
rect 507676 15088 507728 15094
rect 507676 15030 507728 15036
rect 506480 4004 506532 4010
rect 506480 3946 506532 3952
rect 505376 3800 505428 3806
rect 505376 3742 505428 3748
rect 505388 480 505416 3742
rect 506492 480 506520 3946
rect 507688 480 507716 15030
rect 508884 480 508912 16546
rect 511264 15020 511316 15026
rect 511264 14962 511316 14968
rect 510068 4140 510120 4146
rect 510068 4082 510120 4088
rect 510080 480 510108 4082
rect 511276 480 511304 14962
rect 512460 4276 512512 4282
rect 512460 4218 512512 4224
rect 512472 480 512500 4218
rect 512656 3602 512684 53246
rect 519544 53236 519596 53242
rect 519544 53178 519596 53184
rect 519556 16574 519584 53178
rect 520280 53168 520332 53174
rect 520280 53110 520332 53116
rect 520292 16574 520320 53110
rect 526444 53100 526496 53106
rect 526444 53042 526496 53048
rect 519556 16546 519676 16574
rect 520292 16546 520780 16574
rect 514760 14952 514812 14958
rect 514760 14894 514812 14900
rect 513564 3868 513616 3874
rect 513564 3810 513616 3816
rect 512644 3596 512696 3602
rect 512644 3538 512696 3544
rect 513576 480 513604 3810
rect 514772 480 514800 14894
rect 518348 14884 518400 14890
rect 518348 14826 518400 14832
rect 515956 4344 516008 4350
rect 515956 4286 516008 4292
rect 515968 480 515996 4286
rect 517152 4072 517204 4078
rect 517152 4014 517204 4020
rect 517164 480 517192 4014
rect 518360 480 518388 14826
rect 519544 4412 519596 4418
rect 519544 4354 519596 4360
rect 519556 480 519584 4354
rect 519648 3670 519676 16546
rect 519636 3664 519688 3670
rect 519636 3606 519688 3612
rect 520752 480 520780 16546
rect 521844 14816 521896 14822
rect 521844 14758 521896 14764
rect 521856 480 521884 14758
rect 525432 14748 525484 14754
rect 525432 14690 525484 14696
rect 523040 4480 523092 4486
rect 523040 4422 523092 4428
rect 523052 480 523080 4422
rect 524236 3528 524288 3534
rect 524236 3470 524288 3476
rect 524248 480 524276 3470
rect 525444 480 525472 14690
rect 526456 3534 526484 53042
rect 530584 51740 530636 51746
rect 530584 51682 530636 51688
rect 529020 14680 529072 14686
rect 529020 14622 529072 14628
rect 526628 4548 526680 4554
rect 526628 4490 526680 4496
rect 526444 3528 526496 3534
rect 526444 3470 526496 3476
rect 526640 480 526668 4490
rect 527824 3596 527876 3602
rect 527824 3538 527876 3544
rect 527836 480 527864 3538
rect 529032 480 529060 14622
rect 530124 4616 530176 4622
rect 530124 4558 530176 4564
rect 530136 480 530164 4558
rect 530596 3602 530624 51682
rect 533344 50720 533396 50726
rect 533344 50662 533396 50668
rect 532516 14612 532568 14618
rect 532516 14554 532568 14560
rect 531320 3664 531372 3670
rect 531320 3606 531372 3612
rect 530584 3596 530636 3602
rect 530584 3538 530636 3544
rect 531332 480 531360 3606
rect 532528 480 532556 14554
rect 533356 3670 533384 50662
rect 537484 50652 537536 50658
rect 537484 50594 537536 50600
rect 536104 14544 536156 14550
rect 536104 14486 536156 14492
rect 533712 4684 533764 4690
rect 533712 4626 533764 4632
rect 533344 3664 533396 3670
rect 533344 3606 533396 3612
rect 533724 480 533752 4626
rect 534908 3528 534960 3534
rect 534908 3470 534960 3476
rect 534920 480 534948 3470
rect 536116 480 536144 14486
rect 537208 4752 537260 4758
rect 537208 4694 537260 4700
rect 537220 480 537248 4694
rect 537496 3738 537524 50594
rect 542360 50584 542412 50590
rect 542360 50526 542412 50532
rect 542372 16574 542400 50526
rect 542372 16546 543228 16574
rect 539600 14476 539652 14482
rect 539600 14418 539652 14424
rect 538404 10260 538456 10266
rect 538404 10202 538456 10208
rect 537484 3732 537536 3738
rect 537484 3674 537536 3680
rect 538416 480 538444 10202
rect 539612 480 539640 14418
rect 541992 11008 542044 11014
rect 541992 10950 542044 10956
rect 540796 5500 540848 5506
rect 540796 5442 540848 5448
rect 540808 480 540836 5442
rect 542004 480 542032 10950
rect 543200 480 543228 16546
rect 544292 5432 544344 5438
rect 544292 5374 544344 5380
rect 544304 2802 544332 5374
rect 544396 3534 544424 54470
rect 551284 50516 551336 50522
rect 551284 50458 551336 50464
rect 546500 50448 546552 50454
rect 546500 50390 546552 50396
rect 546512 16574 546540 50390
rect 546512 16546 546724 16574
rect 545488 10940 545540 10946
rect 545488 10882 545540 10888
rect 544384 3528 544436 3534
rect 544384 3470 544436 3476
rect 544304 2774 544424 2802
rect 544396 480 544424 2774
rect 545500 480 545528 10882
rect 546696 480 546724 16546
rect 547880 10872 547932 10878
rect 547880 10814 547932 10820
rect 547892 3398 547920 10814
rect 547972 5364 548024 5370
rect 547972 5306 548024 5312
rect 547880 3392 547932 3398
rect 547880 3334 547932 3340
rect 547984 2666 548012 5306
rect 551296 3602 551324 50458
rect 560300 50380 560352 50386
rect 560300 50322 560352 50328
rect 560312 16574 560340 50322
rect 560312 16546 560892 16574
rect 552664 10804 552716 10810
rect 552664 10746 552716 10752
rect 551468 5296 551520 5302
rect 551468 5238 551520 5244
rect 550272 3596 550324 3602
rect 550272 3538 550324 3544
rect 551284 3596 551336 3602
rect 551284 3538 551336 3544
rect 549076 3392 549128 3398
rect 549076 3334 549128 3340
rect 547892 2638 548012 2666
rect 547892 480 547920 2638
rect 549088 480 549116 3334
rect 550284 480 550312 3538
rect 551480 480 551508 5238
rect 552676 480 552704 10746
rect 556160 10736 556212 10742
rect 556160 10678 556212 10684
rect 554964 5228 555016 5234
rect 554964 5170 555016 5176
rect 553768 3664 553820 3670
rect 553768 3606 553820 3612
rect 553780 480 553808 3606
rect 554976 480 555004 5170
rect 556172 480 556200 10678
rect 559748 10668 559800 10674
rect 559748 10610 559800 10616
rect 558552 5160 558604 5166
rect 558552 5102 558604 5108
rect 557356 3732 557408 3738
rect 557356 3674 557408 3680
rect 557368 480 557396 3674
rect 558564 480 558592 5102
rect 559760 480 559788 10610
rect 560864 480 560892 16546
rect 563244 10600 563296 10606
rect 563244 10542 563296 10548
rect 562048 5092 562100 5098
rect 562048 5034 562100 5040
rect 562060 480 562088 5034
rect 563256 480 563284 10542
rect 564452 480 564480 55830
rect 580276 46345 580304 230551
rect 580354 228304 580410 228313
rect 580354 228239 580410 228248
rect 580368 73001 580396 228239
rect 580354 72992 580410 73001
rect 580354 72927 580410 72936
rect 580262 46336 580318 46345
rect 580262 46271 580318 46280
rect 580356 46232 580408 46238
rect 580356 46174 580408 46180
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 580080 20664 580132 20670
rect 580080 20606 580132 20612
rect 580092 19825 580120 20606
rect 580078 19816 580134 19825
rect 580078 19751 580134 19760
rect 575112 15972 575164 15978
rect 575112 15914 575164 15920
rect 566832 10532 566884 10538
rect 566832 10474 566884 10480
rect 565636 5024 565688 5030
rect 565636 4966 565688 4972
rect 565648 480 565676 4966
rect 566844 480 566872 10474
rect 570328 10464 570380 10470
rect 570328 10406 570380 10412
rect 569132 4956 569184 4962
rect 569132 4898 569184 4904
rect 568028 3528 568080 3534
rect 568028 3470 568080 3476
rect 568040 480 568068 3470
rect 569144 480 569172 4898
rect 570340 480 570368 10406
rect 572720 10396 572772 10402
rect 572720 10338 572772 10344
rect 571524 3596 571576 3602
rect 571524 3538 571576 3544
rect 571536 480 571564 3538
rect 572732 3534 572760 10338
rect 572812 4888 572864 4894
rect 572812 4830 572864 4836
rect 572720 3528 572772 3534
rect 572720 3470 572772 3476
rect 572824 2530 572852 4830
rect 573916 3528 573968 3534
rect 573916 3470 573968 3476
rect 572732 2502 572852 2530
rect 572732 480 572760 2502
rect 573928 480 573956 3470
rect 575124 480 575152 15914
rect 578608 15904 578660 15910
rect 578608 15846 578660 15852
rect 577412 10328 577464 10334
rect 577412 10270 577464 10276
rect 576308 4820 576360 4826
rect 576308 4762 576360 4768
rect 576320 480 576348 4762
rect 577424 480 577452 10270
rect 578620 480 578648 15846
rect 580368 6633 580396 46174
rect 582194 11792 582250 11801
rect 582194 11727 582250 11736
rect 580354 6624 580410 6633
rect 580354 6559 580410 6568
rect 581000 3460 581052 3466
rect 581000 3402 581052 3408
rect 581012 480 581040 3402
rect 582208 480 582236 11727
rect 583390 11656 583446 11665
rect 583390 11591 583446 11600
rect 583404 480 583432 11591
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 3422 410488 3478 410544
rect 3514 397468 3516 397488
rect 3516 397468 3568 397488
rect 3568 397468 3570 397488
rect 3514 397432 3570 397468
rect 3422 371320 3478 371376
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3422 319232 3478 319288
rect 3238 306176 3294 306232
rect 3422 293120 3478 293176
rect 3054 267144 3110 267200
rect 53654 488688 53710 488744
rect 53286 488552 53342 488608
rect 3422 254088 3478 254144
rect 4066 241032 4122 241088
rect 3422 236680 3478 236736
rect 4158 233824 4214 233880
rect 17222 233416 17278 233472
rect 3514 232192 3570 232248
rect 3422 228248 3478 228304
rect 3054 214920 3110 214976
rect 3330 188844 3332 188864
rect 3332 188844 3384 188864
rect 3384 188844 3386 188864
rect 3330 188808 3386 188844
rect 3054 162832 3110 162888
rect 3054 136720 3110 136776
rect 3330 110608 3386 110664
rect 3238 97552 3294 97608
rect 2962 84632 3018 84688
rect 3330 71576 3386 71632
rect 3330 45500 3332 45520
rect 3332 45500 3384 45520
rect 3384 45500 3386 45520
rect 3330 45464 3386 45500
rect 2778 32408 2834 32464
rect 4802 232056 4858 232112
rect 3606 228520 3662 228576
rect 3790 228384 3846 228440
rect 3698 227024 3754 227080
rect 3790 201864 3846 201920
rect 3698 149776 3754 149832
rect 3606 58520 3662 58576
rect 3514 19352 3570 19408
rect 3422 6432 3478 6488
rect 4066 57160 4122 57216
rect 11702 231240 11758 231296
rect 7562 229064 7618 229120
rect 14462 231104 14518 231160
rect 15842 230968 15898 231024
rect 21362 233280 21418 233336
rect 18602 229200 18658 229256
rect 12346 57568 12402 57624
rect 10966 57432 11022 57488
rect 9586 57296 9642 57352
rect 15106 57024 15162 57080
rect 13726 56888 13782 56944
rect 32402 232464 32458 232520
rect 29642 232328 29698 232384
rect 53470 486512 53526 486568
rect 53378 483248 53434 483304
rect 53562 483384 53618 483440
rect 58806 487872 58862 487928
rect 54758 487736 54814 487792
rect 54666 487192 54722 487248
rect 53746 485832 53802 485888
rect 54482 242120 54538 242176
rect 58714 487600 58770 487656
rect 54942 487464 54998 487520
rect 54850 485560 54906 485616
rect 56874 487328 56930 487384
rect 55126 484744 55182 484800
rect 55034 484472 55090 484528
rect 56598 432248 56654 432304
rect 22006 56752 22062 56808
rect 55954 235320 56010 235376
rect 55862 206216 55918 206272
rect 56046 136992 56102 137048
rect 55954 121216 56010 121272
rect 56230 239536 56286 239592
rect 56138 108704 56194 108760
rect 56414 236544 56470 236600
rect 56414 215736 56470 215792
rect 56322 184184 56378 184240
rect 56506 165280 56562 165336
rect 56782 227160 56838 227216
rect 56690 226616 56746 226672
rect 56598 105576 56654 105632
rect 56230 83544 56286 83600
rect 56782 149640 56838 149696
rect 56690 77152 56746 77208
rect 58438 485288 58494 485344
rect 57518 483928 57574 483984
rect 57334 435376 57390 435432
rect 57242 433336 57298 433392
rect 57150 429392 57206 429448
rect 57058 407496 57114 407552
rect 57426 427896 57482 427952
rect 57242 243616 57298 243672
rect 57150 243480 57206 243536
rect 57058 226208 57114 226264
rect 57058 187448 57114 187504
rect 57150 102312 57206 102368
rect 57334 239400 57390 239456
rect 57242 96056 57298 96112
rect 57794 436328 57850 436384
rect 57610 430616 57666 430672
rect 57518 221992 57574 222048
rect 57518 212608 57574 212664
rect 57518 196832 57574 196888
rect 57518 193704 57574 193760
rect 57518 190576 57574 190632
rect 57518 181056 57574 181112
rect 57518 177964 57520 177984
rect 57520 177964 57572 177984
rect 57572 177964 57574 177984
rect 57518 177928 57574 177964
rect 57518 174800 57574 174856
rect 57426 159024 57482 159080
rect 57518 155916 57574 155952
rect 57518 155896 57520 155916
rect 57520 155896 57572 155916
rect 57572 155896 57574 155916
rect 57518 152768 57574 152824
rect 57426 146512 57482 146568
rect 57518 143248 57574 143304
rect 57426 133864 57482 133920
rect 57610 130736 57666 130792
rect 57334 89800 57390 89856
rect 57610 118088 57666 118144
rect 57610 111832 57666 111888
rect 57426 86672 57482 86728
rect 57702 74024 57758 74080
rect 57610 70896 57666 70952
rect 56874 64640 56930 64696
rect 57058 61512 57114 61568
rect 57886 409944 57942 410000
rect 58346 250416 58402 250472
rect 58254 240760 58310 240816
rect 58070 238040 58126 238096
rect 57886 226344 57942 226400
rect 57886 209480 57942 209536
rect 58162 235184 58218 235240
rect 58162 218864 58218 218920
rect 58070 162152 58126 162208
rect 58254 124480 58310 124536
rect 58530 485152 58586 485208
rect 58530 230016 58586 230072
rect 58438 229880 58494 229936
rect 58346 114960 58402 115016
rect 58714 199960 58770 200016
rect 59082 489912 59138 489968
rect 58990 484608 59046 484664
rect 58806 168544 58862 168600
rect 58622 140120 58678 140176
rect 58990 127608 59046 127664
rect 59266 488960 59322 489016
rect 59174 488824 59230 488880
rect 59082 99184 59138 99240
rect 59174 92928 59230 92984
rect 59358 408176 59414 408232
rect 88338 485288 88394 485344
rect 118606 490048 118662 490104
rect 158534 488008 158590 488064
rect 133602 487872 133658 487928
rect 118606 486376 118662 486432
rect 138570 487736 138626 487792
rect 143722 487736 143778 487792
rect 153934 487600 153990 487656
rect 133602 485832 133658 485888
rect 138570 485832 138626 485888
rect 143722 485832 143778 485888
rect 153934 485832 153990 485888
rect 158534 485832 158590 485888
rect 104898 485152 104954 485208
rect 59266 80280 59322 80336
rect 85486 398112 85542 398168
rect 92294 398112 92350 398168
rect 95882 398112 95938 398168
rect 59818 226752 59874 226808
rect 59542 203088 59598 203144
rect 59450 171672 59506 171728
rect 61382 227160 61438 227216
rect 76194 397296 76250 397352
rect 78310 397296 78366 397352
rect 79598 397296 79654 397352
rect 80426 397296 80482 397352
rect 82358 397296 82414 397352
rect 83002 397296 83058 397352
rect 60186 226752 60242 226808
rect 61750 226480 61806 226536
rect 62670 226752 62726 226808
rect 77206 396752 77262 396808
rect 89350 397296 89406 397352
rect 90086 397296 90142 397352
rect 91466 397296 91522 397352
rect 85394 396752 85450 396808
rect 86866 396752 86922 396808
rect 88246 396752 88302 396808
rect 89534 396752 89590 396808
rect 77206 245656 77262 245712
rect 67362 234640 67418 234696
rect 65982 230696 66038 230752
rect 63222 229744 63278 229800
rect 64142 229336 64198 229392
rect 65062 227840 65118 227896
rect 75642 231920 75698 231976
rect 68742 230832 68798 230888
rect 70398 230560 70454 230616
rect 70398 229744 70454 229800
rect 74538 229744 74594 229800
rect 70306 229608 70362 229664
rect 71686 229472 71742 229528
rect 71686 228520 71742 228576
rect 74538 228384 74594 228440
rect 73342 228112 73398 228168
rect 70582 227976 70638 228032
rect 70306 227024 70362 227080
rect 70030 226888 70086 226944
rect 72422 227704 72478 227760
rect 74262 227024 74318 227080
rect 76194 228384 76250 228440
rect 79322 237904 79378 237960
rect 84474 228928 84530 228984
rect 85486 228928 85542 228984
rect 87234 228928 87290 228984
rect 90914 396752 90970 396808
rect 93490 397296 93546 397352
rect 95054 397296 95110 397352
rect 92478 396752 92534 396808
rect 88246 228928 88302 228984
rect 90270 230424 90326 230480
rect 91006 230424 91062 230480
rect 98090 397296 98146 397352
rect 102782 397296 102838 397352
rect 104806 397296 104862 397352
rect 106094 397296 106150 397352
rect 106922 397296 106978 397352
rect 108854 397296 108910 397352
rect 109130 397296 109186 397352
rect 96526 396752 96582 396808
rect 97906 396752 97962 396808
rect 92478 239536 92534 239592
rect 93214 230424 93270 230480
rect 93766 230424 93822 230480
rect 95606 228928 95662 228984
rect 96526 233960 96582 234016
rect 96434 228928 96490 228984
rect 101954 396888 102010 396944
rect 99286 396752 99342 396808
rect 100666 396752 100722 396808
rect 100758 396616 100814 396672
rect 98734 230424 98790 230480
rect 99286 230424 99342 230480
rect 102046 396752 102102 396808
rect 101862 246336 101918 246392
rect 103518 396752 103574 396808
rect 102046 246336 102102 246392
rect 100758 238040 100814 238096
rect 106002 396752 106058 396808
rect 104254 230424 104310 230480
rect 107474 396752 107530 396808
rect 107658 396616 107714 396672
rect 106002 240896 106058 240952
rect 104806 230424 104862 230480
rect 106646 253952 106702 254008
rect 111614 396752 111670 396808
rect 111522 396616 111578 396672
rect 107658 235320 107714 235376
rect 110418 253816 110474 253872
rect 110418 251776 110474 251832
rect 111614 239536 111670 239592
rect 113638 398112 113694 398168
rect 112350 397296 112406 397352
rect 113362 397296 113418 397352
rect 113822 397296 113878 397352
rect 115754 396752 115810 396808
rect 113454 227568 113510 227624
rect 115754 236816 115810 236872
rect 118238 397296 118294 397352
rect 118606 397296 118662 397352
rect 117226 396752 117282 396808
rect 115938 396616 115994 396672
rect 119986 396752 120042 396808
rect 121274 396752 121330 396808
rect 114466 227568 114522 227624
rect 118698 251776 118754 251832
rect 118974 227568 119030 227624
rect 121274 247560 121330 247616
rect 136454 397296 136510 397352
rect 124126 396752 124182 396808
rect 126886 396752 126942 396808
rect 129646 396752 129702 396808
rect 131026 396752 131082 396808
rect 133786 396752 133842 396808
rect 121550 230016 121606 230072
rect 119986 227568 120042 227624
rect 124126 238040 124182 238096
rect 124218 233688 124274 233744
rect 123390 229880 123446 229936
rect 124862 233688 124918 233744
rect 126886 235320 126942 235376
rect 126978 233688 127034 233744
rect 139306 396752 139362 396808
rect 129646 249056 129702 249112
rect 127622 233688 127678 233744
rect 129738 233688 129794 233744
rect 130382 233688 130438 233744
rect 132498 233688 132554 233744
rect 133142 233688 133198 233744
rect 135258 233688 135314 233744
rect 135902 233688 135958 233744
rect 138018 233688 138074 233744
rect 138662 233688 138718 233744
rect 154118 397296 154174 397352
rect 163870 397296 163926 397352
rect 142066 396752 142122 396808
rect 144826 396752 144882 396808
rect 145010 396752 145066 396808
rect 148966 396752 149022 396808
rect 151726 396752 151782 396808
rect 140778 233688 140834 233744
rect 141422 233688 141478 233744
rect 155958 396752 156014 396808
rect 158626 396752 158682 396808
rect 161386 396752 161442 396808
rect 150806 236680 150862 236736
rect 149702 233824 149758 233880
rect 155406 233416 155462 233472
rect 152094 231240 152150 231296
rect 154854 231104 154910 231160
rect 153934 229744 153990 229800
rect 153014 229064 153070 229120
rect 161018 233280 161074 233336
rect 158166 232464 158222 232520
rect 158626 232464 158682 232520
rect 157614 230968 157670 231024
rect 156694 229608 156750 229664
rect 155866 229200 155922 229256
rect 155866 228248 155922 228304
rect 160190 232328 160246 232384
rect 158718 232192 158774 232248
rect 158718 229744 158774 229800
rect 159454 229064 159510 229120
rect 162858 232056 162914 232112
rect 162214 229472 162270 229528
rect 164974 229744 165030 229800
rect 164054 229200 164110 229256
rect 166906 396752 166962 396808
rect 168378 233824 168434 233880
rect 166906 233688 166962 233744
rect 167826 229744 167882 229800
rect 169298 233824 169354 233880
rect 171506 229880 171562 229936
rect 174266 230016 174322 230072
rect 177302 233688 177358 233744
rect 183466 397296 183522 397352
rect 182178 396752 182234 396808
rect 177946 233688 178002 233744
rect 181166 233688 181222 233744
rect 179786 230288 179842 230344
rect 182178 250416 182234 250472
rect 182086 233688 182142 233744
rect 183926 233688 183982 233744
rect 182638 230152 182694 230208
rect 182178 229336 182234 229392
rect 182178 228248 182234 228304
rect 184846 233688 184902 233744
rect 186318 229608 186374 229664
rect 188158 230424 188214 230480
rect 192206 233688 192262 233744
rect 190734 230288 190790 230344
rect 190918 230288 190974 230344
rect 190826 230016 190882 230072
rect 190458 229880 190514 229936
rect 190458 229744 190514 229800
rect 190642 229744 190698 229800
rect 190458 229472 190514 229528
rect 193126 233688 193182 233744
rect 197450 485424 197506 485480
rect 196806 485016 196862 485072
rect 196714 484880 196770 484936
rect 197358 484744 197414 484800
rect 196806 230288 196862 230344
rect 197358 230016 197414 230072
rect 197634 484064 197690 484120
rect 197542 483928 197598 483984
rect 197450 229880 197506 229936
rect 197542 229744 197598 229800
rect 196714 229608 196770 229664
rect 197726 417696 197782 417752
rect 201038 486240 201094 486296
rect 200854 485832 200910 485888
rect 200762 485016 200818 485072
rect 198646 484880 198702 484936
rect 197726 239400 197782 239456
rect 198094 230288 198150 230344
rect 197634 229472 197690 229528
rect 199382 479168 199438 479224
rect 198738 416336 198794 416392
rect 198738 243616 198794 243672
rect 199658 419328 199714 419384
rect 199474 414840 199530 414896
rect 199382 234096 199438 234152
rect 199290 230288 199346 230344
rect 199566 413616 199622 413672
rect 200486 233688 200542 233744
rect 199566 232600 199622 232656
rect 199474 228520 199530 228576
rect 201038 322088 201094 322144
rect 202142 487872 202198 487928
rect 201406 233688 201462 233744
rect 200762 230424 200818 230480
rect 204258 487736 204314 487792
rect 202142 230152 202198 230208
rect 206006 230424 206062 230480
rect 209134 486920 209190 486976
rect 209318 486104 209374 486160
rect 209686 484744 209742 484800
rect 209318 260072 209374 260128
rect 209134 239400 209190 239456
rect 206926 230424 206982 230480
rect 208766 230424 208822 230480
rect 210514 486648 210570 486704
rect 209686 230424 209742 230480
rect 211158 485152 211214 485208
rect 210514 229744 210570 229800
rect 213274 486784 213330 486840
rect 211158 230424 211214 230480
rect 211986 230424 212042 230480
rect 214562 487192 214618 487248
rect 213458 486512 213514 486568
rect 213642 486376 213698 486432
rect 213918 485288 213974 485344
rect 213458 250416 213514 250472
rect 214562 484472 214618 484528
rect 215206 484472 215262 484528
rect 213274 234232 213330 234288
rect 214470 230424 214526 230480
rect 218702 490048 218758 490104
rect 217966 487600 218022 487656
rect 216310 487056 216366 487112
rect 216034 485968 216090 486024
rect 215206 230424 215262 230480
rect 216218 483656 216274 483712
rect 217506 436872 217562 436928
rect 216678 431024 216734 431080
rect 217414 429936 217470 429992
rect 217230 409944 217286 410000
rect 216678 408348 216680 408368
rect 216680 408348 216732 408368
rect 216732 408348 216734 408368
rect 216678 408312 216734 408348
rect 217138 408040 217194 408096
rect 216310 232736 216366 232792
rect 216402 230424 216458 230480
rect 216218 230288 216274 230344
rect 216034 229880 216090 229936
rect 217690 435920 217746 435976
rect 217598 428168 217654 428224
rect 217782 433744 217838 433800
rect 217230 242256 217286 242312
rect 217874 432792 217930 432848
rect 217782 238176 217838 238232
rect 217874 231104 217930 231160
rect 218150 486648 218206 486704
rect 218058 483792 218114 483848
rect 218426 486512 218482 486568
rect 218242 486240 218298 486296
rect 218334 483520 218390 483576
rect 218610 485968 218666 486024
rect 218518 484200 218574 484256
rect 218334 231512 218390 231568
rect 260838 489912 260894 489968
rect 218978 489232 219034 489288
rect 218886 488008 218942 488064
rect 218794 486920 218850 486976
rect 218794 398112 218850 398168
rect 219898 489096 219954 489152
rect 219806 487736 219862 487792
rect 219346 486376 219402 486432
rect 219254 485832 219310 485888
rect 219162 485288 219218 485344
rect 219070 483520 219126 483576
rect 218978 397976 219034 398032
rect 218886 231376 218942 231432
rect 218702 231240 218758 231296
rect 218518 230968 218574 231024
rect 217138 228656 217194 228712
rect 217782 230424 217838 230480
rect 219070 230424 219126 230480
rect 219254 227160 219310 227216
rect 62946 226616 63002 226672
rect 71686 226616 71742 226672
rect 62762 226344 62818 226400
rect 68190 226344 68246 226400
rect 219714 485152 219770 485208
rect 219530 483928 219586 483984
rect 219622 483656 219678 483712
rect 253386 488960 253442 489016
rect 219990 486104 220046 486160
rect 219806 398112 219862 398168
rect 258354 488824 258410 488880
rect 288530 489232 288586 489288
rect 278410 488688 278466 488744
rect 266082 487872 266138 487928
rect 260838 486512 260894 486568
rect 273258 486376 273314 486432
rect 253386 485832 253442 485888
rect 258354 485832 258410 485888
rect 266082 485832 266138 485888
rect 295890 489096 295946 489152
rect 288530 486240 288586 486296
rect 310978 488552 311034 488608
rect 301502 487328 301558 487384
rect 301502 486512 301558 486568
rect 295890 486104 295946 486160
rect 313554 487736 313610 487792
rect 320270 487600 320326 487656
rect 340142 487192 340198 487248
rect 340142 486376 340198 486432
rect 278410 485832 278466 485888
rect 310978 485832 311034 485888
rect 313554 485832 313610 485888
rect 320270 485832 320326 485888
rect 273258 485288 273314 485344
rect 356518 484472 356574 484528
rect 222106 251096 222162 251152
rect 222842 251096 222898 251152
rect 220542 230288 220598 230344
rect 219990 227296 220046 227352
rect 223302 230424 223358 230480
rect 224222 233824 224278 233880
rect 223670 228792 223726 228848
rect 61106 226208 61162 226264
rect 62026 226208 62082 226264
rect 219346 226208 219402 226264
rect 58898 67768 58954 67824
rect 58714 57840 58770 57896
rect 58622 57704 58678 57760
rect 58622 57296 58678 57352
rect 58530 57024 58586 57080
rect 58254 56888 58310 56944
rect 58254 56616 58310 56672
rect 60002 57432 60058 57488
rect 60922 57160 60978 57216
rect 62118 57704 62174 57760
rect 62762 57568 62818 57624
rect 63038 57432 63094 57488
rect 62486 57296 62542 57352
rect 63682 56888 63738 56944
rect 63314 56616 63370 56672
rect 65430 56752 65486 56808
rect 97906 3984 97962 4040
rect 99194 3848 99250 3904
rect 99286 3168 99342 3224
rect 100574 3576 100630 3632
rect 102046 3712 102102 3768
rect 101954 3440 102010 3496
rect 104806 3304 104862 3360
rect 127806 57024 127862 57080
rect 132958 57024 133014 57080
rect 149518 3984 149574 4040
rect 151634 6840 151690 6896
rect 151358 6704 151414 6760
rect 150622 3168 150678 3224
rect 153106 6568 153162 6624
rect 153014 3848 153070 3904
rect 157246 6432 157302 6488
rect 157154 6296 157210 6352
rect 161294 3712 161350 3768
rect 160098 3576 160154 3632
rect 165158 6160 165214 6216
rect 164882 3440 164938 3496
rect 169298 3168 169354 3224
rect 170770 3984 170826 4040
rect 180522 57160 180578 57216
rect 176198 3848 176254 3904
rect 175462 3304 175518 3360
rect 180798 57160 180854 57216
rect 181810 9424 181866 9480
rect 180706 3712 180762 3768
rect 181994 3576 182050 3632
rect 182086 3440 182142 3496
rect 183374 9288 183430 9344
rect 184754 9152 184810 9208
rect 184570 9016 184626 9072
rect 183098 3304 183154 3360
rect 187422 8880 187478 8936
rect 206926 57160 206982 57216
rect 208030 57568 208086 57624
rect 210146 58928 210202 58984
rect 211066 57704 211122 57760
rect 211618 56888 211674 56944
rect 208214 11736 208270 11792
rect 212538 59064 212594 59120
rect 212814 57840 212870 57896
rect 213182 57024 213238 57080
rect 211894 56752 211950 56808
rect 213734 57296 213790 57352
rect 216126 59744 216182 59800
rect 215206 57704 215262 57760
rect 214654 57432 214710 57488
rect 217598 59472 217654 59528
rect 218242 59880 218298 59936
rect 217506 56616 217562 56672
rect 208306 11600 208362 11656
rect 219990 59200 220046 59256
rect 219714 58792 219770 58848
rect 221186 59608 221242 59664
rect 219070 6024 219126 6080
rect 222382 59880 222438 59936
rect 222566 59780 222568 59800
rect 222568 59780 222620 59800
rect 222620 59780 222622 59800
rect 222566 59744 222622 59780
rect 222750 59744 222806 59800
rect 223026 59336 223082 59392
rect 223946 59880 224002 59936
rect 224130 59880 224186 59936
rect 224866 223080 224922 223136
rect 225326 249056 225382 249112
rect 225234 198600 225290 198656
rect 225142 193704 225198 193760
rect 225050 58792 225106 58848
rect 225418 238040 225474 238096
rect 225510 220632 225566 220688
rect 225694 228656 225750 228712
rect 225602 93064 225658 93120
rect 224314 57296 224370 57352
rect 225786 228520 225842 228576
rect 225970 247560 226026 247616
rect 226062 235320 226118 235376
rect 226246 233960 226302 234016
rect 226154 232464 226210 232520
rect 226154 213288 226210 213344
rect 226062 164192 226118 164248
rect 225970 151952 226026 152008
rect 225878 134816 225934 134872
rect 226798 227160 226854 227216
rect 226706 183912 226762 183968
rect 226614 176568 226670 176624
rect 226614 175208 226670 175264
rect 226614 174120 226670 174176
rect 226522 159296 226578 159352
rect 226522 150320 226578 150376
rect 226522 149504 226578 149560
rect 226522 140664 226578 140720
rect 226522 139712 226578 139768
rect 226430 120128 226486 120184
rect 226338 88168 226394 88224
rect 226522 84088 226578 84144
rect 226522 83272 226578 83328
rect 226522 77152 226578 77208
rect 226522 75928 226578 75984
rect 227166 250416 227222 250472
rect 226982 231240 227038 231296
rect 226890 154400 226946 154456
rect 227074 225936 227130 225992
rect 226982 144608 227038 144664
rect 227350 239400 227406 239456
rect 227258 227296 227314 227352
rect 227166 171536 227222 171592
rect 227534 234232 227590 234288
rect 227442 229744 227498 229800
rect 227350 188808 227406 188864
rect 227626 231376 227682 231432
rect 227626 215736 227682 215792
rect 227626 209616 227682 209672
rect 227626 208392 227682 208448
rect 227534 196152 227590 196208
rect 227442 181464 227498 181520
rect 227258 166640 227314 166696
rect 227074 142160 227130 142216
rect 226798 71032 226854 71088
rect 226522 64776 226578 64832
rect 226522 63688 226578 63744
rect 227810 179016 227866 179072
rect 228086 240896 228142 240952
rect 227994 210840 228050 210896
rect 227902 68584 227958 68640
rect 228178 234096 228234 234152
rect 228086 57704 228142 57760
rect 228270 232600 228326 232656
rect 228178 57568 228234 57624
rect 226246 56752 226302 56808
rect 228638 186360 228694 186416
rect 228546 169088 228602 169144
rect 228454 112648 228510 112704
rect 228362 105304 228418 105360
rect 229834 239536 229890 239592
rect 229742 231104 229798 231160
rect 229650 147056 229706 147112
rect 229926 236816 229982 236872
rect 229926 218184 229982 218240
rect 229834 203496 229890 203552
rect 229742 117680 229798 117736
rect 230754 61240 230810 61296
rect 230938 60152 230994 60208
rect 231214 238176 231270 238232
rect 231122 78376 231178 78432
rect 231030 59608 231086 59664
rect 230846 59336 230902 59392
rect 231398 205944 231454 206000
rect 231306 161744 231362 161800
rect 232410 242256 232466 242312
rect 232318 137264 232374 137320
rect 232226 129920 232282 129976
rect 232134 127472 232190 127528
rect 232042 122576 232098 122632
rect 231950 97960 232006 98016
rect 231858 85720 231914 85776
rect 232502 140664 232558 140720
rect 235998 398112 236054 398168
rect 233238 95512 233294 95568
rect 232410 66136 232466 66192
rect 231214 57432 231270 57488
rect 234066 226752 234122 226808
rect 233974 110200 234030 110256
rect 229466 56616 229522 56672
rect 234434 228384 234490 228440
rect 234342 227024 234398 227080
rect 234434 218048 234490 218104
rect 235354 230696 235410 230752
rect 235262 209616 235318 209672
rect 234342 205672 234398 205728
rect 234250 191256 234306 191312
rect 234158 175208 234214 175264
rect 235262 120672 235318 120728
rect 235262 100408 235318 100464
rect 235538 226888 235594 226944
rect 235538 151816 235594 151872
rect 235446 150320 235502 150376
rect 235354 85584 235410 85640
rect 236182 397296 236238 397352
rect 239218 397296 239274 397352
rect 237378 396752 237434 396808
rect 240138 396752 240194 396808
rect 241518 396752 241574 396808
rect 236642 230832 236698 230888
rect 236734 228112 236790 228168
rect 236734 178064 236790 178120
rect 236642 125568 236698 125624
rect 238114 226480 238170 226536
rect 238022 125024 238078 125080
rect 239402 227976 239458 228032
rect 238298 201048 238354 201104
rect 239402 138080 239458 138136
rect 238206 102856 238262 102912
rect 240874 227840 240930 227896
rect 240782 157256 240838 157312
rect 241518 120672 241574 120728
rect 242898 396752 242954 396808
rect 244370 396752 244426 396808
rect 244554 396752 244610 396808
rect 242898 242120 242954 242176
rect 242254 91024 242310 91080
rect 242162 84088 242218 84144
rect 265070 398112 265126 398168
rect 300122 398112 300178 398168
rect 315762 398112 315818 398168
rect 325882 398112 325938 398168
rect 247682 397296 247738 397352
rect 247958 397296 248014 397352
rect 248602 397296 248658 397352
rect 250074 397296 250130 397352
rect 250350 397296 250406 397352
rect 252742 397296 252798 397352
rect 259458 397296 259514 397352
rect 260930 397296 260986 397352
rect 261942 397296 261998 397352
rect 262310 397296 262366 397352
rect 263598 397296 263654 397352
rect 245658 396752 245714 396808
rect 244922 64776 244978 64832
rect 246302 226616 246358 226672
rect 246302 165688 246358 165744
rect 251178 397024 251234 397080
rect 249062 132368 249118 132424
rect 251362 396752 251418 396808
rect 252558 396752 252614 396808
rect 251914 257896 251970 257952
rect 251914 237904 251970 237960
rect 258078 396888 258134 396944
rect 254122 396752 254178 396808
rect 255410 396752 255466 396808
rect 256146 396752 256202 396808
rect 256882 396772 256938 396808
rect 256882 396752 256884 396772
rect 256884 396752 256936 396772
rect 256936 396752 256938 396772
rect 253294 234640 253350 234696
rect 253294 111832 253350 111888
rect 258170 396752 258226 396808
rect 259550 396752 259606 396808
rect 255962 57024 256018 57080
rect 260746 245656 260802 245712
rect 263690 396752 263746 396808
rect 268290 397296 268346 397352
rect 268658 397296 268714 397352
rect 272338 397296 272394 397352
rect 275282 397332 275284 397352
rect 275284 397332 275336 397352
rect 275336 397332 275338 397352
rect 275282 397296 275338 397332
rect 277674 397296 277730 397352
rect 278870 397296 278926 397352
rect 290186 397296 290242 397352
rect 298466 397296 298522 397352
rect 265162 396772 265218 396808
rect 265162 396752 265164 396772
rect 265164 396752 265216 396772
rect 265216 396752 265218 396772
rect 266358 396752 266414 396808
rect 266450 396616 266506 396672
rect 269394 396772 269450 396808
rect 269394 396752 269396 396772
rect 269396 396752 269448 396772
rect 269448 396752 269450 396772
rect 270498 396752 270554 396808
rect 266358 59336 266414 59392
rect 270590 396616 270646 396672
rect 273350 396752 273406 396808
rect 273626 396752 273682 396808
rect 276110 396752 276166 396808
rect 277490 396752 277546 396808
rect 273442 396616 273498 396672
rect 276018 396616 276074 396672
rect 270498 240760 270554 240816
rect 271142 227704 271198 227760
rect 280158 396752 280214 396808
rect 283746 396772 283802 396808
rect 283746 396752 283748 396772
rect 283748 396752 283800 396772
rect 283800 396752 283802 396772
rect 285954 396752 286010 396808
rect 287058 396752 287114 396808
rect 292670 396772 292726 396808
rect 292670 396752 292672 396772
rect 292672 396752 292724 396772
rect 292724 396752 292726 396772
rect 295338 396752 295394 396808
rect 308586 397316 308642 397352
rect 308586 397296 308588 397316
rect 308588 397296 308640 397316
rect 308640 397296 308642 397316
rect 302238 396752 302294 396808
rect 304998 396752 305054 396808
rect 310518 396752 310574 396808
rect 313278 396752 313334 396808
rect 317418 396752 317474 396808
rect 320178 396752 320234 396808
rect 322938 396752 322994 396808
rect 320178 236544 320234 236600
rect 342626 397296 342682 397352
rect 342350 396752 342406 396808
rect 322938 235184 322994 235240
rect 357438 418784 357494 418840
rect 356518 77152 356574 77208
rect 357530 414296 357586 414352
rect 359002 478896 359058 478952
rect 358818 415792 358874 415848
rect 357530 243480 357586 243536
rect 358910 413072 358966 413128
rect 359094 417152 359150 417208
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580262 418240 580318 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 579618 365064 579674 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 579986 312024 580042 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 580262 230560 580318 230616
rect 410522 226344 410578 226400
rect 580170 192480 580226 192536
rect 580170 99456 580226 99512
rect 580170 59608 580226 59664
rect 358818 59064 358874 59120
rect 357438 58928 357494 58984
rect 251822 56888 251878 56944
rect 358726 6840 358782 6896
rect 362314 6704 362370 6760
rect 365810 6568 365866 6624
rect 379978 6432 380034 6488
rect 383566 6296 383622 6352
rect 390650 6024 390706 6080
rect 411902 6160 411958 6216
rect 436742 57160 436798 57216
rect 433246 3168 433302 3224
rect 436742 3984 436798 4040
rect 458086 3848 458142 3904
rect 472254 3712 472310 3768
rect 479338 3576 479394 3632
rect 481730 9424 481786 9480
rect 480534 3440 480590 3496
rect 485226 9288 485282 9344
rect 484030 3304 484086 3360
rect 488814 9152 488870 9208
rect 492310 9016 492366 9072
rect 502982 8880 503038 8936
rect 580354 228248 580410 228304
rect 580354 72936 580410 72992
rect 580262 46280 580318 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580078 19760 580134 19816
rect 582194 11736 582250 11792
rect 580354 6568 580410 6624
rect 583390 11600 583446 11656
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect 118601 490106 118667 490109
rect 218697 490106 218763 490109
rect 118601 490104 218763 490106
rect 118601 490048 118606 490104
rect 118662 490048 218702 490104
rect 218758 490048 218763 490104
rect 118601 490046 218763 490048
rect 118601 490043 118667 490046
rect 218697 490043 218763 490046
rect 59077 489970 59143 489973
rect 260833 489970 260899 489973
rect 59077 489968 260899 489970
rect 59077 489912 59082 489968
rect 59138 489912 260838 489968
rect 260894 489912 260899 489968
rect 59077 489910 260899 489912
rect 59077 489907 59143 489910
rect 260833 489907 260899 489910
rect 218973 489290 219039 489293
rect 288525 489290 288591 489293
rect 218973 489288 288591 489290
rect 218973 489232 218978 489288
rect 219034 489232 288530 489288
rect 288586 489232 288591 489288
rect 218973 489230 288591 489232
rect 218973 489227 219039 489230
rect 288525 489227 288591 489230
rect 219893 489154 219959 489157
rect 295885 489154 295951 489157
rect 219893 489152 295951 489154
rect 219893 489096 219898 489152
rect 219954 489096 295890 489152
rect 295946 489096 295951 489152
rect 219893 489094 295951 489096
rect 219893 489091 219959 489094
rect 295885 489091 295951 489094
rect 59261 489018 59327 489021
rect 253381 489018 253447 489021
rect 59261 489016 253447 489018
rect 59261 488960 59266 489016
rect 59322 488960 253386 489016
rect 253442 488960 253447 489016
rect 59261 488958 253447 488960
rect 59261 488955 59327 488958
rect 253381 488955 253447 488958
rect 59169 488882 59235 488885
rect 258349 488882 258415 488885
rect 59169 488880 258415 488882
rect -960 488596 480 488836
rect 59169 488824 59174 488880
rect 59230 488824 258354 488880
rect 258410 488824 258415 488880
rect 59169 488822 258415 488824
rect 59169 488819 59235 488822
rect 258349 488819 258415 488822
rect 53649 488746 53715 488749
rect 278405 488746 278471 488749
rect 53649 488744 278471 488746
rect 53649 488688 53654 488744
rect 53710 488688 278410 488744
rect 278466 488688 278471 488744
rect 53649 488686 278471 488688
rect 53649 488683 53715 488686
rect 278405 488683 278471 488686
rect 53281 488610 53347 488613
rect 310973 488610 311039 488613
rect 53281 488608 311039 488610
rect 53281 488552 53286 488608
rect 53342 488552 310978 488608
rect 311034 488552 311039 488608
rect 53281 488550 311039 488552
rect 53281 488547 53347 488550
rect 310973 488547 311039 488550
rect 158529 488066 158595 488069
rect 218881 488066 218947 488069
rect 158529 488064 218947 488066
rect 158529 488008 158534 488064
rect 158590 488008 218886 488064
rect 218942 488008 218947 488064
rect 158529 488006 218947 488008
rect 158529 488003 158595 488006
rect 218881 488003 218947 488006
rect 58801 487930 58867 487933
rect 133597 487930 133663 487933
rect 58801 487928 133663 487930
rect 58801 487872 58806 487928
rect 58862 487872 133602 487928
rect 133658 487872 133663 487928
rect 58801 487870 133663 487872
rect 58801 487867 58867 487870
rect 133597 487867 133663 487870
rect 202137 487930 202203 487933
rect 266077 487930 266143 487933
rect 202137 487928 266143 487930
rect 202137 487872 202142 487928
rect 202198 487872 266082 487928
rect 266138 487872 266143 487928
rect 202137 487870 266143 487872
rect 202137 487867 202203 487870
rect 266077 487867 266143 487870
rect 54753 487794 54819 487797
rect 138565 487794 138631 487797
rect 54753 487792 138631 487794
rect 54753 487736 54758 487792
rect 54814 487736 138570 487792
rect 138626 487736 138631 487792
rect 54753 487734 138631 487736
rect 54753 487731 54819 487734
rect 138565 487731 138631 487734
rect 143717 487794 143783 487797
rect 204253 487794 204319 487797
rect 143717 487792 204319 487794
rect 143717 487736 143722 487792
rect 143778 487736 204258 487792
rect 204314 487736 204319 487792
rect 143717 487734 204319 487736
rect 143717 487731 143783 487734
rect 204253 487731 204319 487734
rect 219801 487794 219867 487797
rect 313549 487794 313615 487797
rect 219801 487792 313615 487794
rect 219801 487736 219806 487792
rect 219862 487736 313554 487792
rect 313610 487736 313615 487792
rect 219801 487734 313615 487736
rect 219801 487731 219867 487734
rect 313549 487731 313615 487734
rect 58709 487658 58775 487661
rect 153929 487658 153995 487661
rect 58709 487656 153995 487658
rect 58709 487600 58714 487656
rect 58770 487600 153934 487656
rect 153990 487600 153995 487656
rect 58709 487598 153995 487600
rect 58709 487595 58775 487598
rect 153929 487595 153995 487598
rect 217961 487658 218027 487661
rect 320265 487658 320331 487661
rect 217961 487656 320331 487658
rect 217961 487600 217966 487656
rect 218022 487600 320270 487656
rect 320326 487600 320331 487656
rect 217961 487598 320331 487600
rect 217961 487595 218027 487598
rect 320265 487595 320331 487598
rect 54937 487522 55003 487525
rect 268510 487522 268516 487524
rect 54937 487520 268516 487522
rect 54937 487464 54942 487520
rect 54998 487464 268516 487520
rect 54937 487462 268516 487464
rect 54937 487459 55003 487462
rect 268510 487460 268516 487462
rect 268580 487460 268586 487524
rect 56869 487386 56935 487389
rect 301497 487386 301563 487389
rect 56869 487384 301563 487386
rect 56869 487328 56874 487384
rect 56930 487328 301502 487384
rect 301558 487328 301563 487384
rect 56869 487326 301563 487328
rect 56869 487323 56935 487326
rect 301497 487323 301563 487326
rect 54661 487250 54727 487253
rect 150934 487250 150940 487252
rect 54661 487248 150940 487250
rect 54661 487192 54666 487248
rect 54722 487192 150940 487248
rect 54661 487190 150940 487192
rect 54661 487187 54727 487190
rect 150934 487188 150940 487190
rect 151004 487188 151010 487252
rect 214557 487250 214623 487253
rect 340137 487250 340203 487253
rect 214557 487248 340203 487250
rect 214557 487192 214562 487248
rect 214618 487192 340142 487248
rect 340198 487192 340203 487248
rect 214557 487190 340203 487192
rect 214557 487187 214623 487190
rect 340137 487187 340203 487190
rect 90950 487052 90956 487116
rect 91020 487114 91026 487116
rect 216305 487114 216371 487117
rect 91020 487112 216371 487114
rect 91020 487056 216310 487112
rect 216366 487056 216371 487112
rect 91020 487054 216371 487056
rect 91020 487052 91026 487054
rect 216305 487051 216371 487054
rect 140998 486916 141004 486980
rect 141068 486978 141074 486980
rect 209129 486978 209195 486981
rect 141068 486976 209195 486978
rect 141068 486920 209134 486976
rect 209190 486920 209195 486976
rect 141068 486918 209195 486920
rect 141068 486916 141074 486918
rect 209129 486915 209195 486918
rect 218789 486978 218855 486981
rect 318374 486978 318380 486980
rect 218789 486976 318380 486978
rect 218789 486920 218794 486976
rect 218850 486920 318380 486976
rect 218789 486918 318380 486920
rect 218789 486915 218855 486918
rect 318374 486916 318380 486918
rect 318444 486916 318450 486980
rect 145598 486780 145604 486844
rect 145668 486842 145674 486844
rect 213269 486842 213335 486845
rect 145668 486840 213335 486842
rect 145668 486784 213274 486840
rect 213330 486784 213335 486840
rect 145668 486782 213335 486784
rect 145668 486780 145674 486782
rect 213269 486779 213335 486782
rect 136030 486644 136036 486708
rect 136100 486706 136106 486708
rect 210509 486706 210575 486709
rect 136100 486704 210575 486706
rect 136100 486648 210514 486704
rect 210570 486648 210575 486704
rect 136100 486646 210575 486648
rect 136100 486644 136106 486646
rect 210509 486643 210575 486646
rect 218145 486706 218211 486709
rect 256182 486706 256188 486708
rect 218145 486704 256188 486706
rect 218145 486648 218150 486704
rect 218206 486648 256188 486704
rect 218145 486646 256188 486648
rect 218145 486643 218211 486646
rect 256182 486644 256188 486646
rect 256252 486644 256258 486708
rect 263542 486706 263548 486708
rect 258030 486646 263548 486706
rect 53465 486570 53531 486573
rect 128670 486570 128676 486572
rect 53465 486568 128676 486570
rect 53465 486512 53470 486568
rect 53526 486512 128676 486568
rect 53465 486510 128676 486512
rect 53465 486507 53531 486510
rect 128670 486508 128676 486510
rect 128740 486508 128746 486572
rect 131062 486508 131068 486572
rect 131132 486570 131138 486572
rect 213453 486570 213519 486573
rect 131132 486568 213519 486570
rect 131132 486512 213458 486568
rect 213514 486512 213519 486568
rect 131132 486510 213519 486512
rect 131132 486508 131138 486510
rect 213453 486507 213519 486510
rect 218421 486570 218487 486573
rect 258030 486570 258090 486646
rect 263542 486644 263548 486646
rect 263612 486644 263618 486708
rect 218421 486568 258090 486570
rect 218421 486512 218426 486568
rect 218482 486512 258090 486568
rect 218421 486510 258090 486512
rect 260833 486570 260899 486573
rect 260966 486570 260972 486572
rect 260833 486568 260972 486570
rect 260833 486512 260838 486568
rect 260894 486512 260972 486568
rect 260833 486510 260972 486512
rect 218421 486507 218487 486510
rect 260833 486507 260899 486510
rect 260966 486508 260972 486510
rect 261036 486508 261042 486572
rect 273478 486570 273484 486572
rect 267690 486510 273484 486570
rect 118601 486436 118667 486437
rect 118550 486434 118556 486436
rect 118510 486374 118556 486434
rect 118620 486432 118667 486436
rect 118662 486376 118667 486432
rect 118550 486372 118556 486374
rect 118620 486372 118667 486376
rect 120758 486372 120764 486436
rect 120828 486434 120834 486436
rect 213637 486434 213703 486437
rect 120828 486432 213703 486434
rect 120828 486376 213642 486432
rect 213698 486376 213703 486432
rect 120828 486374 213703 486376
rect 120828 486372 120834 486374
rect 118601 486371 118667 486372
rect 213637 486371 213703 486374
rect 219341 486434 219407 486437
rect 267690 486434 267750 486510
rect 273478 486508 273484 486510
rect 273548 486508 273554 486572
rect 301497 486570 301563 486573
rect 339718 486570 339724 486572
rect 301497 486568 339724 486570
rect 301497 486512 301502 486568
rect 301558 486512 339724 486568
rect 301497 486510 339724 486512
rect 301497 486507 301563 486510
rect 339718 486508 339724 486510
rect 339788 486508 339794 486572
rect 219341 486432 267750 486434
rect 219341 486376 219346 486432
rect 219402 486376 267750 486432
rect 219341 486374 267750 486376
rect 273253 486434 273319 486437
rect 323342 486434 323348 486436
rect 273253 486432 323348 486434
rect 273253 486376 273258 486432
rect 273314 486376 323348 486432
rect 273253 486374 323348 486376
rect 219341 486371 219407 486374
rect 273253 486371 273319 486374
rect 323342 486372 323348 486374
rect 323412 486372 323418 486436
rect 340137 486434 340203 486437
rect 350758 486434 350764 486436
rect 340137 486432 350764 486434
rect 340137 486376 340142 486432
rect 340198 486376 350764 486432
rect 340137 486374 350764 486376
rect 340137 486371 340203 486374
rect 350758 486372 350764 486374
rect 350828 486372 350834 486436
rect 101070 486236 101076 486300
rect 101140 486298 101146 486300
rect 201033 486298 201099 486301
rect 101140 486296 201099 486298
rect 101140 486240 201038 486296
rect 201094 486240 201099 486296
rect 101140 486238 201099 486240
rect 101140 486236 101146 486238
rect 201033 486235 201099 486238
rect 218237 486298 218303 486301
rect 288525 486300 288591 486301
rect 283782 486298 283788 486300
rect 218237 486296 283788 486298
rect 218237 486240 218242 486296
rect 218298 486240 283788 486296
rect 218237 486238 283788 486240
rect 218237 486235 218303 486238
rect 283782 486236 283788 486238
rect 283852 486236 283858 486300
rect 288525 486296 288572 486300
rect 288636 486298 288642 486300
rect 288525 486240 288530 486296
rect 288525 486236 288572 486240
rect 288636 486238 288682 486298
rect 288636 486236 288642 486238
rect 288525 486235 288591 486236
rect 98494 486100 98500 486164
rect 98564 486162 98570 486164
rect 209313 486162 209379 486165
rect 98564 486160 209379 486162
rect 98564 486104 209318 486160
rect 209374 486104 209379 486160
rect 98564 486102 209379 486104
rect 98564 486100 98570 486102
rect 209313 486099 209379 486102
rect 219985 486162 220051 486165
rect 295885 486164 295951 486165
rect 290958 486162 290964 486164
rect 219985 486160 290964 486162
rect 219985 486104 219990 486160
rect 220046 486104 290964 486160
rect 219985 486102 290964 486104
rect 219985 486099 220051 486102
rect 290958 486100 290964 486102
rect 291028 486100 291034 486164
rect 295885 486160 295932 486164
rect 295996 486162 296002 486164
rect 295885 486104 295890 486160
rect 295885 486100 295932 486104
rect 295996 486102 296042 486162
rect 295996 486100 296002 486102
rect 295885 486099 295951 486100
rect 93526 485964 93532 486028
rect 93596 486026 93602 486028
rect 216029 486026 216095 486029
rect 93596 486024 216095 486026
rect 93596 485968 216034 486024
rect 216090 485968 216095 486024
rect 93596 485966 216095 485968
rect 93596 485964 93602 485966
rect 216029 485963 216095 485966
rect 218605 486026 218671 486029
rect 300710 486026 300716 486028
rect 218605 486024 300716 486026
rect 218605 485968 218610 486024
rect 218666 485968 300716 486024
rect 218605 485966 300716 485968
rect 218605 485963 218671 485966
rect 300710 485964 300716 485966
rect 300780 485964 300786 486028
rect 53741 485890 53807 485893
rect 133597 485892 133663 485893
rect 138565 485892 138631 485893
rect 111190 485890 111196 485892
rect 53741 485888 111196 485890
rect 53741 485832 53746 485888
rect 53802 485832 111196 485888
rect 53741 485830 111196 485832
rect 53741 485827 53807 485830
rect 111190 485828 111196 485830
rect 111260 485828 111266 485892
rect 133597 485888 133644 485892
rect 133708 485890 133714 485892
rect 133597 485832 133602 485888
rect 133597 485828 133644 485832
rect 133708 485830 133754 485890
rect 138565 485888 138612 485892
rect 138676 485890 138682 485892
rect 138565 485832 138570 485888
rect 133708 485828 133714 485830
rect 138565 485828 138612 485832
rect 138676 485830 138722 485890
rect 138676 485828 138682 485830
rect 143574 485828 143580 485892
rect 143644 485890 143650 485892
rect 143717 485890 143783 485893
rect 143644 485888 143783 485890
rect 143644 485832 143722 485888
rect 143778 485832 143783 485888
rect 143644 485830 143783 485832
rect 143644 485828 143650 485830
rect 133597 485827 133663 485828
rect 138565 485827 138631 485828
rect 143717 485827 143783 485830
rect 153929 485890 153995 485893
rect 158529 485892 158595 485893
rect 154062 485890 154068 485892
rect 153929 485888 154068 485890
rect 153929 485832 153934 485888
rect 153990 485832 154068 485888
rect 153929 485830 154068 485832
rect 153929 485827 153995 485830
rect 154062 485828 154068 485830
rect 154132 485828 154138 485892
rect 158478 485890 158484 485892
rect 158438 485830 158484 485890
rect 158548 485888 158595 485892
rect 158590 485832 158595 485888
rect 158478 485828 158484 485830
rect 158548 485828 158595 485832
rect 161054 485828 161060 485892
rect 161124 485890 161130 485892
rect 200849 485890 200915 485893
rect 161124 485888 200915 485890
rect 161124 485832 200854 485888
rect 200910 485832 200915 485888
rect 161124 485830 200915 485832
rect 161124 485828 161130 485830
rect 158529 485827 158595 485828
rect 200849 485827 200915 485830
rect 219249 485890 219315 485893
rect 253381 485892 253447 485893
rect 258349 485892 258415 485893
rect 266077 485892 266143 485893
rect 278405 485892 278471 485893
rect 310973 485892 311039 485893
rect 313549 485892 313615 485893
rect 251030 485890 251036 485892
rect 219249 485888 251036 485890
rect 219249 485832 219254 485888
rect 219310 485832 251036 485888
rect 219249 485830 251036 485832
rect 219249 485827 219315 485830
rect 251030 485828 251036 485830
rect 251100 485828 251106 485892
rect 253381 485888 253428 485892
rect 253492 485890 253498 485892
rect 253381 485832 253386 485888
rect 253381 485828 253428 485832
rect 253492 485830 253538 485890
rect 258349 485888 258396 485892
rect 258460 485890 258466 485892
rect 258349 485832 258354 485888
rect 253492 485828 253498 485830
rect 258349 485828 258396 485832
rect 258460 485830 258506 485890
rect 266077 485888 266124 485892
rect 266188 485890 266194 485892
rect 266077 485832 266082 485888
rect 258460 485828 258466 485830
rect 266077 485828 266124 485832
rect 266188 485830 266234 485890
rect 278405 485888 278452 485892
rect 278516 485890 278522 485892
rect 278405 485832 278410 485888
rect 266188 485828 266194 485830
rect 278405 485828 278452 485832
rect 278516 485830 278562 485890
rect 310973 485888 311020 485892
rect 311084 485890 311090 485892
rect 310973 485832 310978 485888
rect 278516 485828 278522 485830
rect 310973 485828 311020 485832
rect 311084 485830 311130 485890
rect 313549 485888 313596 485892
rect 313660 485890 313666 485892
rect 320265 485890 320331 485893
rect 320950 485890 320956 485892
rect 313549 485832 313554 485888
rect 311084 485828 311090 485830
rect 313549 485828 313596 485832
rect 313660 485830 313706 485890
rect 320265 485888 320956 485890
rect 320265 485832 320270 485888
rect 320326 485832 320956 485888
rect 320265 485830 320956 485832
rect 313660 485828 313666 485830
rect 253381 485827 253447 485828
rect 258349 485827 258415 485828
rect 266077 485827 266143 485828
rect 278405 485827 278471 485828
rect 310973 485827 311039 485828
rect 313549 485827 313615 485828
rect 320265 485827 320331 485830
rect 320950 485828 320956 485830
rect 321020 485828 321026 485892
rect 54845 485618 54911 485621
rect 126094 485618 126100 485620
rect 54845 485616 126100 485618
rect 54845 485560 54850 485616
rect 54906 485560 126100 485616
rect 54845 485558 126100 485560
rect 54845 485555 54911 485558
rect 126094 485556 126100 485558
rect 126164 485556 126170 485620
rect 96286 485420 96292 485484
rect 96356 485482 96362 485484
rect 197445 485482 197511 485485
rect 96356 485480 197511 485482
rect 96356 485424 197450 485480
rect 197506 485424 197511 485480
rect 96356 485422 197511 485424
rect 96356 485420 96362 485422
rect 197445 485419 197511 485422
rect 58433 485346 58499 485349
rect 88333 485346 88399 485349
rect 58433 485344 88399 485346
rect 58433 485288 58438 485344
rect 58494 485288 88338 485344
rect 88394 485288 88399 485344
rect 58433 485286 88399 485288
rect 58433 485283 58499 485286
rect 88333 485283 88399 485286
rect 156086 485284 156092 485348
rect 156156 485346 156162 485348
rect 213913 485346 213979 485349
rect 156156 485344 213979 485346
rect 156156 485288 213918 485344
rect 213974 485288 213979 485344
rect 156156 485286 213979 485288
rect 156156 485284 156162 485286
rect 213913 485283 213979 485286
rect 219157 485346 219223 485349
rect 273253 485346 273319 485349
rect 219157 485344 273319 485346
rect 219157 485288 219162 485344
rect 219218 485288 273258 485344
rect 273314 485288 273319 485344
rect 219157 485286 273319 485288
rect 219157 485283 219223 485286
rect 273253 485283 273319 485286
rect 58525 485210 58591 485213
rect 104893 485210 104959 485213
rect 58525 485208 104959 485210
rect 58525 485152 58530 485208
rect 58586 485152 104898 485208
rect 104954 485152 104959 485208
rect 58525 485150 104959 485152
rect 58525 485147 58591 485150
rect 104893 485147 104959 485150
rect 148358 485148 148364 485212
rect 148428 485210 148434 485212
rect 211153 485210 211219 485213
rect 148428 485208 211219 485210
rect 148428 485152 211158 485208
rect 211214 485152 211219 485208
rect 148428 485150 211219 485152
rect 148428 485148 148434 485150
rect 211153 485147 211219 485150
rect 219709 485210 219775 485213
rect 285990 485210 285996 485212
rect 219709 485208 285996 485210
rect 219709 485152 219714 485208
rect 219770 485152 285996 485208
rect 219709 485150 285996 485152
rect 219709 485147 219775 485150
rect 285990 485148 285996 485150
rect 286060 485148 286066 485212
rect 123702 485012 123708 485076
rect 123772 485074 123778 485076
rect 196801 485074 196867 485077
rect 123772 485072 196867 485074
rect 123772 485016 196806 485072
rect 196862 485016 196867 485072
rect 123772 485014 196867 485016
rect 123772 485012 123778 485014
rect 196801 485011 196867 485014
rect 200757 485074 200823 485077
rect 276054 485074 276060 485076
rect 200757 485072 276060 485074
rect 200757 485016 200762 485072
rect 200818 485016 276060 485072
rect 200757 485014 276060 485016
rect 200757 485011 200823 485014
rect 276054 485012 276060 485014
rect 276124 485012 276130 485076
rect 113582 484876 113588 484940
rect 113652 484938 113658 484940
rect 196709 484938 196775 484941
rect 113652 484936 196775 484938
rect 113652 484880 196714 484936
rect 196770 484880 196775 484936
rect 113652 484878 196775 484880
rect 113652 484876 113658 484878
rect 196709 484875 196775 484878
rect 198641 484938 198707 484941
rect 293534 484938 293540 484940
rect 198641 484936 293540 484938
rect 198641 484880 198646 484936
rect 198702 484880 293540 484936
rect 198641 484878 293540 484880
rect 198641 484875 198707 484878
rect 293534 484876 293540 484878
rect 293604 484876 293610 484940
rect 55121 484802 55187 484805
rect 88742 484802 88748 484804
rect 55121 484800 88748 484802
rect 55121 484744 55126 484800
rect 55182 484744 88748 484800
rect 55121 484742 88748 484744
rect 55121 484739 55187 484742
rect 88742 484740 88748 484742
rect 88812 484740 88818 484804
rect 103646 484740 103652 484804
rect 103716 484802 103722 484804
rect 197353 484802 197419 484805
rect 103716 484800 197419 484802
rect 103716 484744 197358 484800
rect 197414 484744 197419 484800
rect 103716 484742 197419 484744
rect 103716 484740 103722 484742
rect 197353 484739 197419 484742
rect 209681 484802 209747 484805
rect 305862 484802 305868 484804
rect 209681 484800 305868 484802
rect 209681 484744 209686 484800
rect 209742 484744 305868 484800
rect 209681 484742 305868 484744
rect 209681 484739 209747 484742
rect 305862 484740 305868 484742
rect 305932 484740 305938 484804
rect 58985 484666 59051 484669
rect 271086 484666 271092 484668
rect 58985 484664 271092 484666
rect 58985 484608 58990 484664
rect 59046 484608 271092 484664
rect 58985 484606 271092 484608
rect 58985 484603 59051 484606
rect 271086 484604 271092 484606
rect 271156 484604 271162 484668
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 55029 484530 55095 484533
rect 106038 484530 106044 484532
rect 55029 484528 106044 484530
rect 55029 484472 55034 484528
rect 55090 484472 106044 484528
rect 55029 484470 106044 484472
rect 55029 484467 55095 484470
rect 106038 484468 106044 484470
rect 106108 484468 106114 484532
rect 190862 484468 190868 484532
rect 190932 484530 190938 484532
rect 214557 484530 214623 484533
rect 190932 484528 214623 484530
rect 190932 484472 214562 484528
rect 214618 484472 214623 484528
rect 190932 484470 214623 484472
rect 190932 484468 190938 484470
rect 214557 484467 214623 484470
rect 215201 484530 215267 484533
rect 315798 484530 315804 484532
rect 215201 484528 315804 484530
rect 215201 484472 215206 484528
rect 215262 484472 315804 484528
rect 215201 484470 315804 484472
rect 215201 484467 215267 484470
rect 315798 484468 315804 484470
rect 315868 484468 315874 484532
rect 338430 484468 338436 484532
rect 338500 484530 338506 484532
rect 356513 484530 356579 484533
rect 338500 484528 356579 484530
rect 338500 484472 356518 484528
rect 356574 484472 356579 484528
rect 583520 484516 584960 484606
rect 338500 484470 356579 484472
rect 338500 484468 338506 484470
rect 356513 484467 356579 484470
rect 116158 484196 116164 484260
rect 116228 484258 116234 484260
rect 218513 484258 218579 484261
rect 116228 484256 218579 484258
rect 116228 484200 218518 484256
rect 218574 484200 218579 484256
rect 116228 484198 218579 484200
rect 116228 484196 116234 484198
rect 218513 484195 218579 484198
rect 179638 484060 179644 484124
rect 179708 484122 179714 484124
rect 197629 484122 197695 484125
rect 179708 484120 197695 484122
rect 179708 484064 197634 484120
rect 197690 484064 197695 484120
rect 179708 484062 197695 484064
rect 179708 484060 179714 484062
rect 197629 484059 197695 484062
rect 57513 483986 57579 483989
rect 166022 483986 166028 483988
rect 57513 483984 166028 483986
rect 57513 483928 57518 483984
rect 57574 483928 166028 483984
rect 57513 483926 166028 483928
rect 57513 483923 57579 483926
rect 166022 483924 166028 483926
rect 166092 483924 166098 483988
rect 178534 483924 178540 483988
rect 178604 483986 178610 483988
rect 197537 483986 197603 483989
rect 178604 483984 197603 483986
rect 178604 483928 197542 483984
rect 197598 483928 197603 483984
rect 178604 483926 197603 483928
rect 178604 483924 178610 483926
rect 197537 483923 197603 483926
rect 219525 483986 219591 483989
rect 248638 483986 248644 483988
rect 219525 483984 248644 483986
rect 219525 483928 219530 483984
rect 219586 483928 248644 483984
rect 219525 483926 248644 483928
rect 219525 483923 219591 483926
rect 248638 483924 248644 483926
rect 248708 483924 248714 483988
rect 218053 483850 218119 483853
rect 303470 483850 303476 483852
rect 218053 483848 303476 483850
rect 218053 483792 218058 483848
rect 218114 483792 303476 483848
rect 218053 483790 303476 483792
rect 218053 483787 218119 483790
rect 303470 483788 303476 483790
rect 303540 483788 303546 483852
rect 163360 483652 163366 483716
rect 163430 483714 163436 483716
rect 216213 483714 216279 483717
rect 163430 483712 216279 483714
rect 163430 483656 216218 483712
rect 216274 483656 216279 483712
rect 163430 483654 216279 483656
rect 163430 483652 163436 483654
rect 216213 483651 216279 483654
rect 219617 483714 219683 483717
rect 308400 483714 308406 483716
rect 219617 483712 308406 483714
rect 219617 483656 219622 483712
rect 219678 483656 308406 483712
rect 219617 483654 308406 483656
rect 219617 483651 219683 483654
rect 308400 483652 308406 483654
rect 308470 483652 308476 483716
rect 108552 483516 108558 483580
rect 108622 483578 108628 483580
rect 218329 483578 218395 483581
rect 108622 483576 218395 483578
rect 108622 483520 218334 483576
rect 218390 483520 218395 483576
rect 108622 483518 218395 483520
rect 108622 483516 108628 483518
rect 218329 483515 218395 483518
rect 219065 483578 219131 483581
rect 326080 483578 326086 483580
rect 219065 483576 326086 483578
rect 219065 483520 219070 483576
rect 219126 483520 326086 483576
rect 219065 483518 326086 483520
rect 219065 483515 219131 483518
rect 326080 483516 326086 483518
rect 326150 483516 326156 483580
rect 53557 483442 53623 483445
rect 280928 483442 280934 483444
rect 53557 483440 280934 483442
rect 53557 483384 53562 483440
rect 53618 483384 280934 483440
rect 53557 483382 280934 483384
rect 53557 483379 53623 483382
rect 280928 483380 280934 483382
rect 280998 483380 281004 483444
rect 298608 483380 298614 483444
rect 298678 483380 298684 483444
rect 53373 483306 53439 483309
rect 298616 483306 298676 483380
rect 53373 483304 298676 483306
rect 53373 483248 53378 483304
rect 53434 483248 298676 483304
rect 53373 483246 298676 483248
rect 53373 483243 53439 483246
rect 199377 479226 199443 479229
rect 197126 479224 199443 479226
rect 197126 479220 199382 479224
rect 196604 479168 199382 479220
rect 199438 479168 199443 479224
rect 196604 479166 199443 479168
rect 196604 479160 197186 479166
rect 199377 479163 199443 479166
rect 356562 478954 356622 479190
rect 358997 478954 359063 478957
rect 356562 478952 359063 478954
rect 356562 478896 359002 478952
rect 359058 478896 359063 478952
rect 356562 478894 359063 478896
rect 358997 478891 359063 478894
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect 217501 436930 217567 436933
rect 217501 436928 219450 436930
rect -960 436508 480 436748
rect 57789 436386 57855 436389
rect 60002 436386 60062 436894
rect 217501 436872 217506 436928
rect 217562 436924 219450 436928
rect 217562 436872 220064 436924
rect 217501 436870 220064 436872
rect 217501 436867 217567 436870
rect 219390 436864 220064 436870
rect 57789 436384 60062 436386
rect 57789 436328 57794 436384
rect 57850 436328 60062 436384
rect 57789 436326 60062 436328
rect 57789 436323 57855 436326
rect 217685 435978 217751 435981
rect 217685 435976 219450 435978
rect 57329 435434 57395 435437
rect 60002 435434 60062 435942
rect 217685 435920 217690 435976
rect 217746 435972 219450 435976
rect 217746 435920 220064 435972
rect 217685 435918 220064 435920
rect 217685 435915 217751 435918
rect 219390 435912 220064 435918
rect 57329 435432 60062 435434
rect 57329 435376 57334 435432
rect 57390 435376 60062 435432
rect 57329 435374 60062 435376
rect 57329 435371 57395 435374
rect 217777 433802 217843 433805
rect 217777 433800 219450 433802
rect 57237 433394 57303 433397
rect 60002 433394 60062 433766
rect 217777 433744 217782 433800
rect 217838 433796 219450 433800
rect 217838 433744 220064 433796
rect 217777 433742 220064 433744
rect 217777 433739 217843 433742
rect 219390 433736 220064 433742
rect 57237 433392 60062 433394
rect 57237 433336 57242 433392
rect 57298 433336 60062 433392
rect 57237 433334 60062 433336
rect 57237 433331 57303 433334
rect 217869 432850 217935 432853
rect 217869 432848 219450 432850
rect 56593 432306 56659 432309
rect 60002 432306 60062 432814
rect 217869 432792 217874 432848
rect 217930 432844 219450 432848
rect 217930 432792 220064 432844
rect 217869 432790 220064 432792
rect 217869 432787 217935 432790
rect 219390 432784 220064 432790
rect 56593 432304 60062 432306
rect 56593 432248 56598 432304
rect 56654 432248 60062 432304
rect 56593 432246 60062 432248
rect 56593 432243 56659 432246
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 216673 431082 216739 431085
rect 216673 431080 219450 431082
rect 57605 430674 57671 430677
rect 60002 430674 60062 431046
rect 216673 431024 216678 431080
rect 216734 431076 219450 431080
rect 216734 431024 220064 431076
rect 216673 431022 220064 431024
rect 216673 431019 216739 431022
rect 219390 431016 220064 431022
rect 57605 430672 60062 430674
rect 57605 430616 57610 430672
rect 57666 430616 60062 430672
rect 57605 430614 60062 430616
rect 57605 430611 57671 430614
rect 217409 429994 217475 429997
rect 217409 429992 219450 429994
rect 57145 429450 57211 429453
rect 60002 429450 60062 429958
rect 217409 429936 217414 429992
rect 217470 429988 219450 429992
rect 217470 429936 220064 429988
rect 217409 429934 220064 429936
rect 217409 429931 217475 429934
rect 219390 429928 220064 429934
rect 57145 429448 60062 429450
rect 57145 429392 57150 429448
rect 57206 429392 60062 429448
rect 57145 429390 60062 429392
rect 57145 429387 57211 429390
rect 217593 428226 217659 428229
rect 217593 428224 219450 428226
rect 57421 427954 57487 427957
rect 60002 427954 60062 428190
rect 217593 428168 217598 428224
rect 217654 428220 219450 428224
rect 217654 428168 220064 428220
rect 217593 428166 220064 428168
rect 217593 428163 217659 428166
rect 219390 428160 220064 428166
rect 57421 427952 60062 427954
rect 57421 427896 57426 427952
rect 57482 427896 60062 427952
rect 57421 427894 60062 427896
rect 57421 427891 57487 427894
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 199653 419386 199719 419389
rect 197126 419384 199719 419386
rect 197126 419380 199658 419384
rect 196604 419328 199658 419380
rect 199714 419328 199719 419384
rect 196604 419326 199719 419328
rect 196604 419320 197186 419326
rect 199653 419323 199719 419326
rect 356562 418842 356622 419350
rect 357433 418842 357499 418845
rect 356562 418840 357499 418842
rect 356562 418784 357438 418840
rect 357494 418784 357499 418840
rect 356562 418782 357499 418784
rect 357433 418779 357499 418782
rect 580257 418298 580323 418301
rect 583520 418298 584960 418388
rect 580257 418296 584960 418298
rect 580257 418240 580262 418296
rect 580318 418240 584960 418296
rect 580257 418238 584960 418240
rect 580257 418235 580323 418238
rect 583520 418148 584960 418238
rect 197721 417754 197787 417757
rect 197126 417752 197787 417754
rect 197126 417748 197726 417752
rect 196604 417696 197726 417748
rect 197782 417696 197787 417752
rect 196604 417694 197787 417696
rect 196604 417688 197186 417694
rect 197721 417691 197787 417694
rect 356562 417210 356622 417718
rect 359089 417210 359155 417213
rect 356562 417208 359155 417210
rect 356562 417152 359094 417208
rect 359150 417152 359155 417208
rect 356562 417150 359155 417152
rect 359089 417147 359155 417150
rect 198733 416394 198799 416397
rect 197126 416392 198799 416394
rect 197126 416388 198738 416392
rect 196604 416336 198738 416388
rect 198794 416336 198799 416392
rect 196604 416334 198799 416336
rect 196604 416328 197186 416334
rect 198733 416331 198799 416334
rect 356562 415850 356622 416358
rect 358813 415850 358879 415853
rect 356562 415848 358879 415850
rect 356562 415792 358818 415848
rect 358874 415792 358879 415848
rect 356562 415790 358879 415792
rect 358813 415787 358879 415790
rect 199469 414898 199535 414901
rect 197126 414896 199535 414898
rect 197126 414892 199474 414896
rect 196604 414840 199474 414892
rect 199530 414840 199535 414896
rect 196604 414838 199535 414840
rect 196604 414832 197186 414838
rect 199469 414835 199535 414838
rect 356562 414354 356622 414862
rect 357525 414354 357591 414357
rect 356562 414352 357591 414354
rect 356562 414296 357530 414352
rect 357586 414296 357591 414352
rect 356562 414294 357591 414296
rect 357525 414291 357591 414294
rect 199561 413674 199627 413677
rect 197126 413672 199627 413674
rect 197126 413668 199566 413672
rect 196604 413616 199566 413668
rect 199622 413616 199627 413672
rect 196604 413614 199627 413616
rect 196604 413608 197186 413614
rect 199561 413611 199627 413614
rect 356562 413130 356622 413638
rect 358905 413130 358971 413133
rect 356562 413128 358971 413130
rect 356562 413072 358910 413128
rect 358966 413072 358971 413128
rect 356562 413070 358971 413072
rect 358905 413067 358971 413070
rect -960 410546 480 410636
rect 3417 410546 3483 410549
rect -960 410544 3483 410546
rect -960 410488 3422 410544
rect 3478 410488 3483 410544
rect -960 410486 3483 410488
rect -960 410396 480 410486
rect 3417 410483 3483 410486
rect 57881 410002 57947 410005
rect 217225 410002 217291 410005
rect 57881 410000 60062 410002
rect 57881 409944 57886 410000
rect 57942 409944 60062 410000
rect 57881 409942 60062 409944
rect 217225 410000 219450 410002
rect 217225 409944 217230 410000
rect 217286 409996 219450 410000
rect 217286 409944 220064 409996
rect 217225 409942 220064 409944
rect 57881 409939 57947 409942
rect 217225 409939 217291 409942
rect 219390 409936 220064 409942
rect 216673 408370 216739 408373
rect 216673 408368 219450 408370
rect 59353 408234 59419 408237
rect 60002 408234 60062 408334
rect 216673 408312 216678 408368
rect 216734 408364 219450 408368
rect 216734 408312 220064 408364
rect 216673 408310 220064 408312
rect 216673 408307 216739 408310
rect 219390 408304 220064 408310
rect 59353 408232 60062 408234
rect 59353 408176 59358 408232
rect 59414 408176 60062 408232
rect 59353 408174 60062 408176
rect 59353 408171 59419 408174
rect 217133 408098 217199 408101
rect 217133 408096 220094 408098
rect 57053 407554 57119 407557
rect 60002 407554 60062 408062
rect 217133 408040 217138 408096
rect 217194 408040 220094 408096
rect 217133 408038 220094 408040
rect 217133 408035 217199 408038
rect 57053 407552 60062 407554
rect 57053 407496 57058 407552
rect 57114 407496 60062 407552
rect 57053 407494 60062 407496
rect 57053 407491 57119 407494
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 85481 398172 85547 398173
rect 85430 398170 85436 398172
rect 85390 398110 85436 398170
rect 85500 398168 85547 398172
rect 85542 398112 85547 398168
rect 85430 398108 85436 398110
rect 85500 398108 85547 398112
rect 85481 398107 85547 398108
rect 92289 398170 92355 398173
rect 95877 398172 95943 398173
rect 113633 398172 113699 398173
rect 92422 398170 92428 398172
rect 92289 398168 92428 398170
rect 92289 398112 92294 398168
rect 92350 398112 92428 398168
rect 92289 398110 92428 398112
rect 92289 398107 92355 398110
rect 92422 398108 92428 398110
rect 92492 398108 92498 398172
rect 95877 398168 95924 398172
rect 95988 398170 95994 398172
rect 113582 398170 113588 398172
rect 95877 398112 95882 398168
rect 95877 398108 95924 398112
rect 95988 398110 96034 398170
rect 113542 398110 113588 398170
rect 113652 398168 113699 398172
rect 113694 398112 113699 398168
rect 95988 398108 95994 398110
rect 113582 398108 113588 398110
rect 113652 398108 113699 398112
rect 95877 398107 95943 398108
rect 113633 398107 113699 398108
rect 218789 398170 218855 398173
rect 219801 398170 219867 398173
rect 235993 398172 236059 398173
rect 223798 398170 223804 398172
rect 218789 398168 219634 398170
rect 218789 398112 218794 398168
rect 218850 398112 219634 398168
rect 218789 398110 219634 398112
rect 218789 398107 218855 398110
rect 218973 398034 219039 398037
rect 219574 398034 219634 398110
rect 219801 398168 223804 398170
rect 219801 398112 219806 398168
rect 219862 398112 223804 398168
rect 219801 398110 223804 398112
rect 219801 398107 219867 398110
rect 223798 398108 223804 398110
rect 223868 398108 223874 398172
rect 235942 398170 235948 398172
rect 235902 398110 235948 398170
rect 236012 398168 236059 398172
rect 236054 398112 236059 398168
rect 235942 398108 235948 398110
rect 236012 398108 236059 398112
rect 235993 398107 236059 398108
rect 265065 398170 265131 398173
rect 265198 398170 265204 398172
rect 265065 398168 265204 398170
rect 265065 398112 265070 398168
rect 265126 398112 265204 398168
rect 265065 398110 265204 398112
rect 265065 398107 265131 398110
rect 265198 398108 265204 398110
rect 265268 398108 265274 398172
rect 300117 398170 300183 398173
rect 315757 398172 315823 398173
rect 325877 398172 325943 398173
rect 300894 398170 300900 398172
rect 300117 398168 300900 398170
rect 300117 398112 300122 398168
rect 300178 398112 300900 398168
rect 300117 398110 300900 398112
rect 300117 398107 300183 398110
rect 300894 398108 300900 398110
rect 300964 398108 300970 398172
rect 315757 398168 315804 398172
rect 315868 398170 315874 398172
rect 315757 398112 315762 398168
rect 315757 398108 315804 398112
rect 315868 398110 315914 398170
rect 325877 398168 325924 398172
rect 325988 398170 325994 398172
rect 325877 398112 325882 398168
rect 315868 398108 315874 398110
rect 325877 398108 325924 398112
rect 325988 398110 326034 398170
rect 325988 398108 325994 398110
rect 315757 398107 315823 398108
rect 325877 398107 325943 398108
rect 223614 398034 223620 398036
rect 218973 398032 219450 398034
rect 218973 397976 218978 398032
rect 219034 397976 219450 398032
rect 218973 397974 219450 397976
rect 219574 397974 223620 398034
rect 218973 397971 219039 397974
rect 219390 397898 219450 397974
rect 223614 397972 223620 397974
rect 223684 397972 223690 398036
rect 224902 397898 224908 397900
rect 219390 397838 224908 397898
rect 224902 397836 224908 397838
rect 224972 397836 224978 397900
rect -960 397490 480 397580
rect 3509 397490 3575 397493
rect -960 397488 3575 397490
rect -960 397432 3514 397488
rect 3570 397432 3575 397488
rect -960 397430 3575 397432
rect -960 397340 480 397430
rect 3509 397427 3575 397430
rect 76189 397354 76255 397357
rect 78305 397356 78371 397357
rect 79593 397356 79659 397357
rect 77150 397354 77156 397356
rect 76189 397352 77156 397354
rect 76189 397296 76194 397352
rect 76250 397296 77156 397352
rect 76189 397294 77156 397296
rect 76189 397291 76255 397294
rect 77150 397292 77156 397294
rect 77220 397292 77226 397356
rect 78254 397354 78260 397356
rect 78214 397294 78260 397354
rect 78324 397352 78371 397356
rect 79542 397354 79548 397356
rect 78366 397296 78371 397352
rect 78254 397292 78260 397294
rect 78324 397292 78371 397296
rect 79502 397294 79548 397354
rect 79612 397352 79659 397356
rect 79654 397296 79659 397352
rect 79542 397292 79548 397294
rect 79612 397292 79659 397296
rect 78305 397291 78371 397292
rect 79593 397291 79659 397292
rect 80421 397356 80487 397357
rect 80421 397352 80468 397356
rect 80532 397354 80538 397356
rect 80421 397296 80426 397352
rect 80421 397292 80468 397296
rect 80532 397294 80578 397354
rect 80532 397292 80538 397294
rect 81934 397292 81940 397356
rect 82004 397354 82010 397356
rect 82353 397354 82419 397357
rect 82004 397352 82419 397354
rect 82004 397296 82358 397352
rect 82414 397296 82419 397352
rect 82004 397294 82419 397296
rect 82004 397292 82010 397294
rect 80421 397291 80487 397292
rect 82353 397291 82419 397294
rect 82997 397356 83063 397357
rect 82997 397352 83044 397356
rect 83108 397354 83114 397356
rect 82997 397296 83002 397352
rect 82997 397292 83044 397296
rect 83108 397294 83154 397354
rect 83108 397292 83114 397294
rect 88742 397292 88748 397356
rect 88812 397354 88818 397356
rect 89345 397354 89411 397357
rect 90081 397356 90147 397357
rect 90030 397354 90036 397356
rect 88812 397352 89411 397354
rect 88812 397296 89350 397352
rect 89406 397296 89411 397352
rect 88812 397294 89411 397296
rect 89990 397294 90036 397354
rect 90100 397352 90147 397356
rect 90142 397296 90147 397352
rect 88812 397292 88818 397294
rect 82997 397291 83063 397292
rect 89345 397291 89411 397294
rect 90030 397292 90036 397294
rect 90100 397292 90147 397296
rect 91318 397292 91324 397356
rect 91388 397354 91394 397356
rect 91461 397354 91527 397357
rect 91388 397352 91527 397354
rect 91388 397296 91466 397352
rect 91522 397296 91527 397352
rect 91388 397294 91527 397296
rect 91388 397292 91394 397294
rect 90081 397291 90147 397292
rect 91461 397291 91527 397294
rect 93342 397292 93348 397356
rect 93412 397354 93418 397356
rect 93485 397354 93551 397357
rect 93412 397352 93551 397354
rect 93412 397296 93490 397352
rect 93546 397296 93551 397352
rect 93412 397294 93551 397296
rect 93412 397292 93418 397294
rect 93485 397291 93551 397294
rect 94630 397292 94636 397356
rect 94700 397354 94706 397356
rect 95049 397354 95115 397357
rect 94700 397352 95115 397354
rect 94700 397296 95054 397352
rect 95110 397296 95115 397352
rect 94700 397294 95115 397296
rect 94700 397292 94706 397294
rect 95049 397291 95115 397294
rect 98085 397356 98151 397357
rect 102777 397356 102843 397357
rect 98085 397352 98132 397356
rect 98196 397354 98202 397356
rect 102726 397354 102732 397356
rect 98085 397296 98090 397352
rect 98085 397292 98132 397296
rect 98196 397294 98242 397354
rect 102686 397294 102732 397354
rect 102796 397352 102843 397356
rect 102838 397296 102843 397352
rect 98196 397292 98202 397294
rect 102726 397292 102732 397294
rect 102796 397292 102843 397296
rect 104014 397292 104020 397356
rect 104084 397354 104090 397356
rect 104801 397354 104867 397357
rect 104084 397352 104867 397354
rect 104084 397296 104806 397352
rect 104862 397296 104867 397352
rect 104084 397294 104867 397296
rect 104084 397292 104090 397294
rect 98085 397291 98151 397292
rect 102777 397291 102843 397292
rect 104801 397291 104867 397294
rect 105302 397292 105308 397356
rect 105372 397354 105378 397356
rect 106089 397354 106155 397357
rect 105372 397352 106155 397354
rect 105372 397296 106094 397352
rect 106150 397296 106155 397352
rect 105372 397294 106155 397296
rect 105372 397292 105378 397294
rect 106089 397291 106155 397294
rect 106406 397292 106412 397356
rect 106476 397354 106482 397356
rect 106917 397354 106983 397357
rect 108849 397356 108915 397357
rect 108798 397354 108804 397356
rect 106476 397352 106983 397354
rect 106476 397296 106922 397352
rect 106978 397296 106983 397352
rect 106476 397294 106983 397296
rect 108758 397294 108804 397354
rect 108868 397352 108915 397356
rect 108910 397296 108915 397352
rect 106476 397292 106482 397294
rect 106917 397291 106983 397294
rect 108798 397292 108804 397294
rect 108868 397292 108915 397296
rect 108849 397291 108915 397292
rect 109125 397354 109191 397357
rect 112345 397356 112411 397357
rect 109534 397354 109540 397356
rect 109125 397352 109540 397354
rect 109125 397296 109130 397352
rect 109186 397296 109540 397352
rect 109125 397294 109540 397296
rect 109125 397291 109191 397294
rect 109534 397292 109540 397294
rect 109604 397292 109610 397356
rect 112294 397354 112300 397356
rect 112254 397294 112300 397354
rect 112364 397352 112411 397356
rect 112406 397296 112411 397352
rect 112294 397292 112300 397294
rect 112364 397292 112411 397296
rect 113214 397292 113220 397356
rect 113284 397354 113290 397356
rect 113357 397354 113423 397357
rect 113284 397352 113423 397354
rect 113284 397296 113362 397352
rect 113418 397296 113423 397352
rect 113284 397294 113423 397296
rect 113284 397292 113290 397294
rect 112345 397291 112411 397292
rect 113357 397291 113423 397294
rect 113817 397354 113883 397357
rect 118233 397356 118299 397357
rect 118601 397356 118667 397357
rect 114318 397354 114324 397356
rect 113817 397352 114324 397354
rect 113817 397296 113822 397352
rect 113878 397296 114324 397352
rect 113817 397294 114324 397296
rect 113817 397291 113883 397294
rect 114318 397292 114324 397294
rect 114388 397292 114394 397356
rect 118182 397354 118188 397356
rect 118142 397294 118188 397354
rect 118252 397352 118299 397356
rect 118550 397354 118556 397356
rect 118294 397296 118299 397352
rect 118182 397292 118188 397294
rect 118252 397292 118299 397296
rect 118510 397294 118556 397354
rect 118620 397352 118667 397356
rect 118662 397296 118667 397352
rect 118550 397292 118556 397294
rect 118620 397292 118667 397296
rect 136030 397292 136036 397356
rect 136100 397354 136106 397356
rect 136449 397354 136515 397357
rect 154113 397356 154179 397357
rect 154062 397354 154068 397356
rect 136100 397352 136515 397354
rect 136100 397296 136454 397352
rect 136510 397296 136515 397352
rect 136100 397294 136515 397296
rect 154022 397294 154068 397354
rect 154132 397352 154179 397356
rect 154174 397296 154179 397352
rect 136100 397292 136106 397294
rect 118233 397291 118299 397292
rect 118601 397291 118667 397292
rect 136449 397291 136515 397294
rect 154062 397292 154068 397294
rect 154132 397292 154179 397296
rect 163446 397292 163452 397356
rect 163516 397354 163522 397356
rect 163865 397354 163931 397357
rect 163516 397352 163931 397354
rect 163516 397296 163870 397352
rect 163926 397296 163931 397352
rect 163516 397294 163931 397296
rect 163516 397292 163522 397294
rect 154113 397291 154179 397292
rect 163865 397291 163931 397294
rect 183461 397356 183527 397357
rect 183461 397352 183508 397356
rect 183572 397354 183578 397356
rect 236177 397354 236243 397357
rect 239213 397356 239279 397357
rect 247677 397356 247743 397357
rect 237046 397354 237052 397356
rect 183461 397296 183466 397352
rect 183461 397292 183508 397296
rect 183572 397294 183618 397354
rect 236177 397352 237052 397354
rect 236177 397296 236182 397352
rect 236238 397296 237052 397352
rect 236177 397294 237052 397296
rect 183572 397292 183578 397294
rect 183461 397291 183527 397292
rect 236177 397291 236243 397294
rect 237046 397292 237052 397294
rect 237116 397292 237122 397356
rect 239213 397352 239260 397356
rect 239324 397354 239330 397356
rect 239213 397296 239218 397352
rect 239213 397292 239260 397296
rect 239324 397294 239370 397354
rect 247677 397352 247724 397356
rect 247788 397354 247794 397356
rect 247953 397354 248019 397357
rect 248597 397356 248663 397357
rect 250069 397356 250135 397357
rect 248270 397354 248276 397356
rect 247677 397296 247682 397352
rect 239324 397292 239330 397294
rect 247677 397292 247724 397296
rect 247788 397294 247834 397354
rect 247953 397352 248276 397354
rect 247953 397296 247958 397352
rect 248014 397296 248276 397352
rect 247953 397294 248276 397296
rect 247788 397292 247794 397294
rect 239213 397291 239279 397292
rect 247677 397291 247743 397292
rect 247953 397291 248019 397294
rect 248270 397292 248276 397294
rect 248340 397292 248346 397356
rect 248597 397352 248644 397356
rect 248708 397354 248714 397356
rect 248597 397296 248602 397352
rect 248597 397292 248644 397296
rect 248708 397294 248754 397354
rect 250069 397352 250116 397356
rect 250180 397354 250186 397356
rect 250345 397354 250411 397357
rect 250662 397354 250668 397356
rect 250069 397296 250074 397352
rect 248708 397292 248714 397294
rect 250069 397292 250116 397296
rect 250180 397294 250226 397354
rect 250345 397352 250668 397354
rect 250345 397296 250350 397352
rect 250406 397296 250668 397352
rect 250345 397294 250668 397296
rect 250180 397292 250186 397294
rect 248597 397291 248663 397292
rect 250069 397291 250135 397292
rect 250345 397291 250411 397294
rect 250662 397292 250668 397294
rect 250732 397292 250738 397356
rect 252737 397354 252803 397357
rect 259453 397356 259519 397357
rect 260925 397356 260991 397357
rect 253422 397354 253428 397356
rect 252737 397352 253428 397354
rect 252737 397296 252742 397352
rect 252798 397296 253428 397352
rect 252737 397294 253428 397296
rect 252737 397291 252803 397294
rect 253422 397292 253428 397294
rect 253492 397292 253498 397356
rect 259453 397352 259500 397356
rect 259564 397354 259570 397356
rect 259453 397296 259458 397352
rect 259453 397292 259500 397296
rect 259564 397294 259610 397354
rect 260925 397352 260972 397356
rect 261036 397354 261042 397356
rect 261937 397354 262003 397357
rect 262070 397354 262076 397356
rect 260925 397296 260930 397352
rect 259564 397292 259570 397294
rect 260925 397292 260972 397296
rect 261036 397294 261082 397354
rect 261937 397352 262076 397354
rect 261937 397296 261942 397352
rect 261998 397296 262076 397352
rect 261937 397294 262076 397296
rect 261036 397292 261042 397294
rect 259453 397291 259519 397292
rect 260925 397291 260991 397292
rect 261937 397291 262003 397294
rect 262070 397292 262076 397294
rect 262140 397292 262146 397356
rect 262305 397354 262371 397357
rect 262806 397354 262812 397356
rect 262305 397352 262812 397354
rect 262305 397296 262310 397352
rect 262366 397296 262812 397352
rect 262305 397294 262812 397296
rect 262305 397291 262371 397294
rect 262806 397292 262812 397294
rect 262876 397292 262882 397356
rect 263593 397354 263659 397357
rect 268285 397356 268351 397357
rect 268653 397356 268719 397357
rect 263910 397354 263916 397356
rect 263593 397352 263916 397354
rect 263593 397296 263598 397352
rect 263654 397296 263916 397352
rect 263593 397294 263916 397296
rect 263593 397291 263659 397294
rect 263910 397292 263916 397294
rect 263980 397292 263986 397356
rect 268285 397352 268332 397356
rect 268396 397354 268402 397356
rect 268285 397296 268290 397352
rect 268285 397292 268332 397296
rect 268396 397294 268442 397354
rect 268653 397352 268700 397356
rect 268764 397354 268770 397356
rect 272333 397354 272399 397357
rect 275277 397356 275343 397357
rect 272558 397354 272564 397356
rect 268653 397296 268658 397352
rect 268396 397292 268402 397294
rect 268653 397292 268700 397296
rect 268764 397294 268810 397354
rect 272333 397352 272564 397354
rect 272333 397296 272338 397352
rect 272394 397296 272564 397352
rect 272333 397294 272564 397296
rect 268764 397292 268770 397294
rect 268285 397291 268351 397292
rect 268653 397291 268719 397292
rect 272333 397291 272399 397294
rect 272558 397292 272564 397294
rect 272628 397292 272634 397356
rect 275277 397352 275324 397356
rect 275388 397354 275394 397356
rect 277669 397354 277735 397357
rect 278078 397354 278084 397356
rect 275277 397296 275282 397352
rect 275277 397292 275324 397296
rect 275388 397294 275434 397354
rect 277669 397352 278084 397354
rect 277669 397296 277674 397352
rect 277730 397296 278084 397352
rect 277669 397294 278084 397296
rect 275388 397292 275394 397294
rect 275277 397291 275343 397292
rect 277669 397291 277735 397294
rect 278078 397292 278084 397294
rect 278148 397292 278154 397356
rect 278865 397354 278931 397357
rect 278998 397354 279004 397356
rect 278865 397352 279004 397354
rect 278865 397296 278870 397352
rect 278926 397296 279004 397352
rect 278865 397294 279004 397296
rect 278865 397291 278931 397294
rect 278998 397292 279004 397294
rect 279068 397292 279074 397356
rect 290181 397354 290247 397357
rect 298461 397356 298527 397357
rect 308581 397356 308647 397357
rect 290958 397354 290964 397356
rect 290181 397352 290964 397354
rect 290181 397296 290186 397352
rect 290242 397296 290964 397352
rect 290181 397294 290964 397296
rect 290181 397291 290247 397294
rect 290958 397292 290964 397294
rect 291028 397292 291034 397356
rect 298461 397352 298508 397356
rect 298572 397354 298578 397356
rect 298461 397296 298466 397352
rect 298461 397292 298508 397296
rect 298572 397294 298618 397354
rect 308581 397352 308628 397356
rect 308692 397354 308698 397356
rect 342621 397354 342687 397357
rect 343214 397354 343220 397356
rect 308581 397296 308586 397352
rect 298572 397292 298578 397294
rect 308581 397292 308628 397296
rect 308692 397294 308738 397354
rect 342621 397352 343220 397354
rect 342621 397296 342626 397352
rect 342682 397296 343220 397352
rect 342621 397294 343220 397296
rect 308692 397292 308698 397294
rect 298461 397291 298527 397292
rect 308581 397291 308647 397292
rect 342621 397291 342687 397294
rect 343214 397292 343220 397294
rect 343284 397292 343290 397356
rect 251173 397084 251239 397085
rect 251173 397080 251220 397084
rect 251284 397082 251290 397084
rect 251173 397024 251178 397080
rect 251173 397020 251220 397024
rect 251284 397022 251330 397082
rect 251284 397020 251290 397022
rect 251173 397019 251239 397020
rect 100702 396884 100708 396948
rect 100772 396946 100778 396948
rect 101949 396946 102015 396949
rect 100772 396944 102015 396946
rect 100772 396888 101954 396944
rect 102010 396888 102015 396944
rect 100772 396886 102015 396888
rect 100772 396884 100778 396886
rect 101949 396883 102015 396886
rect 258073 396946 258139 396949
rect 258390 396946 258396 396948
rect 258073 396944 258396 396946
rect 258073 396888 258078 396944
rect 258134 396888 258396 396944
rect 258073 396886 258396 396888
rect 258073 396883 258139 396886
rect 258390 396884 258396 396886
rect 258460 396884 258466 396948
rect 76046 396748 76052 396812
rect 76116 396810 76122 396812
rect 77201 396810 77267 396813
rect 76116 396808 77267 396810
rect 76116 396752 77206 396808
rect 77262 396752 77267 396808
rect 76116 396750 77267 396752
rect 76116 396748 76122 396750
rect 77201 396747 77267 396750
rect 84326 396748 84332 396812
rect 84396 396810 84402 396812
rect 85389 396810 85455 396813
rect 84396 396808 85455 396810
rect 84396 396752 85394 396808
rect 85450 396752 85455 396808
rect 84396 396750 85455 396752
rect 84396 396748 84402 396750
rect 85389 396747 85455 396750
rect 86534 396748 86540 396812
rect 86604 396810 86610 396812
rect 86861 396810 86927 396813
rect 86604 396808 86927 396810
rect 86604 396752 86866 396808
rect 86922 396752 86927 396808
rect 86604 396750 86927 396752
rect 86604 396748 86610 396750
rect 86861 396747 86927 396750
rect 87638 396748 87644 396812
rect 87708 396810 87714 396812
rect 88241 396810 88307 396813
rect 87708 396808 88307 396810
rect 87708 396752 88246 396808
rect 88302 396752 88307 396808
rect 87708 396750 88307 396752
rect 87708 396748 87714 396750
rect 88241 396747 88307 396750
rect 88374 396748 88380 396812
rect 88444 396810 88450 396812
rect 89529 396810 89595 396813
rect 88444 396808 89595 396810
rect 88444 396752 89534 396808
rect 89590 396752 89595 396808
rect 88444 396750 89595 396752
rect 88444 396748 88450 396750
rect 89529 396747 89595 396750
rect 90766 396748 90772 396812
rect 90836 396810 90842 396812
rect 90909 396810 90975 396813
rect 90836 396808 90975 396810
rect 90836 396752 90914 396808
rect 90970 396752 90975 396808
rect 90836 396750 90975 396752
rect 90836 396748 90842 396750
rect 90909 396747 90975 396750
rect 92473 396810 92539 396813
rect 93710 396810 93716 396812
rect 92473 396808 93716 396810
rect 92473 396752 92478 396808
rect 92534 396752 93716 396808
rect 92473 396750 93716 396752
rect 92473 396747 92539 396750
rect 93710 396748 93716 396750
rect 93780 396748 93786 396812
rect 96286 396748 96292 396812
rect 96356 396810 96362 396812
rect 96521 396810 96587 396813
rect 96356 396808 96587 396810
rect 96356 396752 96526 396808
rect 96582 396752 96587 396808
rect 96356 396750 96587 396752
rect 96356 396748 96362 396750
rect 96521 396747 96587 396750
rect 97022 396748 97028 396812
rect 97092 396810 97098 396812
rect 97901 396810 97967 396813
rect 97092 396808 97967 396810
rect 97092 396752 97906 396808
rect 97962 396752 97967 396808
rect 97092 396750 97967 396752
rect 97092 396748 97098 396750
rect 97901 396747 97967 396750
rect 98494 396748 98500 396812
rect 98564 396810 98570 396812
rect 99281 396810 99347 396813
rect 98564 396808 99347 396810
rect 98564 396752 99286 396808
rect 99342 396752 99347 396808
rect 98564 396750 99347 396752
rect 98564 396748 98570 396750
rect 99281 396747 99347 396750
rect 99966 396748 99972 396812
rect 100036 396810 100042 396812
rect 100661 396810 100727 396813
rect 100036 396808 100727 396810
rect 100036 396752 100666 396808
rect 100722 396752 100727 396808
rect 100036 396750 100727 396752
rect 100036 396748 100042 396750
rect 100661 396747 100727 396750
rect 101070 396748 101076 396812
rect 101140 396810 101146 396812
rect 102041 396810 102107 396813
rect 101140 396808 102107 396810
rect 101140 396752 102046 396808
rect 102102 396752 102107 396808
rect 101140 396750 102107 396752
rect 101140 396748 101146 396750
rect 102041 396747 102107 396750
rect 103513 396810 103579 396813
rect 105997 396812 106063 396813
rect 107469 396812 107535 396813
rect 103830 396810 103836 396812
rect 103513 396808 103836 396810
rect 103513 396752 103518 396808
rect 103574 396752 103836 396808
rect 103513 396750 103836 396752
rect 103513 396747 103579 396750
rect 103830 396748 103836 396750
rect 103900 396748 103906 396812
rect 105997 396808 106044 396812
rect 106108 396810 106114 396812
rect 105997 396752 106002 396808
rect 105997 396748 106044 396752
rect 106108 396750 106154 396810
rect 107469 396808 107516 396812
rect 107580 396810 107586 396812
rect 107469 396752 107474 396808
rect 106108 396748 106114 396750
rect 107469 396748 107516 396752
rect 107580 396750 107626 396810
rect 107580 396748 107586 396750
rect 111190 396748 111196 396812
rect 111260 396810 111266 396812
rect 111609 396810 111675 396813
rect 111260 396808 111675 396810
rect 111260 396752 111614 396808
rect 111670 396752 111675 396808
rect 111260 396750 111675 396752
rect 111260 396748 111266 396750
rect 105997 396747 106063 396748
rect 107469 396747 107535 396748
rect 111609 396747 111675 396750
rect 115749 396812 115815 396813
rect 115749 396808 115796 396812
rect 115860 396810 115866 396812
rect 115749 396752 115754 396808
rect 115749 396748 115796 396752
rect 115860 396750 115906 396810
rect 115860 396748 115866 396750
rect 117078 396748 117084 396812
rect 117148 396810 117154 396812
rect 117221 396810 117287 396813
rect 117148 396808 117287 396810
rect 117148 396752 117226 396808
rect 117282 396752 117287 396808
rect 117148 396750 117287 396752
rect 117148 396748 117154 396750
rect 115749 396747 115815 396748
rect 117221 396747 117287 396750
rect 119102 396748 119108 396812
rect 119172 396810 119178 396812
rect 119981 396810 120047 396813
rect 119172 396808 120047 396810
rect 119172 396752 119986 396808
rect 120042 396752 120047 396808
rect 119172 396750 120047 396752
rect 119172 396748 119178 396750
rect 119981 396747 120047 396750
rect 120758 396748 120764 396812
rect 120828 396810 120834 396812
rect 121269 396810 121335 396813
rect 120828 396808 121335 396810
rect 120828 396752 121274 396808
rect 121330 396752 121335 396808
rect 120828 396750 121335 396752
rect 120828 396748 120834 396750
rect 121269 396747 121335 396750
rect 123518 396748 123524 396812
rect 123588 396810 123594 396812
rect 124121 396810 124187 396813
rect 123588 396808 124187 396810
rect 123588 396752 124126 396808
rect 124182 396752 124187 396808
rect 123588 396750 124187 396752
rect 123588 396748 123594 396750
rect 124121 396747 124187 396750
rect 125910 396748 125916 396812
rect 125980 396810 125986 396812
rect 126881 396810 126947 396813
rect 125980 396808 126947 396810
rect 125980 396752 126886 396808
rect 126942 396752 126947 396808
rect 125980 396750 126947 396752
rect 125980 396748 125986 396750
rect 126881 396747 126947 396750
rect 128670 396748 128676 396812
rect 128740 396810 128746 396812
rect 129641 396810 129707 396813
rect 128740 396808 129707 396810
rect 128740 396752 129646 396808
rect 129702 396752 129707 396808
rect 128740 396750 129707 396752
rect 128740 396748 128746 396750
rect 129641 396747 129707 396750
rect 131021 396812 131087 396813
rect 131021 396808 131068 396812
rect 131132 396810 131138 396812
rect 131021 396752 131026 396808
rect 131021 396748 131068 396752
rect 131132 396750 131178 396810
rect 131132 396748 131138 396750
rect 133454 396748 133460 396812
rect 133524 396810 133530 396812
rect 133781 396810 133847 396813
rect 133524 396808 133847 396810
rect 133524 396752 133786 396808
rect 133842 396752 133847 396808
rect 133524 396750 133847 396752
rect 133524 396748 133530 396750
rect 131021 396747 131087 396748
rect 133781 396747 133847 396750
rect 138422 396748 138428 396812
rect 138492 396810 138498 396812
rect 139301 396810 139367 396813
rect 138492 396808 139367 396810
rect 138492 396752 139306 396808
rect 139362 396752 139367 396808
rect 138492 396750 139367 396752
rect 138492 396748 138498 396750
rect 139301 396747 139367 396750
rect 140998 396748 141004 396812
rect 141068 396810 141074 396812
rect 142061 396810 142127 396813
rect 141068 396808 142127 396810
rect 141068 396752 142066 396808
rect 142122 396752 142127 396808
rect 141068 396750 142127 396752
rect 141068 396748 141074 396750
rect 142061 396747 142127 396750
rect 143574 396748 143580 396812
rect 143644 396810 143650 396812
rect 144821 396810 144887 396813
rect 143644 396808 144887 396810
rect 143644 396752 144826 396808
rect 144882 396752 144887 396808
rect 143644 396750 144887 396752
rect 143644 396748 143650 396750
rect 144821 396747 144887 396750
rect 145005 396810 145071 396813
rect 145598 396810 145604 396812
rect 145005 396808 145604 396810
rect 145005 396752 145010 396808
rect 145066 396752 145604 396808
rect 145005 396750 145604 396752
rect 145005 396747 145071 396750
rect 145598 396748 145604 396750
rect 145668 396748 145674 396812
rect 148542 396748 148548 396812
rect 148612 396810 148618 396812
rect 148961 396810 149027 396813
rect 148612 396808 149027 396810
rect 148612 396752 148966 396808
rect 149022 396752 149027 396808
rect 148612 396750 149027 396752
rect 148612 396748 148618 396750
rect 148961 396747 149027 396750
rect 150934 396748 150940 396812
rect 151004 396810 151010 396812
rect 151721 396810 151787 396813
rect 155953 396812 156019 396813
rect 155902 396810 155908 396812
rect 151004 396808 151787 396810
rect 151004 396752 151726 396808
rect 151782 396752 151787 396808
rect 151004 396750 151787 396752
rect 155862 396750 155908 396810
rect 155972 396808 156019 396812
rect 156014 396752 156019 396808
rect 151004 396748 151010 396750
rect 151721 396747 151787 396750
rect 155902 396748 155908 396750
rect 155972 396748 156019 396752
rect 158478 396748 158484 396812
rect 158548 396810 158554 396812
rect 158621 396810 158687 396813
rect 158548 396808 158687 396810
rect 158548 396752 158626 396808
rect 158682 396752 158687 396808
rect 158548 396750 158687 396752
rect 158548 396748 158554 396750
rect 155953 396747 156019 396748
rect 158621 396747 158687 396750
rect 160870 396748 160876 396812
rect 160940 396810 160946 396812
rect 161381 396810 161447 396813
rect 160940 396808 161447 396810
rect 160940 396752 161386 396808
rect 161442 396752 161447 396808
rect 160940 396750 161447 396752
rect 160940 396748 160946 396750
rect 161381 396747 161447 396750
rect 166022 396748 166028 396812
rect 166092 396810 166098 396812
rect 166901 396810 166967 396813
rect 166092 396808 166967 396810
rect 166092 396752 166906 396808
rect 166962 396752 166967 396808
rect 166092 396750 166967 396752
rect 166092 396748 166098 396750
rect 166901 396747 166967 396750
rect 182173 396810 182239 396813
rect 183134 396810 183140 396812
rect 182173 396808 183140 396810
rect 182173 396752 182178 396808
rect 182234 396752 183140 396808
rect 182173 396750 183140 396752
rect 182173 396747 182239 396750
rect 183134 396748 183140 396750
rect 183204 396748 183210 396812
rect 237373 396810 237439 396813
rect 238150 396810 238156 396812
rect 237373 396808 238156 396810
rect 237373 396752 237378 396808
rect 237434 396752 238156 396808
rect 237373 396750 238156 396752
rect 237373 396747 237439 396750
rect 238150 396748 238156 396750
rect 238220 396748 238226 396812
rect 240133 396810 240199 396813
rect 240542 396810 240548 396812
rect 240133 396808 240548 396810
rect 240133 396752 240138 396808
rect 240194 396752 240548 396808
rect 240133 396750 240548 396752
rect 240133 396747 240199 396750
rect 240542 396748 240548 396750
rect 240612 396748 240618 396812
rect 241513 396810 241579 396813
rect 242893 396812 242959 396813
rect 241646 396810 241652 396812
rect 241513 396808 241652 396810
rect 241513 396752 241518 396808
rect 241574 396752 241652 396808
rect 241513 396750 241652 396752
rect 241513 396747 241579 396750
rect 241646 396748 241652 396750
rect 241716 396748 241722 396812
rect 242893 396808 242940 396812
rect 243004 396810 243010 396812
rect 242893 396752 242898 396808
rect 242893 396748 242940 396752
rect 243004 396750 243050 396810
rect 243004 396748 243010 396750
rect 244222 396748 244228 396812
rect 244292 396810 244298 396812
rect 244365 396810 244431 396813
rect 244292 396808 244431 396810
rect 244292 396752 244370 396808
rect 244426 396752 244431 396808
rect 244292 396750 244431 396752
rect 244292 396748 244298 396750
rect 242893 396747 242959 396748
rect 244365 396747 244431 396750
rect 244549 396810 244615 396813
rect 245326 396810 245332 396812
rect 244549 396808 245332 396810
rect 244549 396752 244554 396808
rect 244610 396752 245332 396808
rect 244549 396750 245332 396752
rect 244549 396747 244615 396750
rect 245326 396748 245332 396750
rect 245396 396748 245402 396812
rect 245653 396810 245719 396813
rect 246430 396810 246436 396812
rect 245653 396808 246436 396810
rect 245653 396752 245658 396808
rect 245714 396752 246436 396808
rect 245653 396750 246436 396752
rect 245653 396747 245719 396750
rect 246430 396748 246436 396750
rect 246500 396748 246506 396812
rect 251357 396810 251423 396813
rect 252318 396810 252324 396812
rect 251357 396808 252324 396810
rect 251357 396752 251362 396808
rect 251418 396752 252324 396808
rect 251357 396750 252324 396752
rect 251357 396747 251423 396750
rect 252318 396748 252324 396750
rect 252388 396748 252394 396812
rect 252553 396810 252619 396813
rect 253606 396810 253612 396812
rect 252553 396808 253612 396810
rect 252553 396752 252558 396808
rect 252614 396752 253612 396808
rect 252553 396750 253612 396752
rect 252553 396747 252619 396750
rect 253606 396748 253612 396750
rect 253676 396748 253682 396812
rect 254117 396810 254183 396813
rect 254526 396810 254532 396812
rect 254117 396808 254532 396810
rect 254117 396752 254122 396808
rect 254178 396752 254532 396808
rect 254117 396750 254532 396752
rect 254117 396747 254183 396750
rect 254526 396748 254532 396750
rect 254596 396748 254602 396812
rect 255405 396810 255471 396813
rect 256141 396812 256207 396813
rect 256877 396812 256943 396813
rect 255814 396810 255820 396812
rect 255405 396808 255820 396810
rect 255405 396752 255410 396808
rect 255466 396752 255820 396808
rect 255405 396750 255820 396752
rect 255405 396747 255471 396750
rect 255814 396748 255820 396750
rect 255884 396748 255890 396812
rect 256141 396808 256188 396812
rect 256252 396810 256258 396812
rect 256141 396752 256146 396808
rect 256141 396748 256188 396752
rect 256252 396750 256298 396810
rect 256877 396808 256924 396812
rect 256988 396810 256994 396812
rect 258165 396810 258231 396813
rect 258390 396810 258396 396812
rect 256877 396752 256882 396808
rect 256252 396748 256258 396750
rect 256877 396748 256924 396752
rect 256988 396750 257034 396810
rect 258165 396808 258396 396810
rect 258165 396752 258170 396808
rect 258226 396752 258396 396808
rect 258165 396750 258396 396752
rect 256988 396748 256994 396750
rect 256141 396747 256207 396748
rect 256877 396747 256943 396748
rect 258165 396747 258231 396750
rect 258390 396748 258396 396750
rect 258460 396748 258466 396812
rect 259545 396810 259611 396813
rect 260598 396810 260604 396812
rect 259545 396808 260604 396810
rect 259545 396752 259550 396808
rect 259606 396752 260604 396808
rect 259545 396750 260604 396752
rect 259545 396747 259611 396750
rect 260598 396748 260604 396750
rect 260668 396748 260674 396812
rect 263542 396748 263548 396812
rect 263612 396810 263618 396812
rect 263685 396810 263751 396813
rect 263612 396808 263751 396810
rect 263612 396752 263690 396808
rect 263746 396752 263751 396808
rect 263612 396750 263751 396752
rect 263612 396748 263618 396750
rect 263685 396747 263751 396750
rect 265157 396810 265223 396813
rect 266353 396812 266419 396813
rect 265934 396810 265940 396812
rect 265157 396808 265940 396810
rect 265157 396752 265162 396808
rect 265218 396752 265940 396808
rect 265157 396750 265940 396752
rect 265157 396747 265223 396750
rect 265934 396748 265940 396750
rect 266004 396748 266010 396812
rect 266302 396810 266308 396812
rect 266262 396750 266308 396810
rect 266372 396808 266419 396812
rect 266414 396752 266419 396808
rect 266302 396748 266308 396750
rect 266372 396748 266419 396752
rect 266353 396747 266419 396748
rect 269389 396810 269455 396813
rect 269798 396810 269804 396812
rect 269389 396808 269804 396810
rect 269389 396752 269394 396808
rect 269450 396752 269804 396808
rect 269389 396750 269804 396752
rect 269389 396747 269455 396750
rect 269798 396748 269804 396750
rect 269868 396748 269874 396812
rect 270493 396810 270559 396813
rect 273345 396812 273411 396813
rect 270902 396810 270908 396812
rect 270493 396808 270908 396810
rect 270493 396752 270498 396808
rect 270554 396752 270908 396808
rect 270493 396750 270908 396752
rect 270493 396747 270559 396750
rect 270902 396748 270908 396750
rect 270972 396748 270978 396812
rect 273294 396810 273300 396812
rect 273254 396750 273300 396810
rect 273364 396808 273411 396812
rect 273406 396752 273411 396808
rect 273294 396748 273300 396750
rect 273364 396748 273411 396752
rect 273345 396747 273411 396748
rect 273621 396810 273687 396813
rect 274398 396810 274404 396812
rect 273621 396808 274404 396810
rect 273621 396752 273626 396808
rect 273682 396752 274404 396808
rect 273621 396750 274404 396752
rect 273621 396747 273687 396750
rect 274398 396748 274404 396750
rect 274468 396748 274474 396812
rect 276105 396810 276171 396813
rect 276238 396810 276244 396812
rect 276105 396808 276244 396810
rect 276105 396752 276110 396808
rect 276166 396752 276244 396808
rect 276105 396750 276244 396752
rect 276105 396747 276171 396750
rect 276238 396748 276244 396750
rect 276308 396748 276314 396812
rect 277485 396810 277551 396813
rect 278446 396810 278452 396812
rect 277485 396808 278452 396810
rect 277485 396752 277490 396808
rect 277546 396752 278452 396808
rect 277485 396750 278452 396752
rect 277485 396747 277551 396750
rect 278446 396748 278452 396750
rect 278516 396748 278522 396812
rect 280153 396810 280219 396813
rect 283741 396812 283807 396813
rect 285949 396812 286015 396813
rect 280838 396810 280844 396812
rect 280153 396808 280844 396810
rect 280153 396752 280158 396808
rect 280214 396752 280844 396808
rect 280153 396750 280844 396752
rect 280153 396747 280219 396750
rect 280838 396748 280844 396750
rect 280908 396748 280914 396812
rect 283741 396808 283788 396812
rect 283852 396810 283858 396812
rect 283741 396752 283746 396808
rect 283741 396748 283788 396752
rect 283852 396750 283898 396810
rect 285949 396808 285996 396812
rect 286060 396810 286066 396812
rect 287053 396810 287119 396813
rect 288198 396810 288204 396812
rect 285949 396752 285954 396808
rect 283852 396748 283858 396750
rect 285949 396748 285996 396752
rect 286060 396750 286106 396810
rect 287053 396808 288204 396810
rect 287053 396752 287058 396808
rect 287114 396752 288204 396808
rect 287053 396750 288204 396752
rect 286060 396748 286066 396750
rect 283741 396747 283807 396748
rect 285949 396747 286015 396748
rect 287053 396747 287119 396750
rect 288198 396748 288204 396750
rect 288268 396748 288274 396812
rect 292665 396810 292731 396813
rect 293350 396810 293356 396812
rect 292665 396808 293356 396810
rect 292665 396752 292670 396808
rect 292726 396752 293356 396808
rect 292665 396750 293356 396752
rect 292665 396747 292731 396750
rect 293350 396748 293356 396750
rect 293420 396748 293426 396812
rect 295333 396810 295399 396813
rect 295926 396810 295932 396812
rect 295333 396808 295932 396810
rect 295333 396752 295338 396808
rect 295394 396752 295932 396808
rect 295333 396750 295932 396752
rect 295333 396747 295399 396750
rect 295926 396748 295932 396750
rect 295996 396748 296002 396812
rect 302233 396810 302299 396813
rect 303470 396810 303476 396812
rect 302233 396808 303476 396810
rect 302233 396752 302238 396808
rect 302294 396752 303476 396808
rect 302233 396750 303476 396752
rect 302233 396747 302299 396750
rect 303470 396748 303476 396750
rect 303540 396748 303546 396812
rect 304993 396810 305059 396813
rect 305862 396810 305868 396812
rect 304993 396808 305868 396810
rect 304993 396752 304998 396808
rect 305054 396752 305868 396808
rect 304993 396750 305868 396752
rect 304993 396747 305059 396750
rect 305862 396748 305868 396750
rect 305932 396748 305938 396812
rect 310513 396810 310579 396813
rect 311014 396810 311020 396812
rect 310513 396808 311020 396810
rect 310513 396752 310518 396808
rect 310574 396752 311020 396808
rect 310513 396750 311020 396752
rect 310513 396747 310579 396750
rect 311014 396748 311020 396750
rect 311084 396748 311090 396812
rect 313273 396810 313339 396813
rect 313406 396810 313412 396812
rect 313273 396808 313412 396810
rect 313273 396752 313278 396808
rect 313334 396752 313412 396808
rect 313273 396750 313412 396752
rect 313273 396747 313339 396750
rect 313406 396748 313412 396750
rect 313476 396748 313482 396812
rect 317413 396810 317479 396813
rect 318374 396810 318380 396812
rect 317413 396808 318380 396810
rect 317413 396752 317418 396808
rect 317474 396752 318380 396808
rect 317413 396750 318380 396752
rect 317413 396747 317479 396750
rect 318374 396748 318380 396750
rect 318444 396748 318450 396812
rect 320173 396810 320239 396813
rect 320950 396810 320956 396812
rect 320173 396808 320956 396810
rect 320173 396752 320178 396808
rect 320234 396752 320956 396808
rect 320173 396750 320956 396752
rect 320173 396747 320239 396750
rect 320950 396748 320956 396750
rect 321020 396748 321026 396812
rect 322933 396810 322999 396813
rect 323342 396810 323348 396812
rect 322933 396808 323348 396810
rect 322933 396752 322938 396808
rect 322994 396752 323348 396808
rect 322933 396750 323348 396752
rect 322933 396747 322999 396750
rect 323342 396748 323348 396750
rect 323412 396748 323418 396812
rect 342345 396810 342411 396813
rect 343398 396810 343404 396812
rect 342345 396808 343404 396810
rect 342345 396752 342350 396808
rect 342406 396752 343404 396808
rect 342345 396750 343404 396752
rect 342345 396747 342411 396750
rect 343398 396748 343404 396750
rect 343468 396748 343474 396812
rect 100753 396674 100819 396677
rect 101806 396674 101812 396676
rect 100753 396672 101812 396674
rect 100753 396616 100758 396672
rect 100814 396616 101812 396672
rect 100753 396614 101812 396616
rect 100753 396611 100819 396614
rect 101806 396612 101812 396614
rect 101876 396612 101882 396676
rect 107653 396674 107719 396677
rect 108246 396674 108252 396676
rect 107653 396672 108252 396674
rect 107653 396616 107658 396672
rect 107714 396616 108252 396672
rect 107653 396614 108252 396616
rect 107653 396611 107719 396614
rect 108246 396612 108252 396614
rect 108316 396612 108322 396676
rect 111006 396612 111012 396676
rect 111076 396674 111082 396676
rect 111517 396674 111583 396677
rect 111076 396672 111583 396674
rect 111076 396616 111522 396672
rect 111578 396616 111583 396672
rect 111076 396614 111583 396616
rect 111076 396612 111082 396614
rect 111517 396611 111583 396614
rect 115933 396676 115999 396677
rect 115933 396672 115980 396676
rect 116044 396674 116050 396676
rect 266445 396674 266511 396677
rect 267590 396674 267596 396676
rect 115933 396616 115938 396672
rect 115933 396612 115980 396616
rect 116044 396614 116090 396674
rect 266445 396672 267596 396674
rect 266445 396616 266450 396672
rect 266506 396616 267596 396672
rect 266445 396614 267596 396616
rect 116044 396612 116050 396614
rect 115933 396611 115999 396612
rect 266445 396611 266511 396614
rect 267590 396612 267596 396614
rect 267660 396612 267666 396676
rect 270585 396674 270651 396677
rect 273437 396676 273503 396677
rect 271270 396674 271276 396676
rect 270585 396672 271276 396674
rect 270585 396616 270590 396672
rect 270646 396616 271276 396672
rect 270585 396614 271276 396616
rect 270585 396611 270651 396614
rect 271270 396612 271276 396614
rect 271340 396612 271346 396676
rect 273437 396672 273484 396676
rect 273548 396674 273554 396676
rect 276013 396674 276079 396677
rect 276974 396674 276980 396676
rect 273437 396616 273442 396672
rect 273437 396612 273484 396616
rect 273548 396614 273594 396674
rect 276013 396672 276980 396674
rect 276013 396616 276018 396672
rect 276074 396616 276980 396672
rect 276013 396614 276980 396616
rect 273548 396612 273554 396614
rect 273437 396611 273503 396612
rect 276013 396611 276079 396614
rect 276974 396612 276980 396614
rect 277044 396612 277050 396676
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 579613 365122 579679 365125
rect 583520 365122 584960 365212
rect 579613 365120 584960 365122
rect 579613 365064 579618 365120
rect 579674 365064 584960 365120
rect 579613 365062 584960 365064
rect 579613 365059 579679 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect 201033 322146 201099 322149
rect 226374 322146 226380 322148
rect 201033 322144 226380 322146
rect 201033 322088 201038 322144
rect 201094 322088 226380 322144
rect 201033 322086 226380 322088
rect 201033 322083 201099 322086
rect 226374 322084 226380 322086
rect 226444 322084 226450 322148
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 209313 260130 209379 260133
rect 226742 260130 226748 260132
rect 209313 260128 226748 260130
rect 209313 260072 209318 260128
rect 209374 260072 226748 260128
rect 209313 260070 226748 260072
rect 209313 260067 209379 260070
rect 226742 260068 226748 260070
rect 226812 260068 226818 260132
rect 583520 258906 584960 258996
rect 583342 258846 584960 258906
rect 583342 258770 583402 258846
rect 583520 258770 584960 258846
rect 583342 258756 584960 258770
rect 583342 258710 583586 258756
rect 251909 257954 251975 257957
rect 583526 257954 583586 258710
rect 251909 257952 583586 257954
rect 251909 257896 251914 257952
rect 251970 257896 583586 257952
rect 251909 257894 583586 257896
rect 251909 257891 251975 257894
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 106641 254010 106707 254013
rect 106641 254008 107762 254010
rect 106641 253952 106646 254008
rect 106702 253952 107762 254008
rect 106641 253950 107762 253952
rect 106641 253947 106707 253950
rect 107702 253874 107762 253950
rect 110413 253874 110479 253877
rect 107702 253872 110479 253874
rect 107702 253816 110418 253872
rect 110474 253816 110479 253872
rect 107702 253814 110479 253816
rect 110413 253811 110479 253814
rect 110413 251834 110479 251837
rect 118693 251834 118759 251837
rect 110413 251832 118759 251834
rect 110413 251776 110418 251832
rect 110474 251776 118698 251832
rect 118754 251776 118759 251832
rect 110413 251774 118759 251776
rect 110413 251771 110479 251774
rect 118693 251771 118759 251774
rect 222101 251154 222167 251157
rect 222837 251154 222903 251157
rect 222101 251152 222903 251154
rect 222101 251096 222106 251152
rect 222162 251096 222842 251152
rect 222898 251096 222903 251152
rect 222101 251094 222903 251096
rect 222101 251091 222167 251094
rect 222837 251091 222903 251094
rect 58341 250474 58407 250477
rect 182173 250474 182239 250477
rect 58341 250472 182239 250474
rect 58341 250416 58346 250472
rect 58402 250416 182178 250472
rect 182234 250416 182239 250472
rect 58341 250414 182239 250416
rect 58341 250411 58407 250414
rect 182173 250411 182239 250414
rect 213453 250474 213519 250477
rect 227161 250474 227227 250477
rect 213453 250472 227227 250474
rect 213453 250416 213458 250472
rect 213514 250416 227166 250472
rect 227222 250416 227227 250472
rect 213453 250414 227227 250416
rect 213453 250411 213519 250414
rect 227161 250411 227227 250414
rect 129641 249114 129707 249117
rect 225321 249114 225387 249117
rect 129641 249112 225387 249114
rect 129641 249056 129646 249112
rect 129702 249056 225326 249112
rect 225382 249056 225387 249112
rect 129641 249054 225387 249056
rect 129641 249051 129707 249054
rect 225321 249051 225387 249054
rect 121269 247618 121335 247621
rect 225965 247618 226031 247621
rect 121269 247616 226031 247618
rect 121269 247560 121274 247616
rect 121330 247560 225970 247616
rect 226026 247560 226031 247616
rect 121269 247558 226031 247560
rect 121269 247555 121335 247558
rect 225965 247555 226031 247558
rect 101857 246394 101923 246397
rect 102041 246394 102107 246397
rect 101857 246392 102107 246394
rect 101857 246336 101862 246392
rect 101918 246336 102046 246392
rect 102102 246336 102107 246392
rect 101857 246334 102107 246336
rect 101857 246331 101923 246334
rect 102041 246331 102107 246334
rect 77201 245714 77267 245717
rect 260741 245714 260807 245717
rect 77201 245712 260807 245714
rect 77201 245656 77206 245712
rect 77262 245656 260746 245712
rect 260802 245656 260807 245712
rect 77201 245654 260807 245656
rect 77201 245651 77267 245654
rect 260741 245651 260807 245654
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 57237 243674 57303 243677
rect 198733 243674 198799 243677
rect 57237 243672 198799 243674
rect 57237 243616 57242 243672
rect 57298 243616 198738 243672
rect 198794 243616 198799 243672
rect 57237 243614 198799 243616
rect 57237 243611 57303 243614
rect 198733 243611 198799 243614
rect 57145 243538 57211 243541
rect 357525 243538 357591 243541
rect 57145 243536 357591 243538
rect 57145 243480 57150 243536
rect 57206 243480 357530 243536
rect 357586 243480 357591 243536
rect 57145 243478 357591 243480
rect 57145 243475 57211 243478
rect 357525 243475 357591 243478
rect 217225 242314 217291 242317
rect 232405 242314 232471 242317
rect 217225 242312 232471 242314
rect 217225 242256 217230 242312
rect 217286 242256 232410 242312
rect 232466 242256 232471 242312
rect 217225 242254 232471 242256
rect 217225 242251 217291 242254
rect 232405 242251 232471 242254
rect 54477 242178 54543 242181
rect 242893 242178 242959 242181
rect 54477 242176 242959 242178
rect 54477 242120 54482 242176
rect 54538 242120 242898 242176
rect 242954 242120 242959 242176
rect 54477 242118 242959 242120
rect 54477 242115 54543 242118
rect 242893 242115 242959 242118
rect -960 241090 480 241180
rect 4061 241090 4127 241093
rect -960 241088 4127 241090
rect -960 241032 4066 241088
rect 4122 241032 4127 241088
rect -960 241030 4127 241032
rect -960 240940 480 241030
rect 4061 241027 4127 241030
rect 105997 240954 106063 240957
rect 228081 240954 228147 240957
rect 105997 240952 228147 240954
rect 105997 240896 106002 240952
rect 106058 240896 228086 240952
rect 228142 240896 228147 240952
rect 105997 240894 228147 240896
rect 105997 240891 106063 240894
rect 228081 240891 228147 240894
rect 58249 240818 58315 240821
rect 270493 240818 270559 240821
rect 58249 240816 270559 240818
rect 58249 240760 58254 240816
rect 58310 240760 270498 240816
rect 270554 240760 270559 240816
rect 58249 240758 270559 240760
rect 58249 240755 58315 240758
rect 270493 240755 270559 240758
rect 56225 239594 56291 239597
rect 92473 239594 92539 239597
rect 56225 239592 92539 239594
rect 56225 239536 56230 239592
rect 56286 239536 92478 239592
rect 92534 239536 92539 239592
rect 56225 239534 92539 239536
rect 56225 239531 56291 239534
rect 92473 239531 92539 239534
rect 111609 239594 111675 239597
rect 229829 239594 229895 239597
rect 111609 239592 229895 239594
rect 111609 239536 111614 239592
rect 111670 239536 229834 239592
rect 229890 239536 229895 239592
rect 111609 239534 229895 239536
rect 111609 239531 111675 239534
rect 229829 239531 229895 239534
rect 57329 239458 57395 239461
rect 197721 239458 197787 239461
rect 57329 239456 197787 239458
rect 57329 239400 57334 239456
rect 57390 239400 197726 239456
rect 197782 239400 197787 239456
rect 57329 239398 197787 239400
rect 57329 239395 57395 239398
rect 197721 239395 197787 239398
rect 209129 239458 209195 239461
rect 227345 239458 227411 239461
rect 209129 239456 227411 239458
rect 209129 239400 209134 239456
rect 209190 239400 227350 239456
rect 227406 239400 227411 239456
rect 209129 239398 227411 239400
rect 209129 239395 209195 239398
rect 227345 239395 227411 239398
rect 217777 238234 217843 238237
rect 231209 238234 231275 238237
rect 217777 238232 231275 238234
rect 217777 238176 217782 238232
rect 217838 238176 231214 238232
rect 231270 238176 231275 238232
rect 217777 238174 231275 238176
rect 217777 238171 217843 238174
rect 231209 238171 231275 238174
rect 58065 238098 58131 238101
rect 100753 238098 100819 238101
rect 58065 238096 100819 238098
rect 58065 238040 58070 238096
rect 58126 238040 100758 238096
rect 100814 238040 100819 238096
rect 58065 238038 100819 238040
rect 58065 238035 58131 238038
rect 100753 238035 100819 238038
rect 124121 238098 124187 238101
rect 225413 238098 225479 238101
rect 124121 238096 225479 238098
rect 124121 238040 124126 238096
rect 124182 238040 225418 238096
rect 225474 238040 225479 238096
rect 124121 238038 225479 238040
rect 124121 238035 124187 238038
rect 225413 238035 225479 238038
rect 79317 237962 79383 237965
rect 251909 237962 251975 237965
rect 79317 237960 251975 237962
rect 79317 237904 79322 237960
rect 79378 237904 251914 237960
rect 251970 237904 251975 237960
rect 79317 237902 251975 237904
rect 79317 237899 79383 237902
rect 251909 237899 251975 237902
rect 115749 236874 115815 236877
rect 229921 236874 229987 236877
rect 115749 236872 229987 236874
rect 115749 236816 115754 236872
rect 115810 236816 229926 236872
rect 229982 236816 229987 236872
rect 115749 236814 229987 236816
rect 115749 236811 115815 236814
rect 229921 236811 229987 236814
rect 3417 236738 3483 236741
rect 150801 236738 150867 236741
rect 3417 236736 150867 236738
rect 3417 236680 3422 236736
rect 3478 236680 150806 236736
rect 150862 236680 150867 236736
rect 3417 236678 150867 236680
rect 3417 236675 3483 236678
rect 150801 236675 150867 236678
rect 56409 236602 56475 236605
rect 320173 236602 320239 236605
rect 56409 236600 320239 236602
rect 56409 236544 56414 236600
rect 56470 236544 320178 236600
rect 320234 236544 320239 236600
rect 56409 236542 320239 236544
rect 56409 236539 56475 236542
rect 320173 236539 320239 236542
rect 55949 235378 56015 235381
rect 107653 235378 107719 235381
rect 55949 235376 107719 235378
rect 55949 235320 55954 235376
rect 56010 235320 107658 235376
rect 107714 235320 107719 235376
rect 55949 235318 107719 235320
rect 55949 235315 56015 235318
rect 107653 235315 107719 235318
rect 126881 235378 126947 235381
rect 226057 235378 226123 235381
rect 126881 235376 226123 235378
rect 126881 235320 126886 235376
rect 126942 235320 226062 235376
rect 226118 235320 226123 235376
rect 126881 235318 226123 235320
rect 126881 235315 126947 235318
rect 226057 235315 226123 235318
rect 58157 235242 58223 235245
rect 322933 235242 322999 235245
rect 58157 235240 322999 235242
rect 58157 235184 58162 235240
rect 58218 235184 322938 235240
rect 322994 235184 322999 235240
rect 58157 235182 322999 235184
rect 58157 235179 58223 235182
rect 322933 235179 322999 235182
rect 67357 234698 67423 234701
rect 253289 234698 253355 234701
rect 67357 234696 253355 234698
rect 67357 234640 67362 234696
rect 67418 234640 253294 234696
rect 253350 234640 253355 234696
rect 67357 234638 253355 234640
rect 67357 234635 67423 234638
rect 253289 234635 253355 234638
rect 224902 234500 224908 234564
rect 224972 234562 224978 234564
rect 226006 234562 226012 234564
rect 224972 234502 226012 234562
rect 224972 234500 224978 234502
rect 226006 234500 226012 234502
rect 226076 234500 226082 234564
rect 213269 234290 213335 234293
rect 227529 234290 227595 234293
rect 213269 234288 227595 234290
rect 213269 234232 213274 234288
rect 213330 234232 227534 234288
rect 227590 234232 227595 234288
rect 213269 234230 227595 234232
rect 213269 234227 213335 234230
rect 227529 234227 227595 234230
rect 199377 234154 199443 234157
rect 228173 234154 228239 234157
rect 199377 234152 228239 234154
rect 199377 234096 199382 234152
rect 199438 234096 228178 234152
rect 228234 234096 228239 234152
rect 199377 234094 228239 234096
rect 199377 234091 199443 234094
rect 228173 234091 228239 234094
rect 96521 234018 96587 234021
rect 226241 234018 226307 234021
rect 96521 234016 226307 234018
rect 96521 233960 96526 234016
rect 96582 233960 226246 234016
rect 226302 233960 226307 234016
rect 96521 233958 226307 233960
rect 96521 233955 96587 233958
rect 226241 233955 226307 233958
rect 4153 233882 4219 233885
rect 149697 233882 149763 233885
rect 4153 233880 149763 233882
rect 4153 233824 4158 233880
rect 4214 233824 149702 233880
rect 149758 233824 149763 233880
rect 4153 233822 149763 233824
rect 4153 233819 4219 233822
rect 149697 233819 149763 233822
rect 168373 233882 168439 233885
rect 169293 233882 169359 233885
rect 224217 233882 224283 233885
rect 168373 233880 169359 233882
rect 168373 233824 168378 233880
rect 168434 233824 169298 233880
rect 169354 233824 169359 233880
rect 168373 233822 169359 233824
rect 168373 233819 168439 233822
rect 169293 233819 169359 233822
rect 171090 233880 224283 233882
rect 171090 233824 224222 233880
rect 224278 233824 224283 233880
rect 171090 233822 224283 233824
rect 124213 233746 124279 233749
rect 124857 233746 124923 233749
rect 124213 233744 124923 233746
rect 124213 233688 124218 233744
rect 124274 233688 124862 233744
rect 124918 233688 124923 233744
rect 124213 233686 124923 233688
rect 124213 233683 124279 233686
rect 124857 233683 124923 233686
rect 126973 233746 127039 233749
rect 127617 233746 127683 233749
rect 126973 233744 127683 233746
rect 126973 233688 126978 233744
rect 127034 233688 127622 233744
rect 127678 233688 127683 233744
rect 126973 233686 127683 233688
rect 126973 233683 127039 233686
rect 127617 233683 127683 233686
rect 129733 233746 129799 233749
rect 130377 233746 130443 233749
rect 129733 233744 130443 233746
rect 129733 233688 129738 233744
rect 129794 233688 130382 233744
rect 130438 233688 130443 233744
rect 129733 233686 130443 233688
rect 129733 233683 129799 233686
rect 130377 233683 130443 233686
rect 132493 233746 132559 233749
rect 133137 233746 133203 233749
rect 132493 233744 133203 233746
rect 132493 233688 132498 233744
rect 132554 233688 133142 233744
rect 133198 233688 133203 233744
rect 132493 233686 133203 233688
rect 132493 233683 132559 233686
rect 133137 233683 133203 233686
rect 135253 233746 135319 233749
rect 135897 233746 135963 233749
rect 135253 233744 135963 233746
rect 135253 233688 135258 233744
rect 135314 233688 135902 233744
rect 135958 233688 135963 233744
rect 135253 233686 135963 233688
rect 135253 233683 135319 233686
rect 135897 233683 135963 233686
rect 138013 233746 138079 233749
rect 138657 233746 138723 233749
rect 138013 233744 138723 233746
rect 138013 233688 138018 233744
rect 138074 233688 138662 233744
rect 138718 233688 138723 233744
rect 138013 233686 138723 233688
rect 138013 233683 138079 233686
rect 138657 233683 138723 233686
rect 140773 233746 140839 233749
rect 141417 233746 141483 233749
rect 140773 233744 141483 233746
rect 140773 233688 140778 233744
rect 140834 233688 141422 233744
rect 141478 233688 141483 233744
rect 140773 233686 141483 233688
rect 140773 233683 140839 233686
rect 141417 233683 141483 233686
rect 166901 233746 166967 233749
rect 171090 233746 171150 233822
rect 224217 233819 224283 233822
rect 166901 233744 171150 233746
rect 166901 233688 166906 233744
rect 166962 233688 171150 233744
rect 166901 233686 171150 233688
rect 177297 233746 177363 233749
rect 177941 233746 178007 233749
rect 177297 233744 178007 233746
rect 177297 233688 177302 233744
rect 177358 233688 177946 233744
rect 178002 233688 178007 233744
rect 177297 233686 178007 233688
rect 166901 233683 166967 233686
rect 177297 233683 177363 233686
rect 177941 233683 178007 233686
rect 181161 233746 181227 233749
rect 182081 233746 182147 233749
rect 181161 233744 182147 233746
rect 181161 233688 181166 233744
rect 181222 233688 182086 233744
rect 182142 233688 182147 233744
rect 181161 233686 182147 233688
rect 181161 233683 181227 233686
rect 182081 233683 182147 233686
rect 183921 233746 183987 233749
rect 184841 233746 184907 233749
rect 183921 233744 184907 233746
rect 183921 233688 183926 233744
rect 183982 233688 184846 233744
rect 184902 233688 184907 233744
rect 183921 233686 184907 233688
rect 183921 233683 183987 233686
rect 184841 233683 184907 233686
rect 192201 233746 192267 233749
rect 193121 233746 193187 233749
rect 192201 233744 193187 233746
rect 192201 233688 192206 233744
rect 192262 233688 193126 233744
rect 193182 233688 193187 233744
rect 192201 233686 193187 233688
rect 192201 233683 192267 233686
rect 193121 233683 193187 233686
rect 200481 233746 200547 233749
rect 201401 233746 201467 233749
rect 200481 233744 201467 233746
rect 200481 233688 200486 233744
rect 200542 233688 201406 233744
rect 201462 233688 201467 233744
rect 200481 233686 201467 233688
rect 200481 233683 200547 233686
rect 201401 233683 201467 233686
rect 17217 233474 17283 233477
rect 155401 233474 155467 233477
rect 17217 233472 155467 233474
rect 17217 233416 17222 233472
rect 17278 233416 155406 233472
rect 155462 233416 155467 233472
rect 17217 233414 155467 233416
rect 17217 233411 17283 233414
rect 155401 233411 155467 233414
rect 21357 233338 21423 233341
rect 161013 233338 161079 233341
rect 21357 233336 161079 233338
rect 21357 233280 21362 233336
rect 21418 233280 161018 233336
rect 161074 233280 161079 233336
rect 21357 233278 161079 233280
rect 21357 233275 21423 233278
rect 161013 233275 161079 233278
rect 216305 232794 216371 232797
rect 226558 232794 226564 232796
rect 216305 232792 226564 232794
rect 216305 232736 216310 232792
rect 216366 232736 226564 232792
rect 216305 232734 226564 232736
rect 216305 232731 216371 232734
rect 226558 232732 226564 232734
rect 226628 232732 226634 232796
rect 199561 232658 199627 232661
rect 228265 232658 228331 232661
rect 199561 232656 228331 232658
rect 199561 232600 199566 232656
rect 199622 232600 228270 232656
rect 228326 232600 228331 232656
rect 199561 232598 228331 232600
rect 199561 232595 199627 232598
rect 228265 232595 228331 232598
rect 32397 232522 32463 232525
rect 158161 232522 158227 232525
rect 32397 232520 158227 232522
rect 32397 232464 32402 232520
rect 32458 232464 158166 232520
rect 158222 232464 158227 232520
rect 32397 232462 158227 232464
rect 32397 232459 32463 232462
rect 158161 232459 158227 232462
rect 158621 232522 158687 232525
rect 226149 232522 226215 232525
rect 158621 232520 226215 232522
rect 158621 232464 158626 232520
rect 158682 232464 226154 232520
rect 226210 232464 226215 232520
rect 158621 232462 226215 232464
rect 158621 232459 158687 232462
rect 226149 232459 226215 232462
rect 29637 232386 29703 232389
rect 160185 232386 160251 232389
rect 583520 232386 584960 232476
rect 29637 232384 160251 232386
rect 29637 232328 29642 232384
rect 29698 232328 160190 232384
rect 160246 232328 160251 232384
rect 29637 232326 160251 232328
rect 29637 232323 29703 232326
rect 160185 232323 160251 232326
rect 583342 232326 584960 232386
rect 3509 232250 3575 232253
rect 158713 232250 158779 232253
rect 3509 232248 158779 232250
rect 3509 232192 3514 232248
rect 3570 232192 158718 232248
rect 158774 232192 158779 232248
rect 3509 232190 158779 232192
rect 583342 232250 583402 232326
rect 583520 232250 584960 232326
rect 583342 232236 584960 232250
rect 583342 232190 583586 232236
rect 3509 232187 3575 232190
rect 158713 232187 158779 232190
rect 4797 232114 4863 232117
rect 162853 232114 162919 232117
rect 4797 232112 162919 232114
rect 4797 232056 4802 232112
rect 4858 232056 162858 232112
rect 162914 232056 162919 232112
rect 4797 232054 162919 232056
rect 4797 232051 4863 232054
rect 162853 232051 162919 232054
rect 75637 231978 75703 231981
rect 583526 231978 583586 232190
rect 75637 231976 583586 231978
rect 75637 231920 75642 231976
rect 75698 231920 583586 231976
rect 75637 231918 583586 231920
rect 75637 231915 75703 231918
rect 218329 231570 218395 231573
rect 226190 231570 226196 231572
rect 218329 231568 226196 231570
rect 218329 231512 218334 231568
rect 218390 231512 226196 231568
rect 218329 231510 226196 231512
rect 218329 231507 218395 231510
rect 226190 231508 226196 231510
rect 226260 231508 226266 231572
rect 218881 231434 218947 231437
rect 227621 231434 227687 231437
rect 218881 231432 227687 231434
rect 218881 231376 218886 231432
rect 218942 231376 227626 231432
rect 227682 231376 227687 231432
rect 218881 231374 227687 231376
rect 218881 231371 218947 231374
rect 227621 231371 227687 231374
rect 11697 231298 11763 231301
rect 152089 231298 152155 231301
rect 11697 231296 152155 231298
rect 11697 231240 11702 231296
rect 11758 231240 152094 231296
rect 152150 231240 152155 231296
rect 11697 231238 152155 231240
rect 11697 231235 11763 231238
rect 152089 231235 152155 231238
rect 218697 231298 218763 231301
rect 226977 231298 227043 231301
rect 218697 231296 227043 231298
rect 218697 231240 218702 231296
rect 218758 231240 226982 231296
rect 227038 231240 227043 231296
rect 218697 231238 227043 231240
rect 218697 231235 218763 231238
rect 226977 231235 227043 231238
rect 14457 231162 14523 231165
rect 154849 231162 154915 231165
rect 14457 231160 154915 231162
rect 14457 231104 14462 231160
rect 14518 231104 154854 231160
rect 154910 231104 154915 231160
rect 14457 231102 154915 231104
rect 14457 231099 14523 231102
rect 154849 231099 154915 231102
rect 217869 231162 217935 231165
rect 229737 231162 229803 231165
rect 217869 231160 229803 231162
rect 217869 231104 217874 231160
rect 217930 231104 229742 231160
rect 229798 231104 229803 231160
rect 217869 231102 229803 231104
rect 217869 231099 217935 231102
rect 229737 231099 229803 231102
rect 15837 231026 15903 231029
rect 157609 231026 157675 231029
rect 15837 231024 157675 231026
rect 15837 230968 15842 231024
rect 15898 230968 157614 231024
rect 157670 230968 157675 231024
rect 15837 230966 157675 230968
rect 15837 230963 15903 230966
rect 157609 230963 157675 230966
rect 218513 231026 218579 231029
rect 224718 231026 224724 231028
rect 218513 231024 224724 231026
rect 218513 230968 218518 231024
rect 218574 230968 224724 231024
rect 218513 230966 224724 230968
rect 218513 230963 218579 230966
rect 224718 230964 224724 230966
rect 224788 230964 224794 231028
rect 68737 230890 68803 230893
rect 236637 230890 236703 230893
rect 68737 230888 236703 230890
rect 68737 230832 68742 230888
rect 68798 230832 236642 230888
rect 236698 230832 236703 230888
rect 68737 230830 236703 230832
rect 68737 230827 68803 230830
rect 236637 230827 236703 230830
rect 65977 230754 66043 230757
rect 235349 230754 235415 230757
rect 65977 230752 235415 230754
rect 65977 230696 65982 230752
rect 66038 230696 235354 230752
rect 235410 230696 235415 230752
rect 65977 230694 235415 230696
rect 65977 230691 66043 230694
rect 235349 230691 235415 230694
rect 70393 230618 70459 230621
rect 580257 230618 580323 230621
rect 70393 230616 580323 230618
rect 70393 230560 70398 230616
rect 70454 230560 580262 230616
rect 580318 230560 580323 230616
rect 70393 230558 580323 230560
rect 70393 230555 70459 230558
rect 580257 230555 580323 230558
rect 90265 230482 90331 230485
rect 91001 230482 91067 230485
rect 90265 230480 91067 230482
rect 90265 230424 90270 230480
rect 90326 230424 91006 230480
rect 91062 230424 91067 230480
rect 90265 230422 91067 230424
rect 90265 230419 90331 230422
rect 91001 230419 91067 230422
rect 93209 230482 93275 230485
rect 93761 230482 93827 230485
rect 93209 230480 93827 230482
rect 93209 230424 93214 230480
rect 93270 230424 93766 230480
rect 93822 230424 93827 230480
rect 93209 230422 93827 230424
rect 93209 230419 93275 230422
rect 93761 230419 93827 230422
rect 98729 230482 98795 230485
rect 99281 230482 99347 230485
rect 98729 230480 99347 230482
rect 98729 230424 98734 230480
rect 98790 230424 99286 230480
rect 99342 230424 99347 230480
rect 98729 230422 99347 230424
rect 98729 230419 98795 230422
rect 99281 230419 99347 230422
rect 104249 230482 104315 230485
rect 104801 230482 104867 230485
rect 104249 230480 104867 230482
rect 104249 230424 104254 230480
rect 104310 230424 104806 230480
rect 104862 230424 104867 230480
rect 104249 230422 104867 230424
rect 104249 230419 104315 230422
rect 104801 230419 104867 230422
rect 188153 230482 188219 230485
rect 200757 230482 200823 230485
rect 188153 230480 200823 230482
rect 188153 230424 188158 230480
rect 188214 230424 200762 230480
rect 200818 230424 200823 230480
rect 188153 230422 200823 230424
rect 188153 230419 188219 230422
rect 200757 230419 200823 230422
rect 206001 230482 206067 230485
rect 206921 230482 206987 230485
rect 206001 230480 206987 230482
rect 206001 230424 206006 230480
rect 206062 230424 206926 230480
rect 206982 230424 206987 230480
rect 206001 230422 206987 230424
rect 206001 230419 206067 230422
rect 206921 230419 206987 230422
rect 208761 230482 208827 230485
rect 209681 230482 209747 230485
rect 208761 230480 209747 230482
rect 208761 230424 208766 230480
rect 208822 230424 209686 230480
rect 209742 230424 209747 230480
rect 208761 230422 209747 230424
rect 208761 230419 208827 230422
rect 209681 230419 209747 230422
rect 211153 230482 211219 230485
rect 211981 230482 212047 230485
rect 211153 230480 212047 230482
rect 211153 230424 211158 230480
rect 211214 230424 211986 230480
rect 212042 230424 212047 230480
rect 211153 230422 212047 230424
rect 211153 230419 211219 230422
rect 211981 230419 212047 230422
rect 214465 230482 214531 230485
rect 215201 230482 215267 230485
rect 214465 230480 215267 230482
rect 214465 230424 214470 230480
rect 214526 230424 215206 230480
rect 215262 230424 215267 230480
rect 214465 230422 215267 230424
rect 214465 230419 214531 230422
rect 215201 230419 215267 230422
rect 216397 230482 216463 230485
rect 217777 230482 217843 230485
rect 216397 230480 217843 230482
rect 216397 230424 216402 230480
rect 216458 230424 217782 230480
rect 217838 230424 217843 230480
rect 216397 230422 217843 230424
rect 216397 230419 216463 230422
rect 217777 230419 217843 230422
rect 219065 230482 219131 230485
rect 223297 230482 223363 230485
rect 219065 230480 223363 230482
rect 219065 230424 219070 230480
rect 219126 230424 223302 230480
rect 223358 230424 223363 230480
rect 219065 230422 223363 230424
rect 219065 230419 219131 230422
rect 223297 230419 223363 230422
rect 179781 230346 179847 230349
rect 190729 230346 190795 230349
rect 179781 230344 190795 230346
rect 179781 230288 179786 230344
rect 179842 230288 190734 230344
rect 190790 230288 190795 230344
rect 179781 230286 190795 230288
rect 179781 230283 179847 230286
rect 190729 230283 190795 230286
rect 190913 230346 190979 230349
rect 196801 230346 196867 230349
rect 190913 230344 196867 230346
rect 190913 230288 190918 230344
rect 190974 230288 196806 230344
rect 196862 230288 196867 230344
rect 190913 230286 196867 230288
rect 190913 230283 190979 230286
rect 196801 230283 196867 230286
rect 198089 230346 198155 230349
rect 199285 230346 199351 230349
rect 198089 230344 199351 230346
rect 198089 230288 198094 230344
rect 198150 230288 199290 230344
rect 199346 230288 199351 230344
rect 198089 230286 199351 230288
rect 198089 230283 198155 230286
rect 199285 230283 199351 230286
rect 216213 230346 216279 230349
rect 220537 230346 220603 230349
rect 216213 230344 220603 230346
rect 216213 230288 216218 230344
rect 216274 230288 220542 230344
rect 220598 230288 220603 230344
rect 216213 230286 220603 230288
rect 216213 230283 216279 230286
rect 220537 230283 220603 230286
rect 182633 230210 182699 230213
rect 202137 230210 202203 230213
rect 182633 230208 202203 230210
rect 182633 230152 182638 230208
rect 182694 230152 202142 230208
rect 202198 230152 202203 230208
rect 182633 230150 202203 230152
rect 182633 230147 182699 230150
rect 202137 230147 202203 230150
rect 58525 230074 58591 230077
rect 121545 230074 121611 230077
rect 58525 230072 121611 230074
rect 58525 230016 58530 230072
rect 58586 230016 121550 230072
rect 121606 230016 121611 230072
rect 58525 230014 121611 230016
rect 58525 230011 58591 230014
rect 121545 230011 121611 230014
rect 174261 230074 174327 230077
rect 190821 230074 190887 230077
rect 197353 230074 197419 230077
rect 174261 230072 190746 230074
rect 174261 230016 174266 230072
rect 174322 230016 190746 230072
rect 174261 230014 190746 230016
rect 174261 230011 174327 230014
rect 58433 229938 58499 229941
rect 123385 229938 123451 229941
rect 58433 229936 123451 229938
rect 58433 229880 58438 229936
rect 58494 229880 123390 229936
rect 123446 229880 123451 229936
rect 58433 229878 123451 229880
rect 58433 229875 58499 229878
rect 123385 229875 123451 229878
rect 171501 229938 171567 229941
rect 190453 229938 190519 229941
rect 171501 229936 190519 229938
rect 171501 229880 171506 229936
rect 171562 229880 190458 229936
rect 190514 229880 190519 229936
rect 171501 229878 190519 229880
rect 190686 229938 190746 230014
rect 190821 230072 197419 230074
rect 190821 230016 190826 230072
rect 190882 230016 197358 230072
rect 197414 230016 197419 230072
rect 190821 230014 197419 230016
rect 190821 230011 190887 230014
rect 197353 230011 197419 230014
rect 197445 229938 197511 229941
rect 190686 229936 197511 229938
rect 190686 229880 197450 229936
rect 197506 229880 197511 229936
rect 190686 229878 197511 229880
rect 171501 229875 171567 229878
rect 190453 229875 190519 229878
rect 197445 229875 197511 229878
rect 216029 229938 216095 229941
rect 226926 229938 226932 229940
rect 216029 229936 226932 229938
rect 216029 229880 216034 229936
rect 216090 229880 226932 229936
rect 216029 229878 226932 229880
rect 216029 229875 216095 229878
rect 226926 229876 226932 229878
rect 226996 229876 227002 229940
rect 63217 229802 63283 229805
rect 70393 229802 70459 229805
rect 63217 229800 70459 229802
rect 63217 229744 63222 229800
rect 63278 229744 70398 229800
rect 70454 229744 70459 229800
rect 63217 229742 70459 229744
rect 63217 229739 63283 229742
rect 70393 229739 70459 229742
rect 74533 229802 74599 229805
rect 153929 229802 153995 229805
rect 74533 229800 153995 229802
rect 74533 229744 74538 229800
rect 74594 229744 153934 229800
rect 153990 229744 153995 229800
rect 74533 229742 153995 229744
rect 74533 229739 74599 229742
rect 153929 229739 153995 229742
rect 158713 229802 158779 229805
rect 164969 229802 165035 229805
rect 158713 229800 165035 229802
rect 158713 229744 158718 229800
rect 158774 229744 164974 229800
rect 165030 229744 165035 229800
rect 158713 229742 165035 229744
rect 158713 229739 158779 229742
rect 164969 229739 165035 229742
rect 167821 229802 167887 229805
rect 190453 229802 190519 229805
rect 167821 229800 190519 229802
rect 167821 229744 167826 229800
rect 167882 229744 190458 229800
rect 190514 229744 190519 229800
rect 167821 229742 190519 229744
rect 167821 229739 167887 229742
rect 190453 229739 190519 229742
rect 190637 229802 190703 229805
rect 197537 229802 197603 229805
rect 190637 229800 197603 229802
rect 190637 229744 190642 229800
rect 190698 229744 197542 229800
rect 197598 229744 197603 229800
rect 190637 229742 197603 229744
rect 190637 229739 190703 229742
rect 197537 229739 197603 229742
rect 210509 229802 210575 229805
rect 227437 229802 227503 229805
rect 210509 229800 227503 229802
rect 210509 229744 210514 229800
rect 210570 229744 227442 229800
rect 227498 229744 227503 229800
rect 210509 229742 227503 229744
rect 210509 229739 210575 229742
rect 227437 229739 227503 229742
rect 70301 229666 70367 229669
rect 156689 229666 156755 229669
rect 70301 229664 156755 229666
rect 70301 229608 70306 229664
rect 70362 229608 156694 229664
rect 156750 229608 156755 229664
rect 70301 229606 156755 229608
rect 70301 229603 70367 229606
rect 156689 229603 156755 229606
rect 186313 229666 186379 229669
rect 196709 229666 196775 229669
rect 186313 229664 196775 229666
rect 186313 229608 186318 229664
rect 186374 229608 196714 229664
rect 196770 229608 196775 229664
rect 186313 229606 196775 229608
rect 186313 229603 186379 229606
rect 196709 229603 196775 229606
rect 71681 229530 71747 229533
rect 162209 229530 162275 229533
rect 71681 229528 162275 229530
rect 71681 229472 71686 229528
rect 71742 229472 162214 229528
rect 162270 229472 162275 229528
rect 71681 229470 162275 229472
rect 71681 229467 71747 229470
rect 162209 229467 162275 229470
rect 190453 229530 190519 229533
rect 197629 229530 197695 229533
rect 190453 229528 197695 229530
rect 190453 229472 190458 229528
rect 190514 229472 197634 229528
rect 197690 229472 197695 229528
rect 190453 229470 197695 229472
rect 190453 229467 190519 229470
rect 197629 229467 197695 229470
rect 64137 229394 64203 229397
rect 182173 229394 182239 229397
rect 64137 229392 182239 229394
rect 64137 229336 64142 229392
rect 64198 229336 182178 229392
rect 182234 229336 182239 229392
rect 64137 229334 182239 229336
rect 64137 229331 64203 229334
rect 182173 229331 182239 229334
rect 18597 229258 18663 229261
rect 155861 229258 155927 229261
rect 164049 229258 164115 229261
rect 18597 229256 155602 229258
rect 18597 229200 18602 229256
rect 18658 229200 155602 229256
rect 18597 229198 155602 229200
rect 18597 229195 18663 229198
rect 7557 229122 7623 229125
rect 153009 229122 153075 229125
rect 7557 229120 153075 229122
rect 7557 229064 7562 229120
rect 7618 229064 153014 229120
rect 153070 229064 153075 229120
rect 7557 229062 153075 229064
rect 155542 229122 155602 229198
rect 155861 229256 164115 229258
rect 155861 229200 155866 229256
rect 155922 229200 164054 229256
rect 164110 229200 164115 229256
rect 155861 229198 164115 229200
rect 155861 229195 155927 229198
rect 164049 229195 164115 229198
rect 159449 229122 159515 229125
rect 155542 229120 159515 229122
rect 155542 229064 159454 229120
rect 159510 229064 159515 229120
rect 155542 229062 159515 229064
rect 7557 229059 7623 229062
rect 153009 229059 153075 229062
rect 159449 229059 159515 229062
rect 84469 228986 84535 228989
rect 85481 228986 85547 228989
rect 84469 228984 85547 228986
rect 84469 228928 84474 228984
rect 84530 228928 85486 228984
rect 85542 228928 85547 228984
rect 84469 228926 85547 228928
rect 84469 228923 84535 228926
rect 85481 228923 85547 228926
rect 87229 228986 87295 228989
rect 88241 228986 88307 228989
rect 87229 228984 88307 228986
rect 87229 228928 87234 228984
rect 87290 228928 88246 228984
rect 88302 228928 88307 228984
rect 87229 228926 88307 228928
rect 87229 228923 87295 228926
rect 88241 228923 88307 228926
rect 95601 228986 95667 228989
rect 96429 228986 96495 228989
rect 95601 228984 96495 228986
rect 95601 228928 95606 228984
rect 95662 228928 96434 228984
rect 96490 228928 96495 228984
rect 95601 228926 96495 228928
rect 95601 228923 95667 228926
rect 96429 228923 96495 228926
rect 223665 228850 223731 228853
rect 224166 228850 224172 228852
rect 223665 228848 224172 228850
rect 223665 228792 223670 228848
rect 223726 228792 224172 228848
rect 223665 228790 224172 228792
rect 223665 228787 223731 228790
rect 224166 228788 224172 228790
rect 224236 228788 224242 228852
rect 217133 228714 217199 228717
rect 225689 228714 225755 228717
rect 217133 228712 225755 228714
rect 217133 228656 217138 228712
rect 217194 228656 225694 228712
rect 225750 228656 225755 228712
rect 217133 228654 225755 228656
rect 217133 228651 217199 228654
rect 225689 228651 225755 228654
rect 3601 228578 3667 228581
rect 71681 228578 71747 228581
rect 3601 228576 71747 228578
rect 3601 228520 3606 228576
rect 3662 228520 71686 228576
rect 71742 228520 71747 228576
rect 3601 228518 71747 228520
rect 3601 228515 3667 228518
rect 71681 228515 71747 228518
rect 199469 228578 199535 228581
rect 225781 228578 225847 228581
rect 199469 228576 225847 228578
rect 199469 228520 199474 228576
rect 199530 228520 225786 228576
rect 225842 228520 225847 228576
rect 199469 228518 225847 228520
rect 199469 228515 199535 228518
rect 225781 228515 225847 228518
rect 3785 228442 3851 228445
rect 74533 228442 74599 228445
rect 3785 228440 74599 228442
rect 3785 228384 3790 228440
rect 3846 228384 74538 228440
rect 74594 228384 74599 228440
rect 3785 228382 74599 228384
rect 3785 228379 3851 228382
rect 74533 228379 74599 228382
rect 76189 228442 76255 228445
rect 234429 228442 234495 228445
rect 76189 228440 234495 228442
rect 76189 228384 76194 228440
rect 76250 228384 234434 228440
rect 234490 228384 234495 228440
rect 76189 228382 234495 228384
rect 76189 228379 76255 228382
rect 234429 228379 234495 228382
rect 3417 228306 3483 228309
rect 155861 228306 155927 228309
rect 3417 228304 155927 228306
rect 3417 228248 3422 228304
rect 3478 228248 155866 228304
rect 155922 228248 155927 228304
rect 3417 228246 155927 228248
rect 3417 228243 3483 228246
rect 155861 228243 155927 228246
rect 182173 228306 182239 228309
rect 580349 228306 580415 228309
rect 182173 228304 580415 228306
rect 182173 228248 182178 228304
rect 182234 228248 580354 228304
rect 580410 228248 580415 228304
rect 182173 228246 580415 228248
rect 182173 228243 182239 228246
rect 580349 228243 580415 228246
rect 73337 228170 73403 228173
rect 236729 228170 236795 228173
rect 73337 228168 236795 228170
rect -960 227884 480 228124
rect 73337 228112 73342 228168
rect 73398 228112 236734 228168
rect 236790 228112 236795 228168
rect 73337 228110 236795 228112
rect 73337 228107 73403 228110
rect 236729 228107 236795 228110
rect 70577 228034 70643 228037
rect 239397 228034 239463 228037
rect 70577 228032 239463 228034
rect 70577 227976 70582 228032
rect 70638 227976 239402 228032
rect 239458 227976 239463 228032
rect 70577 227974 239463 227976
rect 70577 227971 70643 227974
rect 239397 227971 239463 227974
rect 65057 227898 65123 227901
rect 240869 227898 240935 227901
rect 65057 227896 240935 227898
rect 65057 227840 65062 227896
rect 65118 227840 240874 227896
rect 240930 227840 240935 227896
rect 65057 227838 240935 227840
rect 65057 227835 65123 227838
rect 240869 227835 240935 227838
rect 72417 227762 72483 227765
rect 271137 227762 271203 227765
rect 72417 227760 271203 227762
rect 72417 227704 72422 227760
rect 72478 227704 271142 227760
rect 271198 227704 271203 227760
rect 72417 227702 271203 227704
rect 72417 227699 72483 227702
rect 271137 227699 271203 227702
rect 113449 227626 113515 227629
rect 114461 227626 114527 227629
rect 113449 227624 114527 227626
rect 113449 227568 113454 227624
rect 113510 227568 114466 227624
rect 114522 227568 114527 227624
rect 113449 227566 114527 227568
rect 113449 227563 113515 227566
rect 114461 227563 114527 227566
rect 118969 227626 119035 227629
rect 119981 227626 120047 227629
rect 118969 227624 120047 227626
rect 118969 227568 118974 227624
rect 119030 227568 119986 227624
rect 120042 227568 120047 227624
rect 118969 227566 120047 227568
rect 118969 227563 119035 227566
rect 119981 227563 120047 227566
rect 219985 227354 220051 227357
rect 227253 227354 227319 227357
rect 219985 227352 227319 227354
rect 219985 227296 219990 227352
rect 220046 227296 227258 227352
rect 227314 227296 227319 227352
rect 219985 227294 227319 227296
rect 219985 227291 220051 227294
rect 227253 227291 227319 227294
rect 56777 227218 56843 227221
rect 61377 227218 61443 227221
rect 56777 227216 61443 227218
rect 56777 227160 56782 227216
rect 56838 227160 61382 227216
rect 61438 227160 61443 227216
rect 56777 227158 61443 227160
rect 56777 227155 56843 227158
rect 61377 227155 61443 227158
rect 219249 227218 219315 227221
rect 226793 227218 226859 227221
rect 219249 227216 226859 227218
rect 219249 227160 219254 227216
rect 219310 227160 226798 227216
rect 226854 227160 226859 227216
rect 219249 227158 226859 227160
rect 219249 227155 219315 227158
rect 226793 227155 226859 227158
rect 3693 227082 3759 227085
rect 70301 227082 70367 227085
rect 3693 227080 70367 227082
rect 3693 227024 3698 227080
rect 3754 227024 70306 227080
rect 70362 227024 70367 227080
rect 3693 227022 70367 227024
rect 3693 227019 3759 227022
rect 70301 227019 70367 227022
rect 74257 227082 74323 227085
rect 234337 227082 234403 227085
rect 74257 227080 234403 227082
rect 74257 227024 74262 227080
rect 74318 227024 234342 227080
rect 234398 227024 234403 227080
rect 74257 227022 234403 227024
rect 74257 227019 74323 227022
rect 234337 227019 234403 227022
rect 70025 226946 70091 226949
rect 235533 226946 235599 226949
rect 70025 226944 235599 226946
rect 70025 226888 70030 226944
rect 70086 226888 235538 226944
rect 235594 226888 235599 226944
rect 70025 226886 235599 226888
rect 70025 226883 70091 226886
rect 235533 226883 235599 226886
rect 59813 226810 59879 226813
rect 60181 226810 60247 226813
rect 59813 226808 60247 226810
rect 59813 226752 59818 226808
rect 59874 226752 60186 226808
rect 60242 226752 60247 226808
rect 59813 226750 60247 226752
rect 59813 226747 59879 226750
rect 60181 226747 60247 226750
rect 62665 226810 62731 226813
rect 234061 226810 234127 226813
rect 62665 226808 234127 226810
rect 62665 226752 62670 226808
rect 62726 226752 234066 226808
rect 234122 226752 234127 226808
rect 62665 226750 234127 226752
rect 62665 226747 62731 226750
rect 234061 226747 234127 226750
rect 56685 226674 56751 226677
rect 62941 226674 63007 226677
rect 56685 226672 63007 226674
rect 56685 226616 56690 226672
rect 56746 226616 62946 226672
rect 63002 226616 63007 226672
rect 56685 226614 63007 226616
rect 56685 226611 56751 226614
rect 62941 226611 63007 226614
rect 71681 226674 71747 226677
rect 246297 226674 246363 226677
rect 71681 226672 246363 226674
rect 71681 226616 71686 226672
rect 71742 226616 246302 226672
rect 246358 226616 246363 226672
rect 71681 226614 246363 226616
rect 71681 226611 71747 226614
rect 246297 226611 246363 226614
rect 61745 226538 61811 226541
rect 238109 226538 238175 226541
rect 61745 226536 238175 226538
rect 61745 226480 61750 226536
rect 61806 226480 238114 226536
rect 238170 226480 238175 226536
rect 61745 226478 238175 226480
rect 61745 226475 61811 226478
rect 238109 226475 238175 226478
rect 57881 226402 57947 226405
rect 62757 226402 62823 226405
rect 57881 226400 62823 226402
rect 57881 226344 57886 226400
rect 57942 226344 62762 226400
rect 62818 226344 62823 226400
rect 57881 226342 62823 226344
rect 57881 226339 57947 226342
rect 62757 226339 62823 226342
rect 68185 226402 68251 226405
rect 410517 226402 410583 226405
rect 68185 226400 410583 226402
rect 68185 226344 68190 226400
rect 68246 226344 410522 226400
rect 410578 226344 410583 226400
rect 68185 226342 410583 226344
rect 68185 226339 68251 226342
rect 410517 226339 410583 226342
rect 57053 226266 57119 226269
rect 61101 226266 61167 226269
rect 57053 226264 61167 226266
rect 57053 226208 57058 226264
rect 57114 226208 61106 226264
rect 61162 226208 61167 226264
rect 57053 226206 61167 226208
rect 57053 226203 57119 226206
rect 61101 226203 61167 226206
rect 62021 226266 62087 226269
rect 219341 226266 219407 226269
rect 62021 226264 62130 226266
rect 62021 226208 62026 226264
rect 62082 226208 62130 226264
rect 62021 226203 62130 226208
rect 219341 226264 219450 226266
rect 219341 226208 219346 226264
rect 219402 226208 219450 226264
rect 219341 226203 219450 226208
rect 62070 225858 62130 226203
rect 59862 225798 62130 225858
rect 219390 225858 219450 226203
rect 227069 225994 227135 225997
rect 222150 225992 227135 225994
rect 222150 225936 227074 225992
rect 227130 225936 227135 225992
rect 222150 225934 227135 225936
rect 222150 225858 222210 225934
rect 227069 225931 227135 225934
rect 219390 225798 222210 225858
rect 59862 225178 59922 225798
rect 224166 225796 224172 225860
rect 224236 225796 224242 225860
rect 224174 225556 224234 225796
rect 59862 225118 60076 225178
rect 224902 224980 224908 225044
rect 224972 225042 224978 225044
rect 225822 225042 225828 225044
rect 224972 224982 225828 225042
rect 224972 224980 224978 224982
rect 225822 224980 225828 224982
rect 225892 224980 225898 225044
rect 224861 223138 224927 223141
rect 224572 223136 224927 223138
rect 224572 223080 224866 223136
rect 224922 223080 224927 223136
rect 224572 223078 224927 223080
rect 224861 223075 224927 223078
rect 57513 222050 57579 222053
rect 57513 222048 60076 222050
rect 57513 221992 57518 222048
rect 57574 221992 60076 222048
rect 57513 221990 60076 221992
rect 57513 221987 57579 221990
rect 225505 220690 225571 220693
rect 224572 220688 225571 220690
rect 224572 220632 225510 220688
rect 225566 220632 225571 220688
rect 224572 220630 225571 220632
rect 225505 220627 225571 220630
rect 583520 219058 584960 219148
rect 583342 218998 584960 219058
rect 58157 218922 58223 218925
rect 583342 218922 583402 218998
rect 583520 218922 584960 218998
rect 58157 218920 60076 218922
rect 58157 218864 58162 218920
rect 58218 218864 60076 218920
rect 58157 218862 60076 218864
rect 583342 218908 584960 218922
rect 583342 218862 583586 218908
rect 58157 218859 58223 218862
rect 229921 218242 229987 218245
rect 224572 218240 229987 218242
rect 224572 218184 229926 218240
rect 229982 218184 229987 218240
rect 224572 218182 229987 218184
rect 229921 218179 229987 218182
rect 234429 218106 234495 218109
rect 583526 218106 583586 218862
rect 234429 218104 583586 218106
rect 234429 218048 234434 218104
rect 234490 218048 583586 218104
rect 234429 218046 583586 218048
rect 234429 218043 234495 218046
rect 56409 215794 56475 215797
rect 227621 215794 227687 215797
rect 56409 215792 60076 215794
rect 56409 215736 56414 215792
rect 56470 215736 60076 215792
rect 56409 215734 60076 215736
rect 224572 215792 227687 215794
rect 224572 215736 227626 215792
rect 227682 215736 227687 215792
rect 224572 215734 227687 215736
rect 56409 215731 56475 215734
rect 227621 215731 227687 215734
rect -960 214978 480 215068
rect 3049 214978 3115 214981
rect -960 214976 3115 214978
rect -960 214920 3054 214976
rect 3110 214920 3115 214976
rect -960 214918 3115 214920
rect -960 214828 480 214918
rect 3049 214915 3115 214918
rect 226149 213346 226215 213349
rect 224572 213344 226215 213346
rect 224572 213288 226154 213344
rect 226210 213288 226215 213344
rect 224572 213286 226215 213288
rect 226149 213283 226215 213286
rect 57513 212666 57579 212669
rect 57513 212664 60076 212666
rect 57513 212608 57518 212664
rect 57574 212608 60076 212664
rect 57513 212606 60076 212608
rect 57513 212603 57579 212606
rect 227989 210898 228055 210901
rect 224572 210896 228055 210898
rect 224572 210840 227994 210896
rect 228050 210840 228055 210896
rect 224572 210838 228055 210840
rect 227989 210835 228055 210838
rect 227621 209674 227687 209677
rect 235257 209674 235323 209677
rect 227621 209672 235323 209674
rect 227621 209616 227626 209672
rect 227682 209616 235262 209672
rect 235318 209616 235323 209672
rect 227621 209614 235323 209616
rect 227621 209611 227687 209614
rect 235257 209611 235323 209614
rect 57881 209538 57947 209541
rect 57881 209536 60076 209538
rect 57881 209480 57886 209536
rect 57942 209480 60076 209536
rect 57881 209478 60076 209480
rect 57881 209475 57947 209478
rect 227621 208450 227687 208453
rect 224572 208448 227687 208450
rect 224572 208392 227626 208448
rect 227682 208392 227687 208448
rect 224572 208390 227687 208392
rect 227621 208387 227687 208390
rect 55857 206274 55923 206277
rect 55857 206272 60076 206274
rect 55857 206216 55862 206272
rect 55918 206216 60076 206272
rect 55857 206214 60076 206216
rect 55857 206211 55923 206214
rect 231393 206002 231459 206005
rect 224572 206000 231459 206002
rect 224572 205944 231398 206000
rect 231454 205944 231459 206000
rect 224572 205942 231459 205944
rect 231393 205939 231459 205942
rect 234337 205730 234403 205733
rect 583520 205730 584960 205820
rect 234337 205728 584960 205730
rect 234337 205672 234342 205728
rect 234398 205672 584960 205728
rect 234337 205670 584960 205672
rect 234337 205667 234403 205670
rect 583520 205580 584960 205670
rect 229829 203554 229895 203557
rect 224572 203552 229895 203554
rect 224572 203496 229834 203552
rect 229890 203496 229895 203552
rect 224572 203494 229895 203496
rect 229829 203491 229895 203494
rect 59537 203146 59603 203149
rect 59537 203144 60076 203146
rect 59537 203088 59542 203144
rect 59598 203088 60076 203144
rect 59537 203086 60076 203088
rect 59537 203083 59603 203086
rect -960 201922 480 202012
rect 3785 201922 3851 201925
rect -960 201920 3851 201922
rect -960 201864 3790 201920
rect 3846 201864 3851 201920
rect -960 201862 3851 201864
rect -960 201772 480 201862
rect 3785 201859 3851 201862
rect 238293 201106 238359 201109
rect 224572 201104 238359 201106
rect 224572 201048 238298 201104
rect 238354 201048 238359 201104
rect 224572 201046 238359 201048
rect 238293 201043 238359 201046
rect 58709 200018 58775 200021
rect 58709 200016 60076 200018
rect 58709 199960 58714 200016
rect 58770 199960 60076 200016
rect 58709 199958 60076 199960
rect 58709 199955 58775 199958
rect 225229 198658 225295 198661
rect 224572 198656 225295 198658
rect 224572 198600 225234 198656
rect 225290 198600 225295 198656
rect 224572 198598 225295 198600
rect 225229 198595 225295 198598
rect 57513 196890 57579 196893
rect 57513 196888 60076 196890
rect 57513 196832 57518 196888
rect 57574 196832 60076 196888
rect 57513 196830 60076 196832
rect 57513 196827 57579 196830
rect 227529 196210 227595 196213
rect 224572 196208 227595 196210
rect 224572 196152 227534 196208
rect 227590 196152 227595 196208
rect 224572 196150 227595 196152
rect 227529 196147 227595 196150
rect 57513 193762 57579 193765
rect 225137 193762 225203 193765
rect 57513 193760 60076 193762
rect 57513 193704 57518 193760
rect 57574 193704 60076 193760
rect 57513 193702 60076 193704
rect 224572 193760 225203 193762
rect 224572 193704 225142 193760
rect 225198 193704 225203 193760
rect 224572 193702 225203 193704
rect 57513 193699 57579 193702
rect 225137 193699 225203 193702
rect 580165 192538 580231 192541
rect 583520 192538 584960 192628
rect 580165 192536 584960 192538
rect 580165 192480 580170 192536
rect 580226 192480 584960 192536
rect 580165 192478 584960 192480
rect 580165 192475 580231 192478
rect 583520 192388 584960 192478
rect 234245 191314 234311 191317
rect 224572 191312 234311 191314
rect 224572 191256 234250 191312
rect 234306 191256 234311 191312
rect 224572 191254 234311 191256
rect 234245 191251 234311 191254
rect 57513 190634 57579 190637
rect 57513 190632 60076 190634
rect 57513 190576 57518 190632
rect 57574 190576 60076 190632
rect 57513 190574 60076 190576
rect 57513 190571 57579 190574
rect -960 188866 480 188956
rect 3325 188866 3391 188869
rect 227345 188866 227411 188869
rect -960 188864 3391 188866
rect -960 188808 3330 188864
rect 3386 188808 3391 188864
rect -960 188806 3391 188808
rect 224572 188864 227411 188866
rect 224572 188808 227350 188864
rect 227406 188808 227411 188864
rect 224572 188806 227411 188808
rect -960 188716 480 188806
rect 3325 188803 3391 188806
rect 227345 188803 227411 188806
rect 57053 187506 57119 187509
rect 57053 187504 60076 187506
rect 57053 187448 57058 187504
rect 57114 187448 60076 187504
rect 57053 187446 60076 187448
rect 57053 187443 57119 187446
rect 228633 186418 228699 186421
rect 224572 186416 228699 186418
rect 224572 186360 228638 186416
rect 228694 186360 228699 186416
rect 224572 186358 228699 186360
rect 228633 186355 228699 186358
rect 56317 184242 56383 184245
rect 56317 184240 60076 184242
rect 56317 184184 56322 184240
rect 56378 184184 60076 184240
rect 56317 184182 60076 184184
rect 56317 184179 56383 184182
rect 226701 183970 226767 183973
rect 224572 183968 226767 183970
rect 224572 183912 226706 183968
rect 226762 183912 226767 183968
rect 224572 183910 226767 183912
rect 226701 183907 226767 183910
rect 227437 181522 227503 181525
rect 224572 181520 227503 181522
rect 224572 181464 227442 181520
rect 227498 181464 227503 181520
rect 224572 181462 227503 181464
rect 227437 181459 227503 181462
rect 57513 181114 57579 181117
rect 57513 181112 60076 181114
rect 57513 181056 57518 181112
rect 57574 181056 60076 181112
rect 57513 181054 60076 181056
rect 57513 181051 57579 181054
rect 583520 179210 584960 179300
rect 583342 179150 584960 179210
rect 227805 179074 227871 179077
rect 224572 179072 227871 179074
rect 224572 179016 227810 179072
rect 227866 179016 227871 179072
rect 224572 179014 227871 179016
rect 583342 179074 583402 179150
rect 583520 179074 584960 179150
rect 583342 179060 584960 179074
rect 583342 179014 583586 179060
rect 227805 179011 227871 179014
rect 236729 178122 236795 178125
rect 583526 178122 583586 179014
rect 236729 178120 583586 178122
rect 236729 178064 236734 178120
rect 236790 178064 583586 178120
rect 236729 178062 583586 178064
rect 236729 178059 236795 178062
rect 57513 177986 57579 177989
rect 57513 177984 60076 177986
rect 57513 177928 57518 177984
rect 57574 177928 60076 177984
rect 57513 177926 60076 177928
rect 57513 177923 57579 177926
rect 226609 176626 226675 176629
rect 224572 176624 226675 176626
rect 224572 176568 226614 176624
rect 226670 176568 226675 176624
rect 224572 176566 226675 176568
rect 226609 176563 226675 176566
rect -960 175796 480 176036
rect 226609 175266 226675 175269
rect 234153 175266 234219 175269
rect 226609 175264 234219 175266
rect 226609 175208 226614 175264
rect 226670 175208 234158 175264
rect 234214 175208 234219 175264
rect 226609 175206 234219 175208
rect 226609 175203 226675 175206
rect 234153 175203 234219 175206
rect 57513 174858 57579 174861
rect 57513 174856 60076 174858
rect 57513 174800 57518 174856
rect 57574 174800 60076 174856
rect 57513 174798 60076 174800
rect 57513 174795 57579 174798
rect 226609 174178 226675 174181
rect 224572 174176 226675 174178
rect 224572 174120 226614 174176
rect 226670 174120 226675 174176
rect 224572 174118 226675 174120
rect 226609 174115 226675 174118
rect 59445 171730 59511 171733
rect 59445 171728 60076 171730
rect 59445 171672 59450 171728
rect 59506 171672 60076 171728
rect 59445 171670 60076 171672
rect 59445 171667 59511 171670
rect 227161 171594 227227 171597
rect 224572 171592 227227 171594
rect 224572 171536 227166 171592
rect 227222 171536 227227 171592
rect 224572 171534 227227 171536
rect 227161 171531 227227 171534
rect 228541 169146 228607 169149
rect 224572 169144 228607 169146
rect 224572 169088 228546 169144
rect 228602 169088 228607 169144
rect 224572 169086 228607 169088
rect 228541 169083 228607 169086
rect 58801 168602 58867 168605
rect 58801 168600 60076 168602
rect 58801 168544 58806 168600
rect 58862 168544 60076 168600
rect 58801 168542 60076 168544
rect 58801 168539 58867 168542
rect 227253 166698 227319 166701
rect 224572 166696 227319 166698
rect 224572 166640 227258 166696
rect 227314 166640 227319 166696
rect 224572 166638 227319 166640
rect 227253 166635 227319 166638
rect 583520 165882 584960 165972
rect 567150 165822 584960 165882
rect 246297 165746 246363 165749
rect 567150 165746 567210 165822
rect 246297 165744 567210 165746
rect 246297 165688 246302 165744
rect 246358 165688 567210 165744
rect 583520 165732 584960 165822
rect 246297 165686 567210 165688
rect 246297 165683 246363 165686
rect 56501 165338 56567 165341
rect 56501 165336 60076 165338
rect 56501 165280 56506 165336
rect 56562 165280 60076 165336
rect 56501 165278 60076 165280
rect 56501 165275 56567 165278
rect 226057 164250 226123 164253
rect 224572 164248 226123 164250
rect 224572 164192 226062 164248
rect 226118 164192 226123 164248
rect 224572 164190 226123 164192
rect 226057 164187 226123 164190
rect -960 162890 480 162980
rect 3049 162890 3115 162893
rect -960 162888 3115 162890
rect -960 162832 3054 162888
rect 3110 162832 3115 162888
rect -960 162830 3115 162832
rect -960 162740 480 162830
rect 3049 162827 3115 162830
rect 58065 162210 58131 162213
rect 58065 162208 60076 162210
rect 58065 162152 58070 162208
rect 58126 162152 60076 162208
rect 58065 162150 60076 162152
rect 58065 162147 58131 162150
rect 231301 161802 231367 161805
rect 224572 161800 231367 161802
rect 224572 161744 231306 161800
rect 231362 161744 231367 161800
rect 224572 161742 231367 161744
rect 231301 161739 231367 161742
rect 226517 159354 226583 159357
rect 224572 159352 226583 159354
rect 224572 159296 226522 159352
rect 226578 159296 226583 159352
rect 224572 159294 226583 159296
rect 226517 159291 226583 159294
rect 57421 159082 57487 159085
rect 57421 159080 60076 159082
rect 57421 159024 57426 159080
rect 57482 159024 60076 159080
rect 57421 159022 60076 159024
rect 57421 159019 57487 159022
rect 240777 157314 240843 157317
rect 229050 157312 240843 157314
rect 229050 157256 240782 157312
rect 240838 157256 240843 157312
rect 229050 157254 240843 157256
rect 229050 156906 229110 157254
rect 240777 157251 240843 157254
rect 224572 156846 229110 156906
rect 57513 155954 57579 155957
rect 57513 155952 60076 155954
rect 57513 155896 57518 155952
rect 57574 155896 60076 155952
rect 57513 155894 60076 155896
rect 57513 155891 57579 155894
rect 226885 154458 226951 154461
rect 224572 154456 226951 154458
rect 224572 154400 226890 154456
rect 226946 154400 226951 154456
rect 224572 154398 226951 154400
rect 226885 154395 226951 154398
rect 57513 152826 57579 152829
rect 57513 152824 60076 152826
rect 57513 152768 57518 152824
rect 57574 152768 60076 152824
rect 57513 152766 60076 152768
rect 57513 152763 57579 152766
rect 583520 152690 584960 152780
rect 583342 152630 584960 152690
rect 583342 152554 583402 152630
rect 583520 152554 584960 152630
rect 583342 152540 584960 152554
rect 583342 152494 583586 152540
rect 225965 152010 226031 152013
rect 224572 152008 226031 152010
rect 224572 151952 225970 152008
rect 226026 151952 226031 152008
rect 224572 151950 226031 151952
rect 225965 151947 226031 151950
rect 235533 151874 235599 151877
rect 583526 151874 583586 152494
rect 235533 151872 583586 151874
rect 235533 151816 235538 151872
rect 235594 151816 583586 151872
rect 235533 151814 583586 151816
rect 235533 151811 235599 151814
rect 226517 150378 226583 150381
rect 235441 150378 235507 150381
rect 226517 150376 235507 150378
rect 226517 150320 226522 150376
rect 226578 150320 235446 150376
rect 235502 150320 235507 150376
rect 226517 150318 235507 150320
rect 226517 150315 226583 150318
rect 235441 150315 235507 150318
rect -960 149834 480 149924
rect 3693 149834 3759 149837
rect -960 149832 3759 149834
rect -960 149776 3698 149832
rect 3754 149776 3759 149832
rect -960 149774 3759 149776
rect -960 149684 480 149774
rect 3693 149771 3759 149774
rect 56777 149698 56843 149701
rect 56777 149696 60076 149698
rect 56777 149640 56782 149696
rect 56838 149640 60076 149696
rect 56777 149638 60076 149640
rect 56777 149635 56843 149638
rect 226517 149562 226583 149565
rect 224572 149560 226583 149562
rect 224572 149504 226522 149560
rect 226578 149504 226583 149560
rect 224572 149502 226583 149504
rect 226517 149499 226583 149502
rect 229645 147114 229711 147117
rect 224572 147112 229711 147114
rect 224572 147056 229650 147112
rect 229706 147056 229711 147112
rect 224572 147054 229711 147056
rect 229645 147051 229711 147054
rect 57421 146570 57487 146573
rect 57421 146568 60076 146570
rect 57421 146512 57426 146568
rect 57482 146512 60076 146568
rect 57421 146510 60076 146512
rect 57421 146507 57487 146510
rect 226977 144666 227043 144669
rect 224572 144664 227043 144666
rect 224572 144608 226982 144664
rect 227038 144608 227043 144664
rect 224572 144606 227043 144608
rect 226977 144603 227043 144606
rect 57513 143306 57579 143309
rect 57513 143304 60076 143306
rect 57513 143248 57518 143304
rect 57574 143248 60076 143304
rect 57513 143246 60076 143248
rect 57513 143243 57579 143246
rect 227069 142218 227135 142221
rect 224572 142216 227135 142218
rect 224572 142160 227074 142216
rect 227130 142160 227135 142216
rect 224572 142158 227135 142160
rect 227069 142155 227135 142158
rect 226517 140722 226583 140725
rect 232497 140722 232563 140725
rect 226517 140720 232563 140722
rect 226517 140664 226522 140720
rect 226578 140664 232502 140720
rect 232558 140664 232563 140720
rect 226517 140662 232563 140664
rect 226517 140659 226583 140662
rect 232497 140659 232563 140662
rect 58617 140178 58683 140181
rect 58617 140176 60076 140178
rect 58617 140120 58622 140176
rect 58678 140120 60076 140176
rect 58617 140118 60076 140120
rect 58617 140115 58683 140118
rect 226517 139770 226583 139773
rect 224572 139768 226583 139770
rect 224572 139712 226522 139768
rect 226578 139712 226583 139768
rect 224572 139710 226583 139712
rect 226517 139707 226583 139710
rect 583520 139362 584960 139452
rect 583342 139302 584960 139362
rect 583342 139226 583402 139302
rect 583520 139226 584960 139302
rect 583342 139212 584960 139226
rect 583342 139166 583586 139212
rect 239397 138138 239463 138141
rect 583526 138138 583586 139166
rect 239397 138136 583586 138138
rect 239397 138080 239402 138136
rect 239458 138080 583586 138136
rect 239397 138078 583586 138080
rect 239397 138075 239463 138078
rect 232313 137322 232379 137325
rect 224572 137320 232379 137322
rect 224572 137264 232318 137320
rect 232374 137264 232379 137320
rect 224572 137262 232379 137264
rect 232313 137259 232379 137262
rect 56041 137050 56107 137053
rect 56041 137048 60076 137050
rect 56041 136992 56046 137048
rect 56102 136992 60076 137048
rect 56041 136990 60076 136992
rect 56041 136987 56107 136990
rect -960 136778 480 136868
rect 3049 136778 3115 136781
rect -960 136776 3115 136778
rect -960 136720 3054 136776
rect 3110 136720 3115 136776
rect -960 136718 3115 136720
rect -960 136628 480 136718
rect 3049 136715 3115 136718
rect 225873 134874 225939 134877
rect 224572 134872 225939 134874
rect 224572 134816 225878 134872
rect 225934 134816 225939 134872
rect 224572 134814 225939 134816
rect 225873 134811 225939 134814
rect 57421 133922 57487 133925
rect 57421 133920 60076 133922
rect 57421 133864 57426 133920
rect 57482 133864 60076 133920
rect 57421 133862 60076 133864
rect 57421 133859 57487 133862
rect 249057 132426 249123 132429
rect 224572 132424 249123 132426
rect 224572 132368 249062 132424
rect 249118 132368 249123 132424
rect 224572 132366 249123 132368
rect 249057 132363 249123 132366
rect 57605 130794 57671 130797
rect 57605 130792 60076 130794
rect 57605 130736 57610 130792
rect 57666 130736 60076 130792
rect 57605 130734 60076 130736
rect 57605 130731 57671 130734
rect 232221 129978 232287 129981
rect 224572 129976 232287 129978
rect 224572 129920 232226 129976
rect 232282 129920 232287 129976
rect 224572 129918 232287 129920
rect 232221 129915 232287 129918
rect 58985 127666 59051 127669
rect 58985 127664 60076 127666
rect 58985 127608 58990 127664
rect 59046 127608 60076 127664
rect 58985 127606 60076 127608
rect 58985 127603 59051 127606
rect 232129 127530 232195 127533
rect 224572 127528 232195 127530
rect 224572 127472 232134 127528
rect 232190 127472 232195 127528
rect 224572 127470 232195 127472
rect 232129 127467 232195 127470
rect 583520 126034 584960 126124
rect 583342 125974 584960 126034
rect 583342 125898 583402 125974
rect 583520 125898 584960 125974
rect 583342 125884 584960 125898
rect 583342 125838 583586 125884
rect 236637 125626 236703 125629
rect 583526 125626 583586 125838
rect 236637 125624 583586 125626
rect 236637 125568 236642 125624
rect 236698 125568 583586 125624
rect 236637 125566 583586 125568
rect 236637 125563 236703 125566
rect 238017 125082 238083 125085
rect 224572 125080 238083 125082
rect 224572 125024 238022 125080
rect 238078 125024 238083 125080
rect 224572 125022 238083 125024
rect 238017 125019 238083 125022
rect 58249 124538 58315 124541
rect 58249 124536 60076 124538
rect 58249 124480 58254 124536
rect 58310 124480 60076 124536
rect 58249 124478 60076 124480
rect 58249 124475 58315 124478
rect -960 123572 480 123812
rect 232037 122634 232103 122637
rect 224572 122632 232103 122634
rect 224572 122576 232042 122632
rect 232098 122576 232103 122632
rect 224572 122574 232103 122576
rect 232037 122571 232103 122574
rect 55949 121274 56015 121277
rect 55949 121272 60076 121274
rect 55949 121216 55954 121272
rect 56010 121216 60076 121272
rect 55949 121214 60076 121216
rect 55949 121211 56015 121214
rect 235257 120730 235323 120733
rect 241513 120730 241579 120733
rect 235257 120728 241579 120730
rect 235257 120672 235262 120728
rect 235318 120672 241518 120728
rect 241574 120672 241579 120728
rect 235257 120670 241579 120672
rect 235257 120667 235323 120670
rect 241513 120667 241579 120670
rect 226425 120186 226491 120189
rect 224572 120184 226491 120186
rect 224572 120128 226430 120184
rect 226486 120128 226491 120184
rect 224572 120126 226491 120128
rect 226425 120123 226491 120126
rect 57605 118146 57671 118149
rect 57605 118144 60076 118146
rect 57605 118088 57610 118144
rect 57666 118088 60076 118144
rect 57605 118086 60076 118088
rect 57605 118083 57671 118086
rect 229737 117738 229803 117741
rect 224572 117736 229803 117738
rect 224572 117680 229742 117736
rect 229798 117680 229803 117736
rect 224572 117678 229803 117680
rect 229737 117675 229803 117678
rect 226374 115154 226380 115156
rect 224572 115094 226380 115154
rect 226374 115092 226380 115094
rect 226444 115092 226450 115156
rect 58341 115018 58407 115021
rect 58341 115016 60076 115018
rect 58341 114960 58346 115016
rect 58402 114960 60076 115016
rect 58341 114958 60076 114960
rect 58341 114955 58407 114958
rect 583520 112842 584960 112932
rect 583342 112782 584960 112842
rect 228449 112706 228515 112709
rect 224572 112704 228515 112706
rect 224572 112648 228454 112704
rect 228510 112648 228515 112704
rect 224572 112646 228515 112648
rect 583342 112706 583402 112782
rect 583520 112706 584960 112782
rect 583342 112692 584960 112706
rect 583342 112646 583586 112692
rect 228449 112643 228515 112646
rect 57605 111890 57671 111893
rect 253289 111890 253355 111893
rect 583526 111890 583586 112646
rect 57605 111888 60076 111890
rect 57605 111832 57610 111888
rect 57666 111832 60076 111888
rect 57605 111830 60076 111832
rect 253289 111888 583586 111890
rect 253289 111832 253294 111888
rect 253350 111832 583586 111888
rect 253289 111830 583586 111832
rect 57605 111827 57671 111830
rect 253289 111827 253355 111830
rect -960 110666 480 110756
rect 3325 110666 3391 110669
rect -960 110664 3391 110666
rect -960 110608 3330 110664
rect 3386 110608 3391 110664
rect -960 110606 3391 110608
rect -960 110516 480 110606
rect 3325 110603 3391 110606
rect 233969 110258 234035 110261
rect 224572 110256 234035 110258
rect 224572 110200 233974 110256
rect 234030 110200 234035 110256
rect 224572 110198 234035 110200
rect 233969 110195 234035 110198
rect 56133 108762 56199 108765
rect 56133 108760 60076 108762
rect 56133 108704 56138 108760
rect 56194 108704 60076 108760
rect 56133 108702 60076 108704
rect 56133 108699 56199 108702
rect 226742 107810 226748 107812
rect 224572 107750 226748 107810
rect 226742 107748 226748 107750
rect 226812 107748 226818 107812
rect 56593 105634 56659 105637
rect 56593 105632 60076 105634
rect 56593 105576 56598 105632
rect 56654 105576 60076 105632
rect 56593 105574 60076 105576
rect 56593 105571 56659 105574
rect 228357 105362 228423 105365
rect 224572 105360 228423 105362
rect 224572 105304 228362 105360
rect 228418 105304 228423 105360
rect 224572 105302 228423 105304
rect 228357 105299 228423 105302
rect 238201 102914 238267 102917
rect 224572 102912 238267 102914
rect 224572 102856 238206 102912
rect 238262 102856 238267 102912
rect 224572 102854 238267 102856
rect 238201 102851 238267 102854
rect 57145 102370 57211 102373
rect 57145 102368 60076 102370
rect 57145 102312 57150 102368
rect 57206 102312 60076 102368
rect 57145 102310 60076 102312
rect 57145 102307 57211 102310
rect 235257 100466 235323 100469
rect 224572 100464 235323 100466
rect 224572 100408 235262 100464
rect 235318 100408 235323 100464
rect 224572 100406 235323 100408
rect 235257 100403 235323 100406
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect 59077 99242 59143 99245
rect 59077 99240 60076 99242
rect 59077 99184 59082 99240
rect 59138 99184 60076 99240
rect 59077 99182 60076 99184
rect 59077 99179 59143 99182
rect 231945 98018 232011 98021
rect 224572 98016 232011 98018
rect 224572 97960 231950 98016
rect 232006 97960 232011 98016
rect 224572 97958 232011 97960
rect 231945 97955 232011 97958
rect -960 97610 480 97700
rect 3233 97610 3299 97613
rect -960 97608 3299 97610
rect -960 97552 3238 97608
rect 3294 97552 3299 97608
rect -960 97550 3299 97552
rect -960 97460 480 97550
rect 3233 97547 3299 97550
rect 57237 96114 57303 96117
rect 57237 96112 60076 96114
rect 57237 96056 57242 96112
rect 57298 96056 60076 96112
rect 57237 96054 60076 96056
rect 57237 96051 57303 96054
rect 233233 95570 233299 95573
rect 224572 95568 233299 95570
rect 224572 95512 233238 95568
rect 233294 95512 233299 95568
rect 224572 95510 233299 95512
rect 233233 95507 233299 95510
rect 225597 93122 225663 93125
rect 224572 93120 225663 93122
rect 224572 93064 225602 93120
rect 225658 93064 225663 93120
rect 224572 93062 225663 93064
rect 225597 93059 225663 93062
rect 59169 92986 59235 92989
rect 59169 92984 60076 92986
rect 59169 92928 59174 92984
rect 59230 92928 60076 92984
rect 59169 92926 60076 92928
rect 59169 92923 59235 92926
rect 242249 91082 242315 91085
rect 229050 91080 242315 91082
rect 229050 91024 242254 91080
rect 242310 91024 242315 91080
rect 229050 91022 242315 91024
rect 229050 90674 229110 91022
rect 242249 91019 242315 91022
rect 224572 90614 229110 90674
rect 57329 89858 57395 89861
rect 57329 89856 60076 89858
rect 57329 89800 57334 89856
rect 57390 89800 60076 89856
rect 57329 89798 60076 89800
rect 57329 89795 57395 89798
rect 226333 88226 226399 88229
rect 224572 88224 226399 88226
rect 224572 88168 226338 88224
rect 226394 88168 226399 88224
rect 224572 88166 226399 88168
rect 226333 88163 226399 88166
rect 57421 86730 57487 86733
rect 57421 86728 60076 86730
rect 57421 86672 57426 86728
rect 57482 86672 60076 86728
rect 57421 86670 60076 86672
rect 57421 86667 57487 86670
rect 583520 86186 584960 86276
rect 583342 86126 584960 86186
rect 583342 86050 583402 86126
rect 583520 86050 584960 86126
rect 583342 86036 584960 86050
rect 583342 85990 583586 86036
rect 231853 85778 231919 85781
rect 224572 85776 231919 85778
rect 224572 85720 231858 85776
rect 231914 85720 231919 85776
rect 224572 85718 231919 85720
rect 231853 85715 231919 85718
rect 235349 85642 235415 85645
rect 583526 85642 583586 85990
rect 235349 85640 583586 85642
rect 235349 85584 235354 85640
rect 235410 85584 583586 85640
rect 235349 85582 583586 85584
rect 235349 85579 235415 85582
rect -960 84690 480 84780
rect 2957 84690 3023 84693
rect -960 84688 3023 84690
rect -960 84632 2962 84688
rect 3018 84632 3023 84688
rect -960 84630 3023 84632
rect -960 84540 480 84630
rect 2957 84627 3023 84630
rect 226517 84146 226583 84149
rect 242157 84146 242223 84149
rect 226517 84144 242223 84146
rect 226517 84088 226522 84144
rect 226578 84088 242162 84144
rect 242218 84088 242223 84144
rect 226517 84086 242223 84088
rect 226517 84083 226583 84086
rect 242157 84083 242223 84086
rect 56225 83602 56291 83605
rect 56225 83600 60076 83602
rect 56225 83544 56230 83600
rect 56286 83544 60076 83600
rect 56225 83542 60076 83544
rect 56225 83539 56291 83542
rect 226517 83330 226583 83333
rect 224572 83328 226583 83330
rect 224572 83272 226522 83328
rect 226578 83272 226583 83328
rect 224572 83270 226583 83272
rect 226517 83267 226583 83270
rect 226926 80882 226932 80884
rect 224572 80822 226932 80882
rect 226926 80820 226932 80822
rect 226996 80820 227002 80884
rect 59261 80338 59327 80341
rect 59261 80336 60076 80338
rect 59261 80280 59266 80336
rect 59322 80280 60076 80336
rect 59261 80278 60076 80280
rect 59261 80275 59327 80278
rect 231117 78434 231183 78437
rect 224572 78432 231183 78434
rect 224572 78376 231122 78432
rect 231178 78376 231183 78432
rect 224572 78374 231183 78376
rect 231117 78371 231183 78374
rect 56685 77210 56751 77213
rect 226517 77210 226583 77213
rect 356513 77210 356579 77213
rect 56685 77208 60076 77210
rect 56685 77152 56690 77208
rect 56746 77152 60076 77208
rect 56685 77150 60076 77152
rect 226517 77208 356579 77210
rect 226517 77152 226522 77208
rect 226578 77152 356518 77208
rect 356574 77152 356579 77208
rect 226517 77150 356579 77152
rect 56685 77147 56751 77150
rect 226517 77147 226583 77150
rect 356513 77147 356579 77150
rect 226517 75986 226583 75989
rect 224572 75984 226583 75986
rect 224572 75928 226522 75984
rect 226578 75928 226583 75984
rect 224572 75926 226583 75928
rect 226517 75923 226583 75926
rect 57697 74082 57763 74085
rect 57697 74080 60076 74082
rect 57697 74024 57702 74080
rect 57758 74024 60076 74080
rect 57697 74022 60076 74024
rect 57697 74019 57763 74022
rect 226558 73538 226564 73540
rect 224572 73478 226564 73538
rect 226558 73476 226564 73478
rect 226628 73476 226634 73540
rect 580349 72994 580415 72997
rect 583520 72994 584960 73084
rect 580349 72992 584960 72994
rect 580349 72936 580354 72992
rect 580410 72936 584960 72992
rect 580349 72934 584960 72936
rect 580349 72931 580415 72934
rect 583520 72844 584960 72934
rect -960 71634 480 71724
rect 3325 71634 3391 71637
rect -960 71632 3391 71634
rect -960 71576 3330 71632
rect 3386 71576 3391 71632
rect -960 71574 3391 71576
rect -960 71484 480 71574
rect 3325 71571 3391 71574
rect 226793 71090 226859 71093
rect 224572 71088 226859 71090
rect 224572 71032 226798 71088
rect 226854 71032 226859 71088
rect 224572 71030 226859 71032
rect 226793 71027 226859 71030
rect 57605 70954 57671 70957
rect 57605 70952 60076 70954
rect 57605 70896 57610 70952
rect 57666 70896 60076 70952
rect 57605 70894 60076 70896
rect 57605 70891 57671 70894
rect 227897 68642 227963 68645
rect 224572 68640 227963 68642
rect 224572 68584 227902 68640
rect 227958 68584 227963 68640
rect 224572 68582 227963 68584
rect 227897 68579 227963 68582
rect 58893 67826 58959 67829
rect 58893 67824 60076 67826
rect 58893 67768 58898 67824
rect 58954 67768 60076 67824
rect 58893 67766 60076 67768
rect 58893 67763 58959 67766
rect 232405 66194 232471 66197
rect 224572 66192 232471 66194
rect 224572 66136 232410 66192
rect 232466 66136 232471 66192
rect 224572 66134 232471 66136
rect 232405 66131 232471 66134
rect 226517 64834 226583 64837
rect 244917 64834 244983 64837
rect 226517 64832 244983 64834
rect 226517 64776 226522 64832
rect 226578 64776 244922 64832
rect 244978 64776 244983 64832
rect 226517 64774 244983 64776
rect 226517 64771 226583 64774
rect 244917 64771 244983 64774
rect 56869 64698 56935 64701
rect 56869 64696 60076 64698
rect 56869 64640 56874 64696
rect 56930 64640 60076 64696
rect 56869 64638 60076 64640
rect 56869 64635 56935 64638
rect 226517 63746 226583 63749
rect 224572 63744 226583 63746
rect 224572 63688 226522 63744
rect 226578 63688 226583 63744
rect 224572 63686 226583 63688
rect 226517 63683 226583 63686
rect 57053 61570 57119 61573
rect 57053 61568 60076 61570
rect 57053 61512 57058 61568
rect 57114 61512 60076 61568
rect 57053 61510 60076 61512
rect 57053 61507 57119 61510
rect 230749 61298 230815 61301
rect 224572 61296 230815 61298
rect 224572 61240 230754 61296
rect 230810 61240 230815 61296
rect 224572 61238 230815 61240
rect 230749 61235 230815 61238
rect 230933 60210 230999 60213
rect 223254 60208 230999 60210
rect 223254 60152 230938 60208
rect 230994 60152 230999 60208
rect 223254 60150 230999 60152
rect 223062 60074 223068 60076
rect 221598 60014 223068 60074
rect 218237 59938 218303 59941
rect 221598 59938 221658 60014
rect 223062 60012 223068 60014
rect 223132 60012 223138 60076
rect 218237 59936 221658 59938
rect 218237 59880 218242 59936
rect 218298 59880 221658 59936
rect 218237 59878 221658 59880
rect 222377 59938 222443 59941
rect 223254 59938 223314 60150
rect 230933 60147 230999 60150
rect 223430 60012 223436 60076
rect 223500 60074 223506 60076
rect 225086 60074 225092 60076
rect 223500 60014 225092 60074
rect 223500 60012 223506 60014
rect 225086 60012 225092 60014
rect 225156 60012 225162 60076
rect 222377 59936 223314 59938
rect 222377 59880 222382 59936
rect 222438 59880 223314 59936
rect 222377 59878 223314 59880
rect 218237 59875 218303 59878
rect 222377 59875 222443 59878
rect 223614 59876 223620 59940
rect 223684 59938 223690 59940
rect 223941 59938 224007 59941
rect 223684 59936 224007 59938
rect 223684 59880 223946 59936
rect 224002 59880 224007 59936
rect 223684 59878 224007 59880
rect 223684 59876 223690 59878
rect 223941 59875 224007 59878
rect 224125 59938 224191 59941
rect 226006 59938 226012 59940
rect 224125 59936 226012 59938
rect 224125 59880 224130 59936
rect 224186 59880 226012 59936
rect 224125 59878 226012 59880
rect 224125 59875 224191 59878
rect 226006 59876 226012 59878
rect 226076 59876 226082 59940
rect 216121 59802 216187 59805
rect 222561 59802 222627 59805
rect 216121 59800 222627 59802
rect 216121 59744 216126 59800
rect 216182 59744 222566 59800
rect 222622 59744 222627 59800
rect 216121 59742 222627 59744
rect 216121 59739 216187 59742
rect 222561 59739 222627 59742
rect 222745 59802 222811 59805
rect 223798 59802 223804 59804
rect 222745 59800 223804 59802
rect 222745 59744 222750 59800
rect 222806 59744 223804 59800
rect 222745 59742 223804 59744
rect 222745 59739 222811 59742
rect 223798 59740 223804 59742
rect 223868 59740 223874 59804
rect 223990 59742 234630 59802
rect 221181 59666 221247 59669
rect 223990 59666 224050 59742
rect 231025 59666 231091 59669
rect 221181 59664 224050 59666
rect 221181 59608 221186 59664
rect 221242 59608 224050 59664
rect 221181 59606 224050 59608
rect 224910 59664 231091 59666
rect 224910 59608 231030 59664
rect 231086 59608 231091 59664
rect 224910 59606 231091 59608
rect 221181 59603 221247 59606
rect 217593 59530 217659 59533
rect 224910 59530 224970 59606
rect 231025 59603 231091 59606
rect 217593 59528 224970 59530
rect 217593 59472 217598 59528
rect 217654 59472 224970 59528
rect 217593 59470 224970 59472
rect 217593 59467 217659 59470
rect 223021 59394 223087 59397
rect 230841 59394 230907 59397
rect 223021 59392 230907 59394
rect 223021 59336 223026 59392
rect 223082 59336 230846 59392
rect 230902 59336 230907 59392
rect 223021 59334 230907 59336
rect 234570 59394 234630 59742
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect 266353 59394 266419 59397
rect 234570 59392 266419 59394
rect 234570 59336 266358 59392
rect 266414 59336 266419 59392
rect 234570 59334 266419 59336
rect 223021 59331 223087 59334
rect 230841 59331 230907 59334
rect 266353 59331 266419 59334
rect 219985 59258 220051 59261
rect 224718 59258 224724 59260
rect 219985 59256 224724 59258
rect 219985 59200 219990 59256
rect 220046 59200 224724 59256
rect 219985 59198 224724 59200
rect 219985 59195 220051 59198
rect 224718 59196 224724 59198
rect 224788 59196 224794 59260
rect 212533 59122 212599 59125
rect 358813 59122 358879 59125
rect 212533 59120 358879 59122
rect 212533 59064 212538 59120
rect 212594 59064 358818 59120
rect 358874 59064 358879 59120
rect 212533 59062 358879 59064
rect 212533 59059 212599 59062
rect 358813 59059 358879 59062
rect 210141 58986 210207 58989
rect 357433 58986 357499 58989
rect 210141 58984 357499 58986
rect 210141 58928 210146 58984
rect 210202 58928 357438 58984
rect 357494 58928 357499 58984
rect 210141 58926 357499 58928
rect 210141 58923 210207 58926
rect 357433 58923 357499 58926
rect 219709 58850 219775 58853
rect 225045 58850 225111 58853
rect 219709 58848 225111 58850
rect 219709 58792 219714 58848
rect 219770 58792 225050 58848
rect 225106 58792 225111 58848
rect 219709 58790 225111 58792
rect 219709 58787 219775 58790
rect 225045 58787 225111 58790
rect -960 58578 480 58668
rect 3601 58578 3667 58581
rect -960 58576 3667 58578
rect -960 58520 3606 58576
rect 3662 58520 3667 58576
rect -960 58518 3667 58520
rect -960 58428 480 58518
rect 3601 58515 3667 58518
rect 58709 57898 58775 57901
rect 212809 57898 212875 57901
rect 58709 57896 212875 57898
rect 58709 57840 58714 57896
rect 58770 57840 212814 57896
rect 212870 57840 212875 57896
rect 58709 57838 212875 57840
rect 58709 57835 58775 57838
rect 212809 57835 212875 57838
rect 58617 57762 58683 57765
rect 62113 57762 62179 57765
rect 211061 57762 211127 57765
rect 58617 57760 62179 57762
rect 58617 57704 58622 57760
rect 58678 57704 62118 57760
rect 62174 57704 62179 57760
rect 58617 57702 62179 57704
rect 58617 57699 58683 57702
rect 62113 57699 62179 57702
rect 64830 57760 211127 57762
rect 64830 57704 211066 57760
rect 211122 57704 211127 57760
rect 64830 57702 211127 57704
rect 12341 57626 12407 57629
rect 62757 57626 62823 57629
rect 12341 57624 62823 57626
rect 12341 57568 12346 57624
rect 12402 57568 62762 57624
rect 62818 57568 62823 57624
rect 12341 57566 62823 57568
rect 12341 57563 12407 57566
rect 62757 57563 62823 57566
rect 10961 57490 11027 57493
rect 59997 57490 60063 57493
rect 63033 57490 63099 57493
rect 10961 57488 58818 57490
rect 10961 57432 10966 57488
rect 11022 57432 58818 57488
rect 10961 57430 58818 57432
rect 10961 57427 11027 57430
rect 9581 57354 9647 57357
rect 58617 57354 58683 57357
rect 9581 57352 58683 57354
rect 9581 57296 9586 57352
rect 9642 57296 58622 57352
rect 58678 57296 58683 57352
rect 9581 57294 58683 57296
rect 58758 57354 58818 57430
rect 59997 57488 63099 57490
rect 59997 57432 60002 57488
rect 60058 57432 63038 57488
rect 63094 57432 63099 57488
rect 59997 57430 63099 57432
rect 59997 57427 60063 57430
rect 63033 57427 63099 57430
rect 62481 57354 62547 57357
rect 58758 57352 62547 57354
rect 58758 57296 62486 57352
rect 62542 57296 62547 57352
rect 58758 57294 62547 57296
rect 9581 57291 9647 57294
rect 58617 57291 58683 57294
rect 62481 57291 62547 57294
rect 4061 57218 4127 57221
rect 60917 57218 60983 57221
rect 4061 57216 60983 57218
rect 4061 57160 4066 57216
rect 4122 57160 60922 57216
rect 60978 57160 60983 57216
rect 4061 57158 60983 57160
rect 4061 57155 4127 57158
rect 60917 57155 60983 57158
rect 15101 57082 15167 57085
rect 58525 57082 58591 57085
rect 64830 57082 64890 57702
rect 211061 57699 211127 57702
rect 215201 57762 215267 57765
rect 228081 57762 228147 57765
rect 215201 57760 228147 57762
rect 215201 57704 215206 57760
rect 215262 57704 228086 57760
rect 228142 57704 228147 57760
rect 215201 57702 228147 57704
rect 215201 57699 215267 57702
rect 228081 57699 228147 57702
rect 208025 57626 208091 57629
rect 228173 57626 228239 57629
rect 208025 57624 228239 57626
rect 208025 57568 208030 57624
rect 208086 57568 228178 57624
rect 228234 57568 228239 57624
rect 208025 57566 228239 57568
rect 208025 57563 208091 57566
rect 228173 57563 228239 57566
rect 214649 57490 214715 57493
rect 231209 57490 231275 57493
rect 214649 57488 231275 57490
rect 214649 57432 214654 57488
rect 214710 57432 231214 57488
rect 231270 57432 231275 57488
rect 214649 57430 231275 57432
rect 214649 57427 214715 57430
rect 231209 57427 231275 57430
rect 213729 57354 213795 57357
rect 224309 57354 224375 57357
rect 213729 57352 224375 57354
rect 213729 57296 213734 57352
rect 213790 57296 224314 57352
rect 224370 57296 224375 57352
rect 213729 57294 224375 57296
rect 213729 57291 213795 57294
rect 224309 57291 224375 57294
rect 180517 57218 180583 57221
rect 180793 57218 180859 57221
rect 180517 57216 180859 57218
rect 180517 57160 180522 57216
rect 180578 57160 180798 57216
rect 180854 57160 180859 57216
rect 180517 57158 180859 57160
rect 180517 57155 180583 57158
rect 180793 57155 180859 57158
rect 206921 57218 206987 57221
rect 436737 57218 436803 57221
rect 206921 57216 436803 57218
rect 206921 57160 206926 57216
rect 206982 57160 436742 57216
rect 436798 57160 436803 57216
rect 206921 57158 436803 57160
rect 206921 57155 206987 57158
rect 436737 57155 436803 57158
rect 15101 57080 58450 57082
rect 15101 57024 15106 57080
rect 15162 57024 58450 57080
rect 15101 57022 58450 57024
rect 15101 57019 15167 57022
rect 13721 56946 13787 56949
rect 58249 56946 58315 56949
rect 13721 56944 58315 56946
rect 13721 56888 13726 56944
rect 13782 56888 58254 56944
rect 58310 56888 58315 56944
rect 13721 56886 58315 56888
rect 58390 56946 58450 57022
rect 58525 57080 64890 57082
rect 58525 57024 58530 57080
rect 58586 57024 64890 57080
rect 58525 57022 64890 57024
rect 127801 57082 127867 57085
rect 132953 57082 133019 57085
rect 127801 57080 133019 57082
rect 127801 57024 127806 57080
rect 127862 57024 132958 57080
rect 133014 57024 133019 57080
rect 127801 57022 133019 57024
rect 58525 57019 58591 57022
rect 127801 57019 127867 57022
rect 132953 57019 133019 57022
rect 213177 57082 213243 57085
rect 255957 57082 256023 57085
rect 213177 57080 256023 57082
rect 213177 57024 213182 57080
rect 213238 57024 255962 57080
rect 256018 57024 256023 57080
rect 213177 57022 256023 57024
rect 213177 57019 213243 57022
rect 255957 57019 256023 57022
rect 63677 56946 63743 56949
rect 58390 56944 63743 56946
rect 58390 56888 63682 56944
rect 63738 56888 63743 56944
rect 58390 56886 63743 56888
rect 13721 56883 13787 56886
rect 58249 56883 58315 56886
rect 63677 56883 63743 56886
rect 211613 56946 211679 56949
rect 251817 56946 251883 56949
rect 211613 56944 251883 56946
rect 211613 56888 211618 56944
rect 211674 56888 251822 56944
rect 251878 56888 251883 56944
rect 211613 56886 251883 56888
rect 211613 56883 211679 56886
rect 251817 56883 251883 56886
rect 22001 56810 22067 56813
rect 65425 56810 65491 56813
rect 22001 56808 65491 56810
rect 22001 56752 22006 56808
rect 22062 56752 65430 56808
rect 65486 56752 65491 56808
rect 22001 56750 65491 56752
rect 22001 56747 22067 56750
rect 65425 56747 65491 56750
rect 211889 56810 211955 56813
rect 226241 56810 226307 56813
rect 211889 56808 226307 56810
rect 211889 56752 211894 56808
rect 211950 56752 226246 56808
rect 226302 56752 226307 56808
rect 211889 56750 226307 56752
rect 211889 56747 211955 56750
rect 226241 56747 226307 56750
rect 58249 56674 58315 56677
rect 63309 56674 63375 56677
rect 58249 56672 63375 56674
rect 58249 56616 58254 56672
rect 58310 56616 63314 56672
rect 63370 56616 63375 56672
rect 58249 56614 63375 56616
rect 58249 56611 58315 56614
rect 63309 56611 63375 56614
rect 217501 56674 217567 56677
rect 229461 56674 229527 56677
rect 217501 56672 229527 56674
rect 217501 56616 217506 56672
rect 217562 56616 229466 56672
rect 229522 56616 229527 56672
rect 217501 56614 229527 56616
rect 217501 56611 217567 56614
rect 229461 56611 229527 56614
rect 580257 46338 580323 46341
rect 583520 46338 584960 46428
rect 580257 46336 584960 46338
rect 580257 46280 580262 46336
rect 580318 46280 584960 46336
rect 580257 46278 584960 46280
rect 580257 46275 580323 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3325 45522 3391 45525
rect -960 45520 3391 45522
rect -960 45464 3330 45520
rect 3386 45464 3391 45520
rect -960 45462 3391 45464
rect -960 45372 480 45462
rect 3325 45459 3391 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2773 32466 2839 32469
rect -960 32464 2839 32466
rect -960 32408 2778 32464
rect 2834 32408 2839 32464
rect -960 32406 2839 32408
rect -960 32316 480 32406
rect 2773 32403 2839 32406
rect 580073 19818 580139 19821
rect 583520 19818 584960 19908
rect 580073 19816 584960 19818
rect 580073 19760 580078 19816
rect 580134 19760 584960 19816
rect 580073 19758 584960 19760
rect 580073 19755 580139 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3509 19410 3575 19413
rect -960 19408 3575 19410
rect -960 19352 3514 19408
rect 3570 19352 3575 19408
rect -960 19350 3575 19352
rect -960 19260 480 19350
rect 3509 19347 3575 19350
rect 208209 11794 208275 11797
rect 582189 11794 582255 11797
rect 208209 11792 582255 11794
rect 208209 11736 208214 11792
rect 208270 11736 582194 11792
rect 582250 11736 582255 11792
rect 208209 11734 582255 11736
rect 208209 11731 208275 11734
rect 582189 11731 582255 11734
rect 208301 11658 208367 11661
rect 583385 11658 583451 11661
rect 208301 11656 583451 11658
rect 208301 11600 208306 11656
rect 208362 11600 583390 11656
rect 583446 11600 583451 11656
rect 208301 11598 583451 11600
rect 208301 11595 208367 11598
rect 583385 11595 583451 11598
rect 181805 9482 181871 9485
rect 481725 9482 481791 9485
rect 181805 9480 481791 9482
rect 181805 9424 181810 9480
rect 181866 9424 481730 9480
rect 481786 9424 481791 9480
rect 181805 9422 481791 9424
rect 181805 9419 181871 9422
rect 481725 9419 481791 9422
rect 183369 9346 183435 9349
rect 485221 9346 485287 9349
rect 183369 9344 485287 9346
rect 183369 9288 183374 9344
rect 183430 9288 485226 9344
rect 485282 9288 485287 9344
rect 183369 9286 485287 9288
rect 183369 9283 183435 9286
rect 485221 9283 485287 9286
rect 184749 9210 184815 9213
rect 488809 9210 488875 9213
rect 184749 9208 488875 9210
rect 184749 9152 184754 9208
rect 184810 9152 488814 9208
rect 488870 9152 488875 9208
rect 184749 9150 488875 9152
rect 184749 9147 184815 9150
rect 488809 9147 488875 9150
rect 184565 9074 184631 9077
rect 492305 9074 492371 9077
rect 184565 9072 492371 9074
rect 184565 9016 184570 9072
rect 184626 9016 492310 9072
rect 492366 9016 492371 9072
rect 184565 9014 492371 9016
rect 184565 9011 184631 9014
rect 492305 9011 492371 9014
rect 187417 8938 187483 8941
rect 502977 8938 503043 8941
rect 187417 8936 503043 8938
rect 187417 8880 187422 8936
rect 187478 8880 502982 8936
rect 503038 8880 503043 8936
rect 187417 8878 503043 8880
rect 187417 8875 187483 8878
rect 502977 8875 503043 8878
rect 151629 6898 151695 6901
rect 358721 6898 358787 6901
rect 151629 6896 358787 6898
rect 151629 6840 151634 6896
rect 151690 6840 358726 6896
rect 358782 6840 358787 6896
rect 151629 6838 358787 6840
rect 151629 6835 151695 6838
rect 358721 6835 358787 6838
rect 151353 6762 151419 6765
rect 362309 6762 362375 6765
rect 151353 6760 362375 6762
rect 151353 6704 151358 6760
rect 151414 6704 362314 6760
rect 362370 6704 362375 6760
rect 151353 6702 362375 6704
rect 151353 6699 151419 6702
rect 362309 6699 362375 6702
rect 153101 6626 153167 6629
rect 365805 6626 365871 6629
rect 153101 6624 365871 6626
rect -960 6490 480 6580
rect 153101 6568 153106 6624
rect 153162 6568 365810 6624
rect 365866 6568 365871 6624
rect 153101 6566 365871 6568
rect 153101 6563 153167 6566
rect 365805 6563 365871 6566
rect 580349 6626 580415 6629
rect 583520 6626 584960 6716
rect 580349 6624 584960 6626
rect 580349 6568 580354 6624
rect 580410 6568 584960 6624
rect 580349 6566 584960 6568
rect 580349 6563 580415 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 157241 6490 157307 6493
rect 379973 6490 380039 6493
rect 157241 6488 380039 6490
rect 157241 6432 157246 6488
rect 157302 6432 379978 6488
rect 380034 6432 380039 6488
rect 583520 6476 584960 6566
rect 157241 6430 380039 6432
rect 157241 6427 157307 6430
rect 379973 6427 380039 6430
rect 157149 6354 157215 6357
rect 383561 6354 383627 6357
rect 157149 6352 383627 6354
rect 157149 6296 157154 6352
rect 157210 6296 383566 6352
rect 383622 6296 383627 6352
rect 157149 6294 383627 6296
rect 157149 6291 157215 6294
rect 383561 6291 383627 6294
rect 165153 6218 165219 6221
rect 411897 6218 411963 6221
rect 165153 6216 411963 6218
rect 165153 6160 165158 6216
rect 165214 6160 411902 6216
rect 411958 6160 411963 6216
rect 165153 6158 411963 6160
rect 165153 6155 165219 6158
rect 411897 6155 411963 6158
rect 219065 6082 219131 6085
rect 390645 6082 390711 6085
rect 219065 6080 390711 6082
rect 219065 6024 219070 6080
rect 219126 6024 390650 6080
rect 390706 6024 390711 6080
rect 219065 6022 390711 6024
rect 219065 6019 219131 6022
rect 390645 6019 390711 6022
rect 97901 4042 97967 4045
rect 149513 4042 149579 4045
rect 97901 4040 149579 4042
rect 97901 3984 97906 4040
rect 97962 3984 149518 4040
rect 149574 3984 149579 4040
rect 97901 3982 149579 3984
rect 97901 3979 97967 3982
rect 149513 3979 149579 3982
rect 170765 4042 170831 4045
rect 436737 4042 436803 4045
rect 170765 4040 436803 4042
rect 170765 3984 170770 4040
rect 170826 3984 436742 4040
rect 436798 3984 436803 4040
rect 170765 3982 436803 3984
rect 170765 3979 170831 3982
rect 436737 3979 436803 3982
rect 99189 3906 99255 3909
rect 153009 3906 153075 3909
rect 99189 3904 153075 3906
rect 99189 3848 99194 3904
rect 99250 3848 153014 3904
rect 153070 3848 153075 3904
rect 99189 3846 153075 3848
rect 99189 3843 99255 3846
rect 153009 3843 153075 3846
rect 176193 3906 176259 3909
rect 458081 3906 458147 3909
rect 176193 3904 458147 3906
rect 176193 3848 176198 3904
rect 176254 3848 458086 3904
rect 458142 3848 458147 3904
rect 176193 3846 458147 3848
rect 176193 3843 176259 3846
rect 458081 3843 458147 3846
rect 102041 3770 102107 3773
rect 161289 3770 161355 3773
rect 102041 3768 161355 3770
rect 102041 3712 102046 3768
rect 102102 3712 161294 3768
rect 161350 3712 161355 3768
rect 102041 3710 161355 3712
rect 102041 3707 102107 3710
rect 161289 3707 161355 3710
rect 180701 3770 180767 3773
rect 472249 3770 472315 3773
rect 180701 3768 472315 3770
rect 180701 3712 180706 3768
rect 180762 3712 472254 3768
rect 472310 3712 472315 3768
rect 180701 3710 472315 3712
rect 180701 3707 180767 3710
rect 472249 3707 472315 3710
rect 100569 3634 100635 3637
rect 160093 3634 160159 3637
rect 100569 3632 160159 3634
rect 100569 3576 100574 3632
rect 100630 3576 160098 3632
rect 160154 3576 160159 3632
rect 100569 3574 160159 3576
rect 100569 3571 100635 3574
rect 160093 3571 160159 3574
rect 181989 3634 182055 3637
rect 479333 3634 479399 3637
rect 181989 3632 479399 3634
rect 181989 3576 181994 3632
rect 182050 3576 479338 3632
rect 479394 3576 479399 3632
rect 181989 3574 479399 3576
rect 181989 3571 182055 3574
rect 479333 3571 479399 3574
rect 101949 3498 102015 3501
rect 164877 3498 164943 3501
rect 101949 3496 164943 3498
rect 101949 3440 101954 3496
rect 102010 3440 164882 3496
rect 164938 3440 164943 3496
rect 101949 3438 164943 3440
rect 101949 3435 102015 3438
rect 164877 3435 164943 3438
rect 182081 3498 182147 3501
rect 480529 3498 480595 3501
rect 182081 3496 480595 3498
rect 182081 3440 182086 3496
rect 182142 3440 480534 3496
rect 480590 3440 480595 3496
rect 182081 3438 480595 3440
rect 182081 3435 182147 3438
rect 480529 3435 480595 3438
rect 104801 3362 104867 3365
rect 175457 3362 175523 3365
rect 104801 3360 175523 3362
rect 104801 3304 104806 3360
rect 104862 3304 175462 3360
rect 175518 3304 175523 3360
rect 104801 3302 175523 3304
rect 104801 3299 104867 3302
rect 175457 3299 175523 3302
rect 183093 3362 183159 3365
rect 484025 3362 484091 3365
rect 183093 3360 484091 3362
rect 183093 3304 183098 3360
rect 183154 3304 484030 3360
rect 484086 3304 484091 3360
rect 183093 3302 484091 3304
rect 183093 3299 183159 3302
rect 484025 3299 484091 3302
rect 99281 3226 99347 3229
rect 150617 3226 150683 3229
rect 99281 3224 150683 3226
rect 99281 3168 99286 3224
rect 99342 3168 150622 3224
rect 150678 3168 150683 3224
rect 99281 3166 150683 3168
rect 99281 3163 99347 3166
rect 150617 3163 150683 3166
rect 169293 3226 169359 3229
rect 433241 3226 433307 3229
rect 169293 3224 433307 3226
rect 169293 3168 169298 3224
rect 169354 3168 433246 3224
rect 433302 3168 433307 3224
rect 169293 3166 433307 3168
rect 169293 3163 169359 3166
rect 433241 3163 433307 3166
<< via3 >>
rect 268516 487460 268580 487524
rect 150940 487188 151004 487252
rect 90956 487052 91020 487116
rect 141004 486916 141068 486980
rect 318380 486916 318444 486980
rect 145604 486780 145668 486844
rect 136036 486644 136100 486708
rect 256188 486644 256252 486708
rect 128676 486508 128740 486572
rect 131068 486508 131132 486572
rect 263548 486644 263612 486708
rect 260972 486508 261036 486572
rect 118556 486432 118620 486436
rect 118556 486376 118606 486432
rect 118606 486376 118620 486432
rect 118556 486372 118620 486376
rect 120764 486372 120828 486436
rect 273484 486508 273548 486572
rect 339724 486508 339788 486572
rect 323348 486372 323412 486436
rect 350764 486372 350828 486436
rect 101076 486236 101140 486300
rect 283788 486236 283852 486300
rect 288572 486296 288636 486300
rect 288572 486240 288586 486296
rect 288586 486240 288636 486296
rect 288572 486236 288636 486240
rect 98500 486100 98564 486164
rect 290964 486100 291028 486164
rect 295932 486160 295996 486164
rect 295932 486104 295946 486160
rect 295946 486104 295996 486160
rect 295932 486100 295996 486104
rect 93532 485964 93596 486028
rect 300716 485964 300780 486028
rect 111196 485828 111260 485892
rect 133644 485888 133708 485892
rect 133644 485832 133658 485888
rect 133658 485832 133708 485888
rect 133644 485828 133708 485832
rect 138612 485888 138676 485892
rect 138612 485832 138626 485888
rect 138626 485832 138676 485888
rect 138612 485828 138676 485832
rect 143580 485828 143644 485892
rect 154068 485828 154132 485892
rect 158484 485888 158548 485892
rect 158484 485832 158534 485888
rect 158534 485832 158548 485888
rect 158484 485828 158548 485832
rect 161060 485828 161124 485892
rect 251036 485828 251100 485892
rect 253428 485888 253492 485892
rect 253428 485832 253442 485888
rect 253442 485832 253492 485888
rect 253428 485828 253492 485832
rect 258396 485888 258460 485892
rect 258396 485832 258410 485888
rect 258410 485832 258460 485888
rect 258396 485828 258460 485832
rect 266124 485888 266188 485892
rect 266124 485832 266138 485888
rect 266138 485832 266188 485888
rect 266124 485828 266188 485832
rect 278452 485888 278516 485892
rect 278452 485832 278466 485888
rect 278466 485832 278516 485888
rect 278452 485828 278516 485832
rect 311020 485888 311084 485892
rect 311020 485832 311034 485888
rect 311034 485832 311084 485888
rect 311020 485828 311084 485832
rect 313596 485888 313660 485892
rect 313596 485832 313610 485888
rect 313610 485832 313660 485888
rect 313596 485828 313660 485832
rect 320956 485828 321020 485892
rect 126100 485556 126164 485620
rect 96292 485420 96356 485484
rect 156092 485284 156156 485348
rect 148364 485148 148428 485212
rect 285996 485148 286060 485212
rect 123708 485012 123772 485076
rect 276060 485012 276124 485076
rect 113588 484876 113652 484940
rect 293540 484876 293604 484940
rect 88748 484740 88812 484804
rect 103652 484740 103716 484804
rect 305868 484740 305932 484804
rect 271092 484604 271156 484668
rect 106044 484468 106108 484532
rect 190868 484468 190932 484532
rect 315804 484468 315868 484532
rect 338436 484468 338500 484532
rect 116164 484196 116228 484260
rect 179644 484060 179708 484124
rect 166028 483924 166092 483988
rect 178540 483924 178604 483988
rect 248644 483924 248708 483988
rect 303476 483788 303540 483852
rect 163366 483652 163430 483716
rect 308406 483652 308470 483716
rect 108558 483516 108622 483580
rect 326086 483516 326150 483580
rect 280934 483380 280998 483444
rect 298614 483380 298678 483444
rect 85436 398168 85500 398172
rect 85436 398112 85486 398168
rect 85486 398112 85500 398168
rect 85436 398108 85500 398112
rect 92428 398108 92492 398172
rect 95924 398168 95988 398172
rect 95924 398112 95938 398168
rect 95938 398112 95988 398168
rect 95924 398108 95988 398112
rect 113588 398168 113652 398172
rect 113588 398112 113638 398168
rect 113638 398112 113652 398168
rect 113588 398108 113652 398112
rect 223804 398108 223868 398172
rect 235948 398168 236012 398172
rect 235948 398112 235998 398168
rect 235998 398112 236012 398168
rect 235948 398108 236012 398112
rect 265204 398108 265268 398172
rect 300900 398108 300964 398172
rect 315804 398168 315868 398172
rect 315804 398112 315818 398168
rect 315818 398112 315868 398168
rect 315804 398108 315868 398112
rect 325924 398168 325988 398172
rect 325924 398112 325938 398168
rect 325938 398112 325988 398168
rect 325924 398108 325988 398112
rect 223620 397972 223684 398036
rect 224908 397836 224972 397900
rect 77156 397292 77220 397356
rect 78260 397352 78324 397356
rect 78260 397296 78310 397352
rect 78310 397296 78324 397352
rect 78260 397292 78324 397296
rect 79548 397352 79612 397356
rect 79548 397296 79598 397352
rect 79598 397296 79612 397352
rect 79548 397292 79612 397296
rect 80468 397352 80532 397356
rect 80468 397296 80482 397352
rect 80482 397296 80532 397352
rect 80468 397292 80532 397296
rect 81940 397292 82004 397356
rect 83044 397352 83108 397356
rect 83044 397296 83058 397352
rect 83058 397296 83108 397352
rect 83044 397292 83108 397296
rect 88748 397292 88812 397356
rect 90036 397352 90100 397356
rect 90036 397296 90086 397352
rect 90086 397296 90100 397352
rect 90036 397292 90100 397296
rect 91324 397292 91388 397356
rect 93348 397292 93412 397356
rect 94636 397292 94700 397356
rect 98132 397352 98196 397356
rect 98132 397296 98146 397352
rect 98146 397296 98196 397352
rect 98132 397292 98196 397296
rect 102732 397352 102796 397356
rect 102732 397296 102782 397352
rect 102782 397296 102796 397352
rect 102732 397292 102796 397296
rect 104020 397292 104084 397356
rect 105308 397292 105372 397356
rect 106412 397292 106476 397356
rect 108804 397352 108868 397356
rect 108804 397296 108854 397352
rect 108854 397296 108868 397352
rect 108804 397292 108868 397296
rect 109540 397292 109604 397356
rect 112300 397352 112364 397356
rect 112300 397296 112350 397352
rect 112350 397296 112364 397352
rect 112300 397292 112364 397296
rect 113220 397292 113284 397356
rect 114324 397292 114388 397356
rect 118188 397352 118252 397356
rect 118188 397296 118238 397352
rect 118238 397296 118252 397352
rect 118188 397292 118252 397296
rect 118556 397352 118620 397356
rect 118556 397296 118606 397352
rect 118606 397296 118620 397352
rect 118556 397292 118620 397296
rect 136036 397292 136100 397356
rect 154068 397352 154132 397356
rect 154068 397296 154118 397352
rect 154118 397296 154132 397352
rect 154068 397292 154132 397296
rect 163452 397292 163516 397356
rect 183508 397352 183572 397356
rect 183508 397296 183522 397352
rect 183522 397296 183572 397352
rect 183508 397292 183572 397296
rect 237052 397292 237116 397356
rect 239260 397352 239324 397356
rect 239260 397296 239274 397352
rect 239274 397296 239324 397352
rect 239260 397292 239324 397296
rect 247724 397352 247788 397356
rect 247724 397296 247738 397352
rect 247738 397296 247788 397352
rect 247724 397292 247788 397296
rect 248276 397292 248340 397356
rect 248644 397352 248708 397356
rect 248644 397296 248658 397352
rect 248658 397296 248708 397352
rect 248644 397292 248708 397296
rect 250116 397352 250180 397356
rect 250116 397296 250130 397352
rect 250130 397296 250180 397352
rect 250116 397292 250180 397296
rect 250668 397292 250732 397356
rect 253428 397292 253492 397356
rect 259500 397352 259564 397356
rect 259500 397296 259514 397352
rect 259514 397296 259564 397352
rect 259500 397292 259564 397296
rect 260972 397352 261036 397356
rect 260972 397296 260986 397352
rect 260986 397296 261036 397352
rect 260972 397292 261036 397296
rect 262076 397292 262140 397356
rect 262812 397292 262876 397356
rect 263916 397292 263980 397356
rect 268332 397352 268396 397356
rect 268332 397296 268346 397352
rect 268346 397296 268396 397352
rect 268332 397292 268396 397296
rect 268700 397352 268764 397356
rect 268700 397296 268714 397352
rect 268714 397296 268764 397352
rect 268700 397292 268764 397296
rect 272564 397292 272628 397356
rect 275324 397352 275388 397356
rect 275324 397296 275338 397352
rect 275338 397296 275388 397352
rect 275324 397292 275388 397296
rect 278084 397292 278148 397356
rect 279004 397292 279068 397356
rect 290964 397292 291028 397356
rect 298508 397352 298572 397356
rect 298508 397296 298522 397352
rect 298522 397296 298572 397352
rect 298508 397292 298572 397296
rect 308628 397352 308692 397356
rect 308628 397296 308642 397352
rect 308642 397296 308692 397352
rect 308628 397292 308692 397296
rect 343220 397292 343284 397356
rect 251220 397080 251284 397084
rect 251220 397024 251234 397080
rect 251234 397024 251284 397080
rect 251220 397020 251284 397024
rect 100708 396884 100772 396948
rect 258396 396884 258460 396948
rect 76052 396748 76116 396812
rect 84332 396748 84396 396812
rect 86540 396748 86604 396812
rect 87644 396748 87708 396812
rect 88380 396748 88444 396812
rect 90772 396748 90836 396812
rect 93716 396748 93780 396812
rect 96292 396748 96356 396812
rect 97028 396748 97092 396812
rect 98500 396748 98564 396812
rect 99972 396748 100036 396812
rect 101076 396748 101140 396812
rect 103836 396748 103900 396812
rect 106044 396808 106108 396812
rect 106044 396752 106058 396808
rect 106058 396752 106108 396808
rect 106044 396748 106108 396752
rect 107516 396808 107580 396812
rect 107516 396752 107530 396808
rect 107530 396752 107580 396808
rect 107516 396748 107580 396752
rect 111196 396748 111260 396812
rect 115796 396808 115860 396812
rect 115796 396752 115810 396808
rect 115810 396752 115860 396808
rect 115796 396748 115860 396752
rect 117084 396748 117148 396812
rect 119108 396748 119172 396812
rect 120764 396748 120828 396812
rect 123524 396748 123588 396812
rect 125916 396748 125980 396812
rect 128676 396748 128740 396812
rect 131068 396808 131132 396812
rect 131068 396752 131082 396808
rect 131082 396752 131132 396808
rect 131068 396748 131132 396752
rect 133460 396748 133524 396812
rect 138428 396748 138492 396812
rect 141004 396748 141068 396812
rect 143580 396748 143644 396812
rect 145604 396748 145668 396812
rect 148548 396748 148612 396812
rect 150940 396748 151004 396812
rect 155908 396808 155972 396812
rect 155908 396752 155958 396808
rect 155958 396752 155972 396808
rect 155908 396748 155972 396752
rect 158484 396748 158548 396812
rect 160876 396748 160940 396812
rect 166028 396748 166092 396812
rect 183140 396748 183204 396812
rect 238156 396748 238220 396812
rect 240548 396748 240612 396812
rect 241652 396748 241716 396812
rect 242940 396808 243004 396812
rect 242940 396752 242954 396808
rect 242954 396752 243004 396808
rect 242940 396748 243004 396752
rect 244228 396748 244292 396812
rect 245332 396748 245396 396812
rect 246436 396748 246500 396812
rect 252324 396748 252388 396812
rect 253612 396748 253676 396812
rect 254532 396748 254596 396812
rect 255820 396748 255884 396812
rect 256188 396808 256252 396812
rect 256188 396752 256202 396808
rect 256202 396752 256252 396808
rect 256188 396748 256252 396752
rect 256924 396808 256988 396812
rect 256924 396752 256938 396808
rect 256938 396752 256988 396808
rect 256924 396748 256988 396752
rect 258396 396748 258460 396812
rect 260604 396748 260668 396812
rect 263548 396748 263612 396812
rect 265940 396748 266004 396812
rect 266308 396808 266372 396812
rect 266308 396752 266358 396808
rect 266358 396752 266372 396808
rect 266308 396748 266372 396752
rect 269804 396748 269868 396812
rect 270908 396748 270972 396812
rect 273300 396808 273364 396812
rect 273300 396752 273350 396808
rect 273350 396752 273364 396808
rect 273300 396748 273364 396752
rect 274404 396748 274468 396812
rect 276244 396748 276308 396812
rect 278452 396748 278516 396812
rect 280844 396748 280908 396812
rect 283788 396808 283852 396812
rect 283788 396752 283802 396808
rect 283802 396752 283852 396808
rect 283788 396748 283852 396752
rect 285996 396808 286060 396812
rect 285996 396752 286010 396808
rect 286010 396752 286060 396808
rect 285996 396748 286060 396752
rect 288204 396748 288268 396812
rect 293356 396748 293420 396812
rect 295932 396748 295996 396812
rect 303476 396748 303540 396812
rect 305868 396748 305932 396812
rect 311020 396748 311084 396812
rect 313412 396748 313476 396812
rect 318380 396748 318444 396812
rect 320956 396748 321020 396812
rect 323348 396748 323412 396812
rect 343404 396748 343468 396812
rect 101812 396612 101876 396676
rect 108252 396612 108316 396676
rect 111012 396612 111076 396676
rect 115980 396672 116044 396676
rect 115980 396616 115994 396672
rect 115994 396616 116044 396672
rect 115980 396612 116044 396616
rect 267596 396612 267660 396676
rect 271276 396612 271340 396676
rect 273484 396672 273548 396676
rect 273484 396616 273498 396672
rect 273498 396616 273548 396672
rect 273484 396612 273548 396616
rect 276980 396612 277044 396676
rect 226380 322084 226444 322148
rect 226748 260068 226812 260132
rect 224908 234500 224972 234564
rect 226012 234500 226076 234564
rect 226564 232732 226628 232796
rect 226196 231508 226260 231572
rect 224724 230964 224788 231028
rect 226932 229876 226996 229940
rect 224172 228788 224236 228852
rect 224172 225796 224236 225860
rect 224908 224980 224972 225044
rect 225828 224980 225892 225044
rect 226380 115092 226444 115156
rect 226748 107748 226812 107812
rect 226932 80820 226996 80884
rect 226564 73476 226628 73540
rect 223068 60012 223132 60076
rect 223436 60012 223500 60076
rect 225092 60012 225156 60076
rect 223620 59876 223684 59940
rect 226012 59876 226076 59940
rect 223804 59740 223868 59804
rect 224724 59196 224788 59260
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 485308 60134 492618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 485308 63854 496338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 485308 67574 500058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 485308 74414 506898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 485308 78134 510618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 485308 81854 514338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 485308 85574 518058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 90955 487116 91021 487117
rect 90955 487052 90956 487116
rect 91020 487052 91021 487116
rect 90955 487051 91021 487052
rect 88747 484804 88813 484805
rect 88747 484740 88748 484804
rect 88812 484740 88813 484804
rect 88747 484739 88813 484740
rect 88750 483850 88810 484739
rect 88704 483790 88810 483850
rect 90958 483850 91018 487051
rect 91794 485308 92414 488898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 93531 486028 93597 486029
rect 93531 485964 93532 486028
rect 93596 485964 93597 486028
rect 93531 485963 93597 485964
rect 93534 483850 93594 485963
rect 95514 485308 96134 492618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 98499 486164 98565 486165
rect 98499 486100 98500 486164
rect 98564 486100 98565 486164
rect 98499 486099 98565 486100
rect 96291 485484 96357 485485
rect 96291 485420 96292 485484
rect 96356 485420 96357 485484
rect 96291 485419 96357 485420
rect 96294 483850 96354 485419
rect 98502 483850 98562 486099
rect 99234 485308 99854 496338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 101075 486300 101141 486301
rect 101075 486236 101076 486300
rect 101140 486236 101141 486300
rect 101075 486235 101141 486236
rect 90958 483790 91076 483850
rect 88704 483202 88764 483790
rect 91016 483202 91076 483790
rect 93464 483790 93594 483850
rect 96184 483790 96354 483850
rect 98496 483790 98562 483850
rect 101078 483850 101138 486235
rect 102954 485308 103574 500058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 109794 485308 110414 506898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 111195 485892 111261 485893
rect 111195 485828 111196 485892
rect 111260 485828 111261 485892
rect 111195 485827 111261 485828
rect 103651 484804 103717 484805
rect 103651 484740 103652 484804
rect 103716 484740 103717 484804
rect 103651 484739 103717 484740
rect 103654 483850 103714 484739
rect 106043 484532 106109 484533
rect 106043 484468 106044 484532
rect 106108 484468 106109 484532
rect 106043 484467 106109 484468
rect 101078 483790 101140 483850
rect 93464 483202 93524 483790
rect 96184 483202 96244 483790
rect 98496 483202 98556 483790
rect 101080 483202 101140 483790
rect 103528 483790 103714 483850
rect 106046 483850 106106 484467
rect 111198 483850 111258 485827
rect 113514 485308 114134 510618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 117234 485308 117854 514338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 118555 486436 118621 486437
rect 118555 486372 118556 486436
rect 118620 486372 118621 486436
rect 118555 486371 118621 486372
rect 120763 486436 120829 486437
rect 120763 486372 120764 486436
rect 120828 486372 120829 486436
rect 120763 486371 120829 486372
rect 113587 484940 113653 484941
rect 113587 484876 113588 484940
rect 113652 484876 113653 484940
rect 113587 484875 113653 484876
rect 106046 483790 106172 483850
rect 103528 483202 103588 483790
rect 106112 483202 106172 483790
rect 111144 483790 111258 483850
rect 113590 483850 113650 484875
rect 116163 484260 116229 484261
rect 116163 484196 116164 484260
rect 116228 484196 116229 484260
rect 116163 484195 116229 484196
rect 116166 483850 116226 484195
rect 118558 483850 118618 486371
rect 113590 483790 113652 483850
rect 116166 483790 116236 483850
rect 108557 483580 108623 483581
rect 108557 483516 108558 483580
rect 108622 483516 108623 483580
rect 108557 483515 108623 483516
rect 108560 483202 108620 483515
rect 111144 483202 111204 483790
rect 113592 483202 113652 483790
rect 116176 483202 116236 483790
rect 118488 483790 118618 483850
rect 120766 483850 120826 486371
rect 120954 485308 121574 518058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 126099 485620 126165 485621
rect 126099 485556 126100 485620
rect 126164 485556 126165 485620
rect 126099 485555 126165 485556
rect 123707 485076 123773 485077
rect 123707 485012 123708 485076
rect 123772 485012 123773 485076
rect 123707 485011 123773 485012
rect 123710 483850 123770 485011
rect 120766 483790 120996 483850
rect 118488 483202 118548 483790
rect 120936 483202 120996 483790
rect 123656 483790 123770 483850
rect 126102 483850 126162 485555
rect 127794 485308 128414 488898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 128675 486572 128741 486573
rect 128675 486508 128676 486572
rect 128740 486508 128741 486572
rect 128675 486507 128741 486508
rect 131067 486572 131133 486573
rect 131067 486508 131068 486572
rect 131132 486508 131133 486572
rect 131067 486507 131133 486508
rect 128678 483850 128738 486507
rect 131070 483850 131130 486507
rect 131514 485308 132134 492618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 133643 485892 133709 485893
rect 133643 485828 133644 485892
rect 133708 485828 133709 485892
rect 133643 485827 133709 485828
rect 133646 483850 133706 485827
rect 135234 485308 135854 496338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 136035 486708 136101 486709
rect 136035 486644 136036 486708
rect 136100 486644 136101 486708
rect 136035 486643 136101 486644
rect 136038 483850 136098 486643
rect 138611 485892 138677 485893
rect 138611 485828 138612 485892
rect 138676 485828 138677 485892
rect 138611 485827 138677 485828
rect 126102 483790 126164 483850
rect 123656 483202 123716 483790
rect 126104 483202 126164 483790
rect 128552 483790 128738 483850
rect 131000 483790 131130 483850
rect 133584 483790 133706 483850
rect 135896 483790 136098 483850
rect 138614 483850 138674 485827
rect 138954 485308 139574 500058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 141003 486980 141069 486981
rect 141003 486916 141004 486980
rect 141068 486916 141069 486980
rect 141003 486915 141069 486916
rect 141006 483850 141066 486915
rect 145603 486844 145669 486845
rect 145603 486780 145604 486844
rect 145668 486780 145669 486844
rect 145603 486779 145669 486780
rect 143579 485892 143645 485893
rect 143579 485828 143580 485892
rect 143644 485828 143645 485892
rect 143579 485827 143645 485828
rect 143582 483850 143642 485827
rect 138614 483790 138676 483850
rect 141006 483790 141124 483850
rect 128552 483202 128612 483790
rect 131000 483202 131060 483790
rect 133584 483202 133644 483790
rect 135896 483202 135956 483790
rect 138616 483202 138676 483790
rect 141064 483202 141124 483790
rect 143512 483790 143642 483850
rect 145606 483850 145666 486779
rect 145794 485308 146414 506898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 485308 150134 510618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 150939 487252 151005 487253
rect 150939 487188 150940 487252
rect 151004 487188 151005 487252
rect 150939 487187 151005 487188
rect 148363 485212 148429 485213
rect 148363 485148 148364 485212
rect 148428 485148 148429 485212
rect 148363 485147 148429 485148
rect 148366 483850 148426 485147
rect 150942 483850 151002 487187
rect 153234 485308 153854 514338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 154067 485892 154133 485893
rect 154067 485828 154068 485892
rect 154132 485828 154133 485892
rect 154067 485827 154133 485828
rect 154070 483850 154130 485827
rect 156091 485348 156157 485349
rect 156091 485284 156092 485348
rect 156156 485284 156157 485348
rect 156954 485308 157574 518058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 158483 485892 158549 485893
rect 158483 485828 158484 485892
rect 158548 485828 158549 485892
rect 158483 485827 158549 485828
rect 161059 485892 161125 485893
rect 161059 485828 161060 485892
rect 161124 485828 161125 485892
rect 161059 485827 161125 485828
rect 156091 485283 156157 485284
rect 156094 483850 156154 485283
rect 158486 483850 158546 485827
rect 161062 483850 161122 485827
rect 163794 485308 164414 488898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 167514 485308 168134 492618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 485308 171854 496338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 485308 175574 500058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 181794 485308 182414 506898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 485308 186134 510618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 485308 189854 514338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 485308 193574 518058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 190867 484532 190933 484533
rect 190867 484468 190868 484532
rect 190932 484468 190933 484532
rect 190867 484467 190933 484468
rect 179643 484124 179709 484125
rect 179643 484060 179644 484124
rect 179708 484060 179709 484124
rect 179643 484059 179709 484060
rect 166027 483988 166093 483989
rect 166027 483924 166028 483988
rect 166092 483924 166093 483988
rect 166027 483923 166093 483924
rect 178539 483988 178605 483989
rect 178539 483924 178540 483988
rect 178604 483924 178605 483988
rect 178539 483923 178605 483924
rect 145606 483790 146020 483850
rect 148366 483790 148468 483850
rect 150942 483790 151052 483850
rect 143512 483202 143572 483790
rect 145960 483202 146020 483790
rect 148408 483202 148468 483790
rect 150992 483202 151052 483790
rect 153576 483790 154130 483850
rect 156024 483790 156154 483850
rect 158472 483790 158546 483850
rect 161056 483790 161122 483850
rect 166030 483850 166090 483923
rect 178542 483850 178602 483923
rect 166030 483790 166148 483850
rect 153576 483202 153636 483790
rect 156024 483202 156084 483790
rect 158472 483202 158532 483790
rect 161056 483202 161116 483790
rect 163365 483716 163431 483717
rect 163365 483652 163366 483716
rect 163430 483652 163431 483716
rect 163365 483651 163431 483652
rect 163368 483202 163428 483651
rect 166088 483202 166148 483790
rect 178464 483790 178602 483850
rect 179646 483850 179706 484059
rect 190870 483850 190930 484467
rect 179646 483790 179748 483850
rect 178464 483202 178524 483790
rect 179688 483202 179748 483790
rect 190840 483790 190930 483850
rect 190840 483202 190900 483790
rect 60952 471454 61300 471486
rect 60952 471218 61008 471454
rect 61244 471218 61300 471454
rect 60952 471134 61300 471218
rect 60952 470898 61008 471134
rect 61244 470898 61300 471134
rect 60952 470866 61300 470898
rect 195320 471454 195668 471486
rect 195320 471218 195376 471454
rect 195612 471218 195668 471454
rect 195320 471134 195668 471218
rect 195320 470898 195376 471134
rect 195612 470898 195668 471134
rect 195320 470866 195668 470898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 60272 453454 60620 453486
rect 60272 453218 60328 453454
rect 60564 453218 60620 453454
rect 60272 453134 60620 453218
rect 60272 452898 60328 453134
rect 60564 452898 60620 453134
rect 60272 452866 60620 452898
rect 196000 453454 196348 453486
rect 196000 453218 196056 453454
rect 196292 453218 196348 453454
rect 196000 453134 196348 453218
rect 196000 452898 196056 453134
rect 196292 452898 196348 453134
rect 196000 452866 196348 452898
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 60952 435454 61300 435486
rect 60952 435218 61008 435454
rect 61244 435218 61300 435454
rect 60952 435134 61300 435218
rect 60952 434898 61008 435134
rect 61244 434898 61300 435134
rect 60952 434866 61300 434898
rect 195320 435454 195668 435486
rect 195320 435218 195376 435454
rect 195612 435218 195668 435454
rect 195320 435134 195668 435218
rect 195320 434898 195376 435134
rect 195612 434898 195668 435134
rect 195320 434866 195668 434898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 60272 417454 60620 417486
rect 60272 417218 60328 417454
rect 60564 417218 60620 417454
rect 60272 417134 60620 417218
rect 60272 416898 60328 417134
rect 60564 416898 60620 417134
rect 60272 416866 60620 416898
rect 196000 417454 196348 417486
rect 196000 417218 196056 417454
rect 196292 417218 196348 417454
rect 196000 417134 196348 417218
rect 196000 416898 196056 417134
rect 196292 416898 196348 417134
rect 196000 416866 196348 416898
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 76056 399530 76116 400106
rect 76054 399470 76116 399530
rect 77144 399530 77204 400106
rect 78232 399530 78292 400106
rect 79592 399530 79652 400106
rect 80544 399530 80604 400106
rect 77144 399470 77218 399530
rect 78232 399470 78322 399530
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 59514 385174 60134 398000
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 228924 60134 240618
rect 63234 388894 63854 398000
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 228924 63854 244338
rect 66954 392614 67574 398000
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 228924 67574 248058
rect 73794 363454 74414 398000
rect 76054 396813 76114 399470
rect 77158 397357 77218 399470
rect 77155 397356 77221 397357
rect 77155 397292 77156 397356
rect 77220 397292 77221 397356
rect 77155 397291 77221 397292
rect 76051 396812 76117 396813
rect 76051 396748 76052 396812
rect 76116 396748 76117 396812
rect 76051 396747 76117 396748
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 228924 74414 254898
rect 77514 367174 78134 398000
rect 78262 397357 78322 399470
rect 79550 399470 79652 399530
rect 80470 399470 80604 399530
rect 81768 399530 81828 400106
rect 83128 399530 83188 400106
rect 81768 399470 82002 399530
rect 79550 397357 79610 399470
rect 80470 397357 80530 399470
rect 78259 397356 78325 397357
rect 78259 397292 78260 397356
rect 78324 397292 78325 397356
rect 78259 397291 78325 397292
rect 79547 397356 79613 397357
rect 79547 397292 79548 397356
rect 79612 397292 79613 397356
rect 79547 397291 79613 397292
rect 80467 397356 80533 397357
rect 80467 397292 80468 397356
rect 80532 397292 80533 397356
rect 80467 397291 80533 397292
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 228924 78134 258618
rect 81234 370894 81854 398000
rect 81942 397357 82002 399470
rect 83046 399470 83188 399530
rect 84216 399530 84276 400106
rect 85440 399530 85500 400106
rect 84216 399470 84394 399530
rect 83046 397357 83106 399470
rect 81939 397356 82005 397357
rect 81939 397292 81940 397356
rect 82004 397292 82005 397356
rect 81939 397291 82005 397292
rect 83043 397356 83109 397357
rect 83043 397292 83044 397356
rect 83108 397292 83109 397356
rect 83043 397291 83109 397292
rect 84334 396813 84394 399470
rect 85438 399470 85500 399530
rect 86528 399530 86588 400106
rect 87616 399530 87676 400106
rect 88296 399530 88356 400106
rect 88704 399530 88764 400106
rect 90064 399530 90124 400106
rect 86528 399470 86602 399530
rect 87616 399470 87706 399530
rect 88296 399470 88442 399530
rect 88704 399470 88810 399530
rect 85438 398173 85498 399470
rect 85435 398172 85501 398173
rect 85435 398108 85436 398172
rect 85500 398108 85501 398172
rect 85435 398107 85501 398108
rect 84331 396812 84397 396813
rect 84331 396748 84332 396812
rect 84396 396748 84397 396812
rect 84331 396747 84397 396748
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 228924 81854 262338
rect 84954 374614 85574 398000
rect 86542 396813 86602 399470
rect 87646 396813 87706 399470
rect 88382 396813 88442 399470
rect 88750 397357 88810 399470
rect 90038 399470 90124 399530
rect 90744 399530 90804 400106
rect 91288 399530 91348 400106
rect 92376 399530 92436 400106
rect 93464 399530 93524 400106
rect 90744 399470 90834 399530
rect 91288 399470 91386 399530
rect 92376 399470 92490 399530
rect 90038 397357 90098 399470
rect 88747 397356 88813 397357
rect 88747 397292 88748 397356
rect 88812 397292 88813 397356
rect 88747 397291 88813 397292
rect 90035 397356 90101 397357
rect 90035 397292 90036 397356
rect 90100 397292 90101 397356
rect 90035 397291 90101 397292
rect 90774 396813 90834 399470
rect 91326 397357 91386 399470
rect 92430 398173 92490 399470
rect 93350 399470 93524 399530
rect 93600 399530 93660 400106
rect 94552 399530 94612 400106
rect 95912 399530 95972 400106
rect 96048 399530 96108 400106
rect 97000 399530 97060 400106
rect 98088 399530 98148 400106
rect 98496 399530 98556 400106
rect 99448 399530 99508 400106
rect 100672 399530 100732 400106
rect 101080 399530 101140 400106
rect 93600 399470 93778 399530
rect 94552 399470 94698 399530
rect 95912 399470 95986 399530
rect 96048 399470 96354 399530
rect 97000 399470 97090 399530
rect 98088 399470 98194 399530
rect 98496 399470 98562 399530
rect 99448 399470 100034 399530
rect 100672 399470 100770 399530
rect 92427 398172 92493 398173
rect 92427 398108 92428 398172
rect 92492 398108 92493 398172
rect 92427 398107 92493 398108
rect 91323 397356 91389 397357
rect 91323 397292 91324 397356
rect 91388 397292 91389 397356
rect 91323 397291 91389 397292
rect 86539 396812 86605 396813
rect 86539 396748 86540 396812
rect 86604 396748 86605 396812
rect 86539 396747 86605 396748
rect 87643 396812 87709 396813
rect 87643 396748 87644 396812
rect 87708 396748 87709 396812
rect 87643 396747 87709 396748
rect 88379 396812 88445 396813
rect 88379 396748 88380 396812
rect 88444 396748 88445 396812
rect 88379 396747 88445 396748
rect 90771 396812 90837 396813
rect 90771 396748 90772 396812
rect 90836 396748 90837 396812
rect 90771 396747 90837 396748
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 228924 85574 230058
rect 91794 381454 92414 398000
rect 93350 397357 93410 399470
rect 93347 397356 93413 397357
rect 93347 397292 93348 397356
rect 93412 397292 93413 397356
rect 93347 397291 93413 397292
rect 93718 396813 93778 399470
rect 94638 397357 94698 399470
rect 95926 398173 95986 399470
rect 95923 398172 95989 398173
rect 95923 398108 95924 398172
rect 95988 398108 95989 398172
rect 95923 398107 95989 398108
rect 94635 397356 94701 397357
rect 94635 397292 94636 397356
rect 94700 397292 94701 397356
rect 94635 397291 94701 397292
rect 93715 396812 93781 396813
rect 93715 396748 93716 396812
rect 93780 396748 93781 396812
rect 93715 396747 93781 396748
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 228924 92414 236898
rect 95514 385174 96134 398000
rect 96294 396813 96354 399470
rect 97030 396813 97090 399470
rect 98134 397357 98194 399470
rect 98131 397356 98197 397357
rect 98131 397292 98132 397356
rect 98196 397292 98197 397356
rect 98131 397291 98197 397292
rect 98502 396813 98562 399470
rect 96291 396812 96357 396813
rect 96291 396748 96292 396812
rect 96356 396748 96357 396812
rect 96291 396747 96357 396748
rect 97027 396812 97093 396813
rect 97027 396748 97028 396812
rect 97092 396748 97093 396812
rect 97027 396747 97093 396748
rect 98499 396812 98565 396813
rect 98499 396748 98500 396812
rect 98564 396748 98565 396812
rect 98499 396747 98565 396748
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 228924 96134 240618
rect 99234 388894 99854 398000
rect 99974 396813 100034 399470
rect 100710 396949 100770 399470
rect 101078 399470 101140 399530
rect 101760 399530 101820 400106
rect 102848 399530 102908 400106
rect 101760 399470 101874 399530
rect 100707 396948 100773 396949
rect 100707 396884 100708 396948
rect 100772 396884 100773 396948
rect 100707 396883 100773 396884
rect 101078 396813 101138 399470
rect 99971 396812 100037 396813
rect 99971 396748 99972 396812
rect 100036 396748 100037 396812
rect 99971 396747 100037 396748
rect 101075 396812 101141 396813
rect 101075 396748 101076 396812
rect 101140 396748 101141 396812
rect 101075 396747 101141 396748
rect 101814 396677 101874 399470
rect 102734 399470 102908 399530
rect 103528 399530 103588 400106
rect 103936 399530 103996 400106
rect 105296 399530 105356 400106
rect 105976 399530 106036 400106
rect 106384 399530 106444 400106
rect 107608 399530 107668 400106
rect 108288 399530 108348 400106
rect 103528 399470 103714 399530
rect 103936 399470 104082 399530
rect 105296 399470 105370 399530
rect 105976 399470 106106 399530
rect 106384 399470 106474 399530
rect 102734 397357 102794 399470
rect 102731 397356 102797 397357
rect 102731 397292 102732 397356
rect 102796 397292 102797 397356
rect 102731 397291 102797 397292
rect 101811 396676 101877 396677
rect 101811 396612 101812 396676
rect 101876 396612 101877 396676
rect 101811 396611 101877 396612
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 228924 99854 244338
rect 102954 392614 103574 398000
rect 103654 396810 103714 399470
rect 104022 397357 104082 399470
rect 105310 397357 105370 399470
rect 104019 397356 104085 397357
rect 104019 397292 104020 397356
rect 104084 397292 104085 397356
rect 104019 397291 104085 397292
rect 105307 397356 105373 397357
rect 105307 397292 105308 397356
rect 105372 397292 105373 397356
rect 105307 397291 105373 397292
rect 106046 396813 106106 399470
rect 106414 397357 106474 399470
rect 107518 399470 107668 399530
rect 108254 399470 108348 399530
rect 108696 399530 108756 400106
rect 109784 399530 109844 400106
rect 108696 399470 108866 399530
rect 106411 397356 106477 397357
rect 106411 397292 106412 397356
rect 106476 397292 106477 397356
rect 106411 397291 106477 397292
rect 107518 396813 107578 399470
rect 103835 396812 103901 396813
rect 103835 396810 103836 396812
rect 103654 396750 103836 396810
rect 103835 396748 103836 396750
rect 103900 396748 103901 396812
rect 103835 396747 103901 396748
rect 106043 396812 106109 396813
rect 106043 396748 106044 396812
rect 106108 396748 106109 396812
rect 106043 396747 106109 396748
rect 107515 396812 107581 396813
rect 107515 396748 107516 396812
rect 107580 396748 107581 396812
rect 107515 396747 107581 396748
rect 108254 396677 108314 399470
rect 108806 397357 108866 399470
rect 109542 399470 109844 399530
rect 111008 399530 111068 400106
rect 111144 399530 111204 400106
rect 112232 399530 112292 400106
rect 113320 399530 113380 400106
rect 111008 399470 111074 399530
rect 111144 399470 111258 399530
rect 112232 399470 112362 399530
rect 109542 397357 109602 399470
rect 108803 397356 108869 397357
rect 108803 397292 108804 397356
rect 108868 397292 108869 397356
rect 108803 397291 108869 397292
rect 109539 397356 109605 397357
rect 109539 397292 109540 397356
rect 109604 397292 109605 397356
rect 109539 397291 109605 397292
rect 108251 396676 108317 396677
rect 108251 396612 108252 396676
rect 108316 396612 108317 396676
rect 108251 396611 108317 396612
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 228924 103574 248058
rect 109794 363454 110414 398000
rect 111014 396677 111074 399470
rect 111198 396813 111258 399470
rect 112302 397357 112362 399470
rect 113222 399470 113380 399530
rect 113222 397357 113282 399470
rect 113590 398173 113650 400136
rect 114408 399530 114468 400106
rect 114326 399470 114468 399530
rect 113587 398172 113653 398173
rect 113587 398108 113588 398172
rect 113652 398108 113653 398172
rect 113587 398107 113653 398108
rect 112299 397356 112365 397357
rect 112299 397292 112300 397356
rect 112364 397292 112365 397356
rect 112299 397291 112365 397292
rect 113219 397356 113285 397357
rect 113219 397292 113220 397356
rect 113284 397292 113285 397356
rect 113219 397291 113285 397292
rect 111195 396812 111261 396813
rect 111195 396748 111196 396812
rect 111260 396748 111261 396812
rect 111195 396747 111261 396748
rect 111011 396676 111077 396677
rect 111011 396612 111012 396676
rect 111076 396612 111077 396676
rect 111011 396611 111077 396612
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 228924 110414 254898
rect 113514 367174 114134 398000
rect 114326 397357 114386 399470
rect 114323 397356 114389 397357
rect 114323 397292 114324 397356
rect 114388 397292 114389 397356
rect 114323 397291 114389 397292
rect 115798 396813 115858 400136
rect 115982 400076 116070 400136
rect 115795 396812 115861 396813
rect 115795 396748 115796 396812
rect 115860 396748 115861 396812
rect 115795 396747 115861 396748
rect 115982 396677 116042 400076
rect 116992 399530 117052 400106
rect 118080 399530 118140 400106
rect 118488 399530 118548 400106
rect 119168 399530 119228 400106
rect 120936 399530 120996 400106
rect 116992 399470 117146 399530
rect 118080 399470 118250 399530
rect 118488 399470 118618 399530
rect 117086 396813 117146 399470
rect 117083 396812 117149 396813
rect 117083 396748 117084 396812
rect 117148 396748 117149 396812
rect 117083 396747 117149 396748
rect 115979 396676 116045 396677
rect 115979 396612 115980 396676
rect 116044 396612 116045 396676
rect 115979 396611 116045 396612
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 228924 114134 258618
rect 117234 370894 117854 398000
rect 118190 397357 118250 399470
rect 118558 397357 118618 399470
rect 119110 399470 119228 399530
rect 120766 399470 120996 399530
rect 123520 399530 123580 400106
rect 125968 399530 126028 400106
rect 123520 399470 123586 399530
rect 118187 397356 118253 397357
rect 118187 397292 118188 397356
rect 118252 397292 118253 397356
rect 118187 397291 118253 397292
rect 118555 397356 118621 397357
rect 118555 397292 118556 397356
rect 118620 397292 118621 397356
rect 118555 397291 118621 397292
rect 119110 396813 119170 399470
rect 120766 396813 120826 399470
rect 119107 396812 119173 396813
rect 119107 396748 119108 396812
rect 119172 396748 119173 396812
rect 119107 396747 119173 396748
rect 120763 396812 120829 396813
rect 120763 396748 120764 396812
rect 120828 396748 120829 396812
rect 120763 396747 120829 396748
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 228924 117854 262338
rect 120954 374614 121574 398000
rect 123526 396813 123586 399470
rect 125918 399470 126028 399530
rect 128280 399530 128340 400106
rect 131000 399530 131060 400106
rect 133448 399530 133508 400106
rect 135896 399530 135956 400106
rect 138480 399530 138540 400106
rect 128280 399470 128554 399530
rect 131000 399470 131130 399530
rect 133448 399470 133522 399530
rect 135896 399470 136098 399530
rect 125918 396813 125978 399470
rect 123523 396812 123589 396813
rect 123523 396748 123524 396812
rect 123588 396748 123589 396812
rect 123523 396747 123589 396748
rect 125915 396812 125981 396813
rect 125915 396748 125916 396812
rect 125980 396748 125981 396812
rect 125915 396747 125981 396748
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 228924 121574 230058
rect 127794 381454 128414 398000
rect 128494 396810 128554 399470
rect 131070 396813 131130 399470
rect 128675 396812 128741 396813
rect 128675 396810 128676 396812
rect 128494 396750 128676 396810
rect 128675 396748 128676 396750
rect 128740 396748 128741 396812
rect 128675 396747 128741 396748
rect 131067 396812 131133 396813
rect 131067 396748 131068 396812
rect 131132 396748 131133 396812
rect 131067 396747 131133 396748
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 228924 128414 236898
rect 131514 385174 132134 398000
rect 133462 396813 133522 399470
rect 133459 396812 133525 396813
rect 133459 396748 133460 396812
rect 133524 396748 133525 396812
rect 133459 396747 133525 396748
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 228924 132134 240618
rect 135234 388894 135854 398000
rect 136038 397357 136098 399470
rect 138430 399470 138540 399530
rect 140928 399530 140988 400106
rect 143512 399530 143572 400106
rect 145960 399530 146020 400106
rect 140928 399470 141066 399530
rect 143512 399470 143642 399530
rect 136035 397356 136101 397357
rect 136035 397292 136036 397356
rect 136100 397292 136101 397356
rect 136035 397291 136101 397292
rect 138430 396813 138490 399470
rect 138427 396812 138493 396813
rect 138427 396748 138428 396812
rect 138492 396748 138493 396812
rect 138427 396747 138493 396748
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 228924 135854 244338
rect 138954 392614 139574 398000
rect 141006 396813 141066 399470
rect 143582 396813 143642 399470
rect 145606 399470 146020 399530
rect 148544 399530 148604 400106
rect 150992 399530 151052 400106
rect 148544 399470 148610 399530
rect 145606 396813 145666 399470
rect 141003 396812 141069 396813
rect 141003 396748 141004 396812
rect 141068 396748 141069 396812
rect 141003 396747 141069 396748
rect 143579 396812 143645 396813
rect 143579 396748 143580 396812
rect 143644 396748 143645 396812
rect 143579 396747 143645 396748
rect 145603 396812 145669 396813
rect 145603 396748 145604 396812
rect 145668 396748 145669 396812
rect 145603 396747 145669 396748
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 228924 139574 248058
rect 145794 363454 146414 398000
rect 148550 396813 148610 399470
rect 150942 399470 151052 399530
rect 153440 399530 153500 400106
rect 155888 399530 155948 400106
rect 158472 399530 158532 400106
rect 160920 399530 160980 400106
rect 153440 399470 154130 399530
rect 155888 399470 155970 399530
rect 158472 399470 158546 399530
rect 148547 396812 148613 396813
rect 148547 396748 148548 396812
rect 148612 396748 148613 396812
rect 148547 396747 148613 396748
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 228924 146414 254898
rect 149514 367174 150134 398000
rect 150942 396813 151002 399470
rect 150939 396812 151005 396813
rect 150939 396748 150940 396812
rect 151004 396748 151005 396812
rect 150939 396747 151005 396748
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 228924 150134 258618
rect 153234 370894 153854 398000
rect 154070 397357 154130 399470
rect 154067 397356 154133 397357
rect 154067 397292 154068 397356
rect 154132 397292 154133 397356
rect 154067 397291 154133 397292
rect 155910 396813 155970 399470
rect 155907 396812 155973 396813
rect 155907 396748 155908 396812
rect 155972 396748 155973 396812
rect 155907 396747 155973 396748
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 228924 153854 262338
rect 156954 374614 157574 398000
rect 158486 396813 158546 399470
rect 160878 399470 160980 399530
rect 163368 399530 163428 400106
rect 165952 399530 166012 400106
rect 183224 399530 183284 400106
rect 163368 399470 163514 399530
rect 165952 399470 166090 399530
rect 160878 396813 160938 399470
rect 163454 397357 163514 399470
rect 163451 397356 163517 397357
rect 163451 397292 163452 397356
rect 163516 397292 163517 397356
rect 163451 397291 163517 397292
rect 158483 396812 158549 396813
rect 158483 396748 158484 396812
rect 158548 396748 158549 396812
rect 158483 396747 158549 396748
rect 160875 396812 160941 396813
rect 160875 396748 160876 396812
rect 160940 396748 160941 396812
rect 160875 396747 160941 396748
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 228924 157574 230058
rect 163794 381454 164414 398000
rect 166030 396813 166090 399470
rect 183142 399470 183284 399530
rect 183360 399530 183420 400106
rect 183360 399470 183570 399530
rect 166027 396812 166093 396813
rect 166027 396748 166028 396812
rect 166092 396748 166093 396812
rect 166027 396747 166093 396748
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 228924 164414 236898
rect 167514 385174 168134 398000
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 228924 168134 240618
rect 171234 388894 171854 398000
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 228924 171854 244338
rect 174954 392614 175574 398000
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 228924 175574 248058
rect 181794 363454 182414 398000
rect 183142 396813 183202 399470
rect 183510 397357 183570 399470
rect 183507 397356 183573 397357
rect 183507 397292 183508 397356
rect 183572 397292 183573 397356
rect 183507 397291 183573 397292
rect 183139 396812 183205 396813
rect 183139 396748 183140 396812
rect 183204 396748 183205 396812
rect 183139 396747 183205 396748
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 228924 182414 254898
rect 185514 367174 186134 398000
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 228924 186134 258618
rect 189234 370894 189854 398000
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 228924 189854 262338
rect 192954 374614 193574 398000
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 228924 193574 230058
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 228924 200414 236898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 228924 204134 240618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 228924 207854 244338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217794 485308 218414 506898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 221514 485308 222134 510618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 485308 225854 514338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 485308 229574 518058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 485308 236414 488898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 485308 240134 492618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 485308 243854 496338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 485308 247574 500058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 251035 485892 251101 485893
rect 251035 485828 251036 485892
rect 251100 485828 251101 485892
rect 251035 485827 251101 485828
rect 253427 485892 253493 485893
rect 253427 485828 253428 485892
rect 253492 485828 253493 485892
rect 253427 485827 253493 485828
rect 248643 483988 248709 483989
rect 248643 483924 248644 483988
rect 248708 483924 248709 483988
rect 248643 483923 248709 483924
rect 248646 483850 248706 483923
rect 251038 483850 251098 485827
rect 248646 483790 248764 483850
rect 248704 483202 248764 483790
rect 251016 483790 251098 483850
rect 253430 483850 253490 485827
rect 253794 485308 254414 506898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 256187 486708 256253 486709
rect 256187 486644 256188 486708
rect 256252 486644 256253 486708
rect 256187 486643 256253 486644
rect 256190 483850 256250 486643
rect 257514 485308 258134 510618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 260971 486572 261037 486573
rect 260971 486508 260972 486572
rect 261036 486508 261037 486572
rect 260971 486507 261037 486508
rect 258395 485892 258461 485893
rect 258395 485828 258396 485892
rect 258460 485828 258461 485892
rect 258395 485827 258461 485828
rect 253430 483790 253524 483850
rect 251016 483202 251076 483790
rect 253464 483202 253524 483790
rect 256184 483790 256250 483850
rect 258398 483850 258458 485827
rect 260974 483850 261034 486507
rect 261234 485308 261854 514338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 263547 486708 263613 486709
rect 263547 486644 263548 486708
rect 263612 486644 263613 486708
rect 263547 486643 263613 486644
rect 263550 483850 263610 486643
rect 264954 485308 265574 518058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 268515 487524 268581 487525
rect 268515 487460 268516 487524
rect 268580 487460 268581 487524
rect 268515 487459 268581 487460
rect 266123 485892 266189 485893
rect 266123 485828 266124 485892
rect 266188 485828 266189 485892
rect 266123 485827 266189 485828
rect 266126 483850 266186 485827
rect 258398 483790 258556 483850
rect 260974 483790 261140 483850
rect 256184 483202 256244 483790
rect 258496 483202 258556 483790
rect 261080 483202 261140 483790
rect 263528 483790 263610 483850
rect 266112 483790 266186 483850
rect 268518 483850 268578 487459
rect 271794 485308 272414 488898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 273483 486572 273549 486573
rect 273483 486508 273484 486572
rect 273548 486508 273549 486572
rect 273483 486507 273549 486508
rect 271091 484668 271157 484669
rect 271091 484604 271092 484668
rect 271156 484604 271157 484668
rect 271091 484603 271157 484604
rect 271094 483850 271154 484603
rect 273486 483850 273546 486507
rect 275514 485308 276134 492618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 278451 485892 278517 485893
rect 278451 485828 278452 485892
rect 278516 485828 278517 485892
rect 278451 485827 278517 485828
rect 276059 485076 276125 485077
rect 276059 485012 276060 485076
rect 276124 485012 276125 485076
rect 276059 485011 276125 485012
rect 276062 483850 276122 485011
rect 278454 483850 278514 485827
rect 279234 485308 279854 496338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 485308 283574 500058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 283787 486300 283853 486301
rect 283787 486236 283788 486300
rect 283852 486236 283853 486300
rect 283787 486235 283853 486236
rect 288571 486300 288637 486301
rect 288571 486236 288572 486300
rect 288636 486236 288637 486300
rect 288571 486235 288637 486236
rect 283790 483850 283850 486235
rect 285995 485212 286061 485213
rect 285995 485148 285996 485212
rect 286060 485148 286061 485212
rect 285995 485147 286061 485148
rect 268518 483790 268620 483850
rect 271094 483790 271204 483850
rect 273486 483790 273652 483850
rect 276062 483790 276236 483850
rect 278454 483790 278548 483850
rect 263528 483202 263588 483790
rect 266112 483202 266172 483790
rect 268560 483202 268620 483790
rect 271144 483202 271204 483790
rect 273592 483202 273652 483790
rect 276176 483202 276236 483790
rect 278488 483202 278548 483790
rect 283656 483790 283850 483850
rect 285998 483850 286058 485147
rect 288574 483850 288634 486235
rect 289794 485308 290414 506898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 290963 486164 291029 486165
rect 290963 486100 290964 486164
rect 291028 486100 291029 486164
rect 290963 486099 291029 486100
rect 285998 483790 286164 483850
rect 280933 483444 280999 483445
rect 280933 483380 280934 483444
rect 280998 483380 280999 483444
rect 280933 483379 280999 483380
rect 280936 483202 280996 483379
rect 283656 483202 283716 483790
rect 286104 483202 286164 483790
rect 288552 483790 288634 483850
rect 290966 483850 291026 486099
rect 293514 485308 294134 510618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 295931 486164 295997 486165
rect 295931 486100 295932 486164
rect 295996 486100 295997 486164
rect 295931 486099 295997 486100
rect 293539 484940 293605 484941
rect 293539 484876 293540 484940
rect 293604 484876 293605 484940
rect 293539 484875 293605 484876
rect 293542 483850 293602 484875
rect 295934 483850 295994 486099
rect 297234 485308 297854 514338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300715 486028 300781 486029
rect 300715 485964 300716 486028
rect 300780 485964 300781 486028
rect 300715 485963 300781 485964
rect 300718 485210 300778 485963
rect 300954 485308 301574 518058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 307794 485308 308414 488898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311019 485892 311085 485893
rect 311019 485828 311020 485892
rect 311084 485828 311085 485892
rect 311019 485827 311085 485828
rect 300718 485150 300962 485210
rect 290966 483790 291060 483850
rect 293542 483790 293644 483850
rect 288552 483202 288612 483790
rect 291000 483202 291060 483790
rect 293584 483202 293644 483790
rect 295896 483790 295994 483850
rect 300902 483850 300962 485150
rect 305867 484804 305933 484805
rect 305867 484740 305868 484804
rect 305932 484740 305933 484804
rect 305867 484739 305933 484740
rect 303475 483852 303541 483853
rect 300902 483790 301124 483850
rect 295896 483202 295956 483790
rect 298613 483444 298679 483445
rect 298613 483380 298614 483444
rect 298678 483380 298679 483444
rect 298613 483379 298679 483380
rect 298616 483202 298676 483379
rect 301064 483202 301124 483790
rect 303475 483788 303476 483852
rect 303540 483850 303541 483852
rect 305870 483850 305930 484739
rect 311022 483850 311082 485827
rect 311514 485308 312134 492618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 313595 485892 313661 485893
rect 313595 485828 313596 485892
rect 313660 485828 313661 485892
rect 313595 485827 313661 485828
rect 313598 483850 313658 485827
rect 315234 485308 315854 496338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318379 486980 318445 486981
rect 318379 486916 318380 486980
rect 318444 486916 318445 486980
rect 318379 486915 318445 486916
rect 315803 484532 315869 484533
rect 315803 484468 315804 484532
rect 315868 484468 315869 484532
rect 315803 484467 315869 484468
rect 303540 483788 303572 483850
rect 305870 483790 306020 483850
rect 303475 483787 303572 483788
rect 303512 483202 303572 483787
rect 305960 483202 306020 483790
rect 310992 483790 311082 483850
rect 313576 483790 313658 483850
rect 315806 483850 315866 484467
rect 318382 483850 318442 486915
rect 318954 485308 319574 500058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 323347 486436 323413 486437
rect 323347 486372 323348 486436
rect 323412 486372 323413 486436
rect 323347 486371 323413 486372
rect 320955 485892 321021 485893
rect 320955 485828 320956 485892
rect 321020 485828 321021 485892
rect 320955 485827 321021 485828
rect 320958 483850 321018 485827
rect 323350 483850 323410 486371
rect 325794 485308 326414 506898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 329514 485308 330134 510618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 485308 333854 514338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 485308 337574 518058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 339723 486572 339789 486573
rect 339723 486508 339724 486572
rect 339788 486508 339789 486572
rect 339723 486507 339789 486508
rect 338435 484532 338501 484533
rect 338435 484468 338436 484532
rect 338500 484468 338501 484532
rect 338435 484467 338501 484468
rect 338438 483850 338498 484467
rect 339726 483850 339786 486507
rect 343794 485308 344414 488898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 485308 348134 492618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 350763 486436 350829 486437
rect 350763 486372 350764 486436
rect 350828 486372 350829 486436
rect 350763 486371 350829 486372
rect 315806 483790 316084 483850
rect 318382 483790 318532 483850
rect 320958 483790 321116 483850
rect 323350 483790 323428 483850
rect 338438 483790 338524 483850
rect 308405 483716 308471 483717
rect 308405 483652 308406 483716
rect 308470 483652 308471 483716
rect 308405 483651 308471 483652
rect 308408 483202 308468 483651
rect 310992 483202 311052 483790
rect 313576 483202 313636 483790
rect 316024 483202 316084 483790
rect 318472 483202 318532 483790
rect 321056 483202 321116 483790
rect 323368 483202 323428 483790
rect 326085 483580 326151 483581
rect 326085 483516 326086 483580
rect 326150 483516 326151 483580
rect 326085 483515 326151 483516
rect 326088 483202 326148 483515
rect 338464 483202 338524 483790
rect 339688 483790 339786 483850
rect 350766 483850 350826 486371
rect 351234 485308 351854 496338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 485308 355574 500058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 350766 483790 350900 483850
rect 339688 483202 339748 483790
rect 350840 483202 350900 483790
rect 220952 471454 221300 471486
rect 220952 471218 221008 471454
rect 221244 471218 221300 471454
rect 220952 471134 221300 471218
rect 220952 470898 221008 471134
rect 221244 470898 221300 471134
rect 220952 470866 221300 470898
rect 355320 471454 355668 471486
rect 355320 471218 355376 471454
rect 355612 471218 355668 471454
rect 355320 471134 355668 471218
rect 355320 470898 355376 471134
rect 355612 470898 355668 471134
rect 355320 470866 355668 470898
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 220272 453454 220620 453486
rect 220272 453218 220328 453454
rect 220564 453218 220620 453454
rect 220272 453134 220620 453218
rect 220272 452898 220328 453134
rect 220564 452898 220620 453134
rect 220272 452866 220620 452898
rect 356000 453454 356348 453486
rect 356000 453218 356056 453454
rect 356292 453218 356348 453454
rect 356000 453134 356348 453218
rect 356000 452898 356056 453134
rect 356292 452898 356348 453134
rect 356000 452866 356348 452898
rect 220952 435454 221300 435486
rect 220952 435218 221008 435454
rect 221244 435218 221300 435454
rect 220952 435134 221300 435218
rect 220952 434898 221008 435134
rect 221244 434898 221300 435134
rect 220952 434866 221300 434898
rect 355320 435454 355668 435486
rect 355320 435218 355376 435454
rect 355612 435218 355668 435454
rect 355320 435134 355668 435218
rect 355320 434898 355376 435134
rect 355612 434898 355668 435134
rect 355320 434866 355668 434898
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 220272 417454 220620 417486
rect 220272 417218 220328 417454
rect 220564 417218 220620 417454
rect 220272 417134 220620 417218
rect 220272 416898 220328 417134
rect 220564 416898 220620 417134
rect 220272 416866 220620 416898
rect 356000 417454 356348 417486
rect 356000 417218 356056 417454
rect 356292 417218 356348 417454
rect 356000 417134 356348 417218
rect 356000 416898 356056 417134
rect 356292 416898 356348 417134
rect 356000 416866 356348 416898
rect 236056 399530 236116 400106
rect 237144 399530 237204 400106
rect 238232 399530 238292 400106
rect 239592 399530 239652 400106
rect 235950 399470 236116 399530
rect 237054 399470 237204 399530
rect 238158 399470 238292 399530
rect 239262 399470 239652 399530
rect 240544 399530 240604 400106
rect 241768 399530 241828 400106
rect 243128 399530 243188 400106
rect 240544 399470 240610 399530
rect 235950 398173 236010 399470
rect 223803 398172 223869 398173
rect 223803 398108 223804 398172
rect 223868 398108 223869 398172
rect 223803 398107 223869 398108
rect 235947 398172 236013 398173
rect 235947 398108 235948 398172
rect 236012 398108 236013 398172
rect 235947 398107 236013 398108
rect 223619 398036 223685 398037
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 228924 211574 248058
rect 217794 363454 218414 398000
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 228924 218414 254898
rect 221514 367174 222134 398000
rect 223619 397972 223620 398036
rect 223684 397972 223685 398036
rect 223619 397971 223685 397972
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 221514 228924 222134 258618
rect 64208 219454 64528 219486
rect 64208 219218 64250 219454
rect 64486 219218 64528 219454
rect 64208 219134 64528 219218
rect 64208 218898 64250 219134
rect 64486 218898 64528 219134
rect 64208 218866 64528 218898
rect 94928 219454 95248 219486
rect 94928 219218 94970 219454
rect 95206 219218 95248 219454
rect 94928 219134 95248 219218
rect 94928 218898 94970 219134
rect 95206 218898 95248 219134
rect 94928 218866 95248 218898
rect 125648 219454 125968 219486
rect 125648 219218 125690 219454
rect 125926 219218 125968 219454
rect 125648 219134 125968 219218
rect 125648 218898 125690 219134
rect 125926 218898 125968 219134
rect 125648 218866 125968 218898
rect 156368 219454 156688 219486
rect 156368 219218 156410 219454
rect 156646 219218 156688 219454
rect 156368 219134 156688 219218
rect 156368 218898 156410 219134
rect 156646 218898 156688 219134
rect 156368 218866 156688 218898
rect 187088 219454 187408 219486
rect 187088 219218 187130 219454
rect 187366 219218 187408 219454
rect 187088 219134 187408 219218
rect 187088 218898 187130 219134
rect 187366 218898 187408 219134
rect 187088 218866 187408 218898
rect 217808 219454 218128 219486
rect 217808 219218 217850 219454
rect 218086 219218 218128 219454
rect 217808 219134 218128 219218
rect 217808 218898 217850 219134
rect 218086 218898 218128 219134
rect 217808 218866 218128 218898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 79568 201454 79888 201486
rect 79568 201218 79610 201454
rect 79846 201218 79888 201454
rect 79568 201134 79888 201218
rect 79568 200898 79610 201134
rect 79846 200898 79888 201134
rect 79568 200866 79888 200898
rect 110288 201454 110608 201486
rect 110288 201218 110330 201454
rect 110566 201218 110608 201454
rect 110288 201134 110608 201218
rect 110288 200898 110330 201134
rect 110566 200898 110608 201134
rect 110288 200866 110608 200898
rect 141008 201454 141328 201486
rect 141008 201218 141050 201454
rect 141286 201218 141328 201454
rect 141008 201134 141328 201218
rect 141008 200898 141050 201134
rect 141286 200898 141328 201134
rect 141008 200866 141328 200898
rect 171728 201454 172048 201486
rect 171728 201218 171770 201454
rect 172006 201218 172048 201454
rect 171728 201134 172048 201218
rect 171728 200898 171770 201134
rect 172006 200898 172048 201134
rect 171728 200866 172048 200898
rect 202448 201454 202768 201486
rect 202448 201218 202490 201454
rect 202726 201218 202768 201454
rect 202448 201134 202768 201218
rect 202448 200898 202490 201134
rect 202726 200898 202768 201134
rect 202448 200866 202768 200898
rect 64208 183454 64528 183486
rect 64208 183218 64250 183454
rect 64486 183218 64528 183454
rect 64208 183134 64528 183218
rect 64208 182898 64250 183134
rect 64486 182898 64528 183134
rect 64208 182866 64528 182898
rect 94928 183454 95248 183486
rect 94928 183218 94970 183454
rect 95206 183218 95248 183454
rect 94928 183134 95248 183218
rect 94928 182898 94970 183134
rect 95206 182898 95248 183134
rect 94928 182866 95248 182898
rect 125648 183454 125968 183486
rect 125648 183218 125690 183454
rect 125926 183218 125968 183454
rect 125648 183134 125968 183218
rect 125648 182898 125690 183134
rect 125926 182898 125968 183134
rect 125648 182866 125968 182898
rect 156368 183454 156688 183486
rect 156368 183218 156410 183454
rect 156646 183218 156688 183454
rect 156368 183134 156688 183218
rect 156368 182898 156410 183134
rect 156646 182898 156688 183134
rect 156368 182866 156688 182898
rect 187088 183454 187408 183486
rect 187088 183218 187130 183454
rect 187366 183218 187408 183454
rect 187088 183134 187408 183218
rect 187088 182898 187130 183134
rect 187366 182898 187408 183134
rect 187088 182866 187408 182898
rect 217808 183454 218128 183486
rect 217808 183218 217850 183454
rect 218086 183218 218128 183454
rect 217808 183134 218128 183218
rect 217808 182898 217850 183134
rect 218086 182898 218128 183134
rect 217808 182866 218128 182898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 79568 165454 79888 165486
rect 79568 165218 79610 165454
rect 79846 165218 79888 165454
rect 79568 165134 79888 165218
rect 79568 164898 79610 165134
rect 79846 164898 79888 165134
rect 79568 164866 79888 164898
rect 110288 165454 110608 165486
rect 110288 165218 110330 165454
rect 110566 165218 110608 165454
rect 110288 165134 110608 165218
rect 110288 164898 110330 165134
rect 110566 164898 110608 165134
rect 110288 164866 110608 164898
rect 141008 165454 141328 165486
rect 141008 165218 141050 165454
rect 141286 165218 141328 165454
rect 141008 165134 141328 165218
rect 141008 164898 141050 165134
rect 141286 164898 141328 165134
rect 141008 164866 141328 164898
rect 171728 165454 172048 165486
rect 171728 165218 171770 165454
rect 172006 165218 172048 165454
rect 171728 165134 172048 165218
rect 171728 164898 171770 165134
rect 172006 164898 172048 165134
rect 171728 164866 172048 164898
rect 202448 165454 202768 165486
rect 202448 165218 202490 165454
rect 202726 165218 202768 165454
rect 202448 165134 202768 165218
rect 202448 164898 202490 165134
rect 202726 164898 202768 165134
rect 202448 164866 202768 164898
rect 64208 147454 64528 147486
rect 64208 147218 64250 147454
rect 64486 147218 64528 147454
rect 64208 147134 64528 147218
rect 64208 146898 64250 147134
rect 64486 146898 64528 147134
rect 64208 146866 64528 146898
rect 94928 147454 95248 147486
rect 94928 147218 94970 147454
rect 95206 147218 95248 147454
rect 94928 147134 95248 147218
rect 94928 146898 94970 147134
rect 95206 146898 95248 147134
rect 94928 146866 95248 146898
rect 125648 147454 125968 147486
rect 125648 147218 125690 147454
rect 125926 147218 125968 147454
rect 125648 147134 125968 147218
rect 125648 146898 125690 147134
rect 125926 146898 125968 147134
rect 125648 146866 125968 146898
rect 156368 147454 156688 147486
rect 156368 147218 156410 147454
rect 156646 147218 156688 147454
rect 156368 147134 156688 147218
rect 156368 146898 156410 147134
rect 156646 146898 156688 147134
rect 156368 146866 156688 146898
rect 187088 147454 187408 147486
rect 187088 147218 187130 147454
rect 187366 147218 187408 147454
rect 187088 147134 187408 147218
rect 187088 146898 187130 147134
rect 187366 146898 187408 147134
rect 187088 146866 187408 146898
rect 217808 147454 218128 147486
rect 217808 147218 217850 147454
rect 218086 147218 218128 147454
rect 217808 147134 218128 147218
rect 217808 146898 217850 147134
rect 218086 146898 218128 147134
rect 217808 146866 218128 146898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 79568 129454 79888 129486
rect 79568 129218 79610 129454
rect 79846 129218 79888 129454
rect 79568 129134 79888 129218
rect 79568 128898 79610 129134
rect 79846 128898 79888 129134
rect 79568 128866 79888 128898
rect 110288 129454 110608 129486
rect 110288 129218 110330 129454
rect 110566 129218 110608 129454
rect 110288 129134 110608 129218
rect 110288 128898 110330 129134
rect 110566 128898 110608 129134
rect 110288 128866 110608 128898
rect 141008 129454 141328 129486
rect 141008 129218 141050 129454
rect 141286 129218 141328 129454
rect 141008 129134 141328 129218
rect 141008 128898 141050 129134
rect 141286 128898 141328 129134
rect 141008 128866 141328 128898
rect 171728 129454 172048 129486
rect 171728 129218 171770 129454
rect 172006 129218 172048 129454
rect 171728 129134 172048 129218
rect 171728 128898 171770 129134
rect 172006 128898 172048 129134
rect 171728 128866 172048 128898
rect 202448 129454 202768 129486
rect 202448 129218 202490 129454
rect 202726 129218 202768 129454
rect 202448 129134 202768 129218
rect 202448 128898 202490 129134
rect 202726 128898 202768 129134
rect 202448 128866 202768 128898
rect 64208 111454 64528 111486
rect 64208 111218 64250 111454
rect 64486 111218 64528 111454
rect 64208 111134 64528 111218
rect 64208 110898 64250 111134
rect 64486 110898 64528 111134
rect 64208 110866 64528 110898
rect 94928 111454 95248 111486
rect 94928 111218 94970 111454
rect 95206 111218 95248 111454
rect 94928 111134 95248 111218
rect 94928 110898 94970 111134
rect 95206 110898 95248 111134
rect 94928 110866 95248 110898
rect 125648 111454 125968 111486
rect 125648 111218 125690 111454
rect 125926 111218 125968 111454
rect 125648 111134 125968 111218
rect 125648 110898 125690 111134
rect 125926 110898 125968 111134
rect 125648 110866 125968 110898
rect 156368 111454 156688 111486
rect 156368 111218 156410 111454
rect 156646 111218 156688 111454
rect 156368 111134 156688 111218
rect 156368 110898 156410 111134
rect 156646 110898 156688 111134
rect 156368 110866 156688 110898
rect 187088 111454 187408 111486
rect 187088 111218 187130 111454
rect 187366 111218 187408 111454
rect 187088 111134 187408 111218
rect 187088 110898 187130 111134
rect 187366 110898 187408 111134
rect 187088 110866 187408 110898
rect 217808 111454 218128 111486
rect 217808 111218 217850 111454
rect 218086 111218 218128 111454
rect 217808 111134 218128 111218
rect 217808 110898 217850 111134
rect 218086 110898 218128 111134
rect 217808 110866 218128 110898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 79568 93454 79888 93486
rect 79568 93218 79610 93454
rect 79846 93218 79888 93454
rect 79568 93134 79888 93218
rect 79568 92898 79610 93134
rect 79846 92898 79888 93134
rect 79568 92866 79888 92898
rect 110288 93454 110608 93486
rect 110288 93218 110330 93454
rect 110566 93218 110608 93454
rect 110288 93134 110608 93218
rect 110288 92898 110330 93134
rect 110566 92898 110608 93134
rect 110288 92866 110608 92898
rect 141008 93454 141328 93486
rect 141008 93218 141050 93454
rect 141286 93218 141328 93454
rect 141008 93134 141328 93218
rect 141008 92898 141050 93134
rect 141286 92898 141328 93134
rect 141008 92866 141328 92898
rect 171728 93454 172048 93486
rect 171728 93218 171770 93454
rect 172006 93218 172048 93454
rect 171728 93134 172048 93218
rect 171728 92898 171770 93134
rect 172006 92898 172048 93134
rect 171728 92866 172048 92898
rect 202448 93454 202768 93486
rect 202448 93218 202490 93454
rect 202726 93218 202768 93454
rect 202448 93134 202768 93218
rect 202448 92898 202490 93134
rect 202726 92898 202768 93134
rect 202448 92866 202768 92898
rect 64208 75454 64528 75486
rect 64208 75218 64250 75454
rect 64486 75218 64528 75454
rect 64208 75134 64528 75218
rect 64208 74898 64250 75134
rect 64486 74898 64528 75134
rect 64208 74866 64528 74898
rect 94928 75454 95248 75486
rect 94928 75218 94970 75454
rect 95206 75218 95248 75454
rect 94928 75134 95248 75218
rect 94928 74898 94970 75134
rect 95206 74898 95248 75134
rect 94928 74866 95248 74898
rect 125648 75454 125968 75486
rect 125648 75218 125690 75454
rect 125926 75218 125968 75454
rect 125648 75134 125968 75218
rect 125648 74898 125690 75134
rect 125926 74898 125968 75134
rect 125648 74866 125968 74898
rect 156368 75454 156688 75486
rect 156368 75218 156410 75454
rect 156646 75218 156688 75454
rect 156368 75134 156688 75218
rect 156368 74898 156410 75134
rect 156646 74898 156688 75134
rect 156368 74866 156688 74898
rect 187088 75454 187408 75486
rect 187088 75218 187130 75454
rect 187366 75218 187408 75454
rect 187088 75134 187408 75218
rect 187088 74898 187130 75134
rect 187366 74898 187408 75134
rect 187088 74866 187408 74898
rect 217808 75454 218128 75486
rect 217808 75218 217850 75454
rect 218086 75218 218128 75454
rect 217808 75134 218128 75218
rect 217808 74898 217850 75134
rect 218086 74898 218128 75134
rect 217808 74866 218128 74898
rect 223067 60076 223133 60077
rect 223067 60012 223068 60076
rect 223132 60074 223133 60076
rect 223435 60076 223501 60077
rect 223435 60074 223436 60076
rect 223132 60014 223436 60074
rect 223132 60012 223133 60014
rect 223067 60011 223133 60012
rect 223435 60012 223436 60014
rect 223500 60012 223501 60076
rect 223435 60011 223501 60012
rect 223622 59941 223682 397971
rect 223619 59940 223685 59941
rect 223619 59876 223620 59940
rect 223684 59876 223685 59940
rect 223619 59875 223685 59876
rect 223806 59805 223866 398107
rect 224907 397900 224973 397901
rect 224907 397836 224908 397900
rect 224972 397836 224973 397900
rect 224907 397835 224973 397836
rect 224910 234565 224970 397835
rect 225234 370894 225854 398000
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 228954 374614 229574 398000
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 226379 322148 226445 322149
rect 226379 322084 226380 322148
rect 226444 322084 226445 322148
rect 226379 322083 226445 322084
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 224907 234564 224973 234565
rect 224907 234500 224908 234564
rect 224972 234500 224973 234564
rect 224907 234499 224973 234500
rect 224723 231028 224789 231029
rect 224723 230964 224724 231028
rect 224788 230964 224789 231028
rect 224723 230963 224789 230964
rect 224726 230210 224786 230963
rect 224726 230150 225154 230210
rect 224171 228852 224237 228853
rect 224171 228788 224172 228852
rect 224236 228788 224237 228852
rect 224171 228787 224237 228788
rect 224174 225861 224234 228787
rect 224171 225860 224237 225861
rect 224171 225796 224172 225860
rect 224236 225796 224237 225860
rect 224171 225795 224237 225796
rect 224907 225044 224973 225045
rect 224907 224980 224908 225044
rect 224972 224980 224973 225044
rect 224907 224979 224973 224980
rect 224910 60750 224970 224979
rect 224726 60690 224970 60750
rect 223803 59804 223869 59805
rect 223803 59740 223804 59804
rect 223868 59740 223869 59804
rect 223803 59739 223869 59740
rect 224726 59261 224786 60690
rect 225094 60077 225154 230150
rect 225234 228924 225854 262338
rect 226011 234564 226077 234565
rect 226011 234500 226012 234564
rect 226076 234500 226077 234564
rect 226011 234499 226077 234500
rect 226014 225450 226074 234499
rect 226195 231572 226261 231573
rect 226195 231508 226196 231572
rect 226260 231508 226261 231572
rect 226195 231507 226261 231508
rect 225830 225390 226074 225450
rect 225830 225045 225890 225390
rect 225827 225044 225893 225045
rect 225827 224980 225828 225044
rect 225892 224980 225893 225044
rect 225827 224979 225893 224980
rect 226198 224970 226258 231507
rect 226014 224910 226258 224970
rect 225091 60076 225157 60077
rect 225091 60012 225092 60076
rect 225156 60012 225157 60076
rect 225091 60011 225157 60012
rect 226014 59941 226074 224910
rect 226382 115157 226442 322083
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 226747 260132 226813 260133
rect 226747 260068 226748 260132
rect 226812 260068 226813 260132
rect 226747 260067 226813 260068
rect 226563 232796 226629 232797
rect 226563 232732 226564 232796
rect 226628 232732 226629 232796
rect 226563 232731 226629 232732
rect 226379 115156 226445 115157
rect 226379 115092 226380 115156
rect 226444 115092 226445 115156
rect 226379 115091 226445 115092
rect 226566 73541 226626 232731
rect 226750 107813 226810 260067
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 226931 229940 226997 229941
rect 226931 229876 226932 229940
rect 226996 229876 226997 229940
rect 226931 229875 226997 229876
rect 226747 107812 226813 107813
rect 226747 107748 226748 107812
rect 226812 107748 226813 107812
rect 226747 107747 226813 107748
rect 226934 80885 226994 229875
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 226931 80884 226997 80885
rect 226931 80820 226932 80884
rect 226996 80820 226997 80884
rect 226931 80819 226997 80820
rect 226563 73540 226629 73541
rect 226563 73476 226564 73540
rect 226628 73476 226629 73540
rect 226563 73475 226629 73476
rect 226011 59940 226077 59941
rect 226011 59876 226012 59940
rect 226076 59876 226077 59940
rect 226011 59875 226077 59876
rect 224723 59260 224789 59261
rect 224723 59196 224724 59260
rect 224788 59196 224789 59260
rect 224723 59195 224789 59196
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 58000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 58000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 58000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 58000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 58000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 381454 236414 398000
rect 237054 397357 237114 399470
rect 237051 397356 237117 397357
rect 237051 397292 237052 397356
rect 237116 397292 237117 397356
rect 237051 397291 237117 397292
rect 238158 396813 238218 399470
rect 239262 397357 239322 399470
rect 239259 397356 239325 397357
rect 239259 397292 239260 397356
rect 239324 397292 239325 397356
rect 239259 397291 239325 397292
rect 238155 396812 238221 396813
rect 238155 396748 238156 396812
rect 238220 396748 238221 396812
rect 238155 396747 238221 396748
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 385174 240134 398000
rect 240550 396813 240610 399470
rect 241654 399470 241828 399530
rect 242942 399470 243188 399530
rect 244216 399530 244276 400106
rect 245440 399530 245500 400106
rect 246528 399530 246588 400106
rect 244216 399470 244290 399530
rect 241654 396813 241714 399470
rect 242942 396813 243002 399470
rect 240547 396812 240613 396813
rect 240547 396748 240548 396812
rect 240612 396748 240613 396812
rect 240547 396747 240613 396748
rect 241651 396812 241717 396813
rect 241651 396748 241652 396812
rect 241716 396748 241717 396812
rect 241651 396747 241717 396748
rect 242939 396812 243005 396813
rect 242939 396748 242940 396812
rect 243004 396748 243005 396812
rect 242939 396747 243005 396748
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 277174 240134 312618
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 388894 243854 398000
rect 244230 396813 244290 399470
rect 245334 399470 245500 399530
rect 246438 399470 246588 399530
rect 247616 399530 247676 400106
rect 248296 399530 248356 400106
rect 248704 399530 248764 400106
rect 247616 399470 247786 399530
rect 245334 396813 245394 399470
rect 246438 396813 246498 399470
rect 244227 396812 244293 396813
rect 244227 396748 244228 396812
rect 244292 396748 244293 396812
rect 244227 396747 244293 396748
rect 245331 396812 245397 396813
rect 245331 396748 245332 396812
rect 245396 396748 245397 396812
rect 245331 396747 245397 396748
rect 246435 396812 246501 396813
rect 246435 396748 246436 396812
rect 246500 396748 246501 396812
rect 246435 396747 246501 396748
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 280894 243854 316338
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 392614 247574 398000
rect 247726 397357 247786 399470
rect 248278 399470 248356 399530
rect 248646 399470 248764 399530
rect 250064 399530 250124 400106
rect 250744 399530 250804 400106
rect 251288 399530 251348 400106
rect 252376 399530 252436 400106
rect 253464 399530 253524 400106
rect 250064 399470 250178 399530
rect 248278 397357 248338 399470
rect 248646 397357 248706 399470
rect 250118 397357 250178 399470
rect 250670 399470 250804 399530
rect 251222 399470 251348 399530
rect 252326 399470 252436 399530
rect 253430 399470 253524 399530
rect 253600 399530 253660 400106
rect 254552 399530 254612 400106
rect 255912 399530 255972 400106
rect 253600 399470 253674 399530
rect 250670 397357 250730 399470
rect 247723 397356 247789 397357
rect 247723 397292 247724 397356
rect 247788 397292 247789 397356
rect 247723 397291 247789 397292
rect 248275 397356 248341 397357
rect 248275 397292 248276 397356
rect 248340 397292 248341 397356
rect 248275 397291 248341 397292
rect 248643 397356 248709 397357
rect 248643 397292 248644 397356
rect 248708 397292 248709 397356
rect 248643 397291 248709 397292
rect 250115 397356 250181 397357
rect 250115 397292 250116 397356
rect 250180 397292 250181 397356
rect 250115 397291 250181 397292
rect 250667 397356 250733 397357
rect 250667 397292 250668 397356
rect 250732 397292 250733 397356
rect 250667 397291 250733 397292
rect 251222 397085 251282 399470
rect 251219 397084 251285 397085
rect 251219 397020 251220 397084
rect 251284 397020 251285 397084
rect 251219 397019 251285 397020
rect 252326 396813 252386 399470
rect 253430 397357 253490 399470
rect 253427 397356 253493 397357
rect 253427 397292 253428 397356
rect 253492 397292 253493 397356
rect 253427 397291 253493 397292
rect 253614 396813 253674 399470
rect 254534 399470 254612 399530
rect 255822 399470 255972 399530
rect 256048 399530 256108 400106
rect 257000 399530 257060 400106
rect 256048 399470 256250 399530
rect 252323 396812 252389 396813
rect 252323 396748 252324 396812
rect 252388 396748 252389 396812
rect 252323 396747 252389 396748
rect 253611 396812 253677 396813
rect 253611 396748 253612 396812
rect 253676 396748 253677 396812
rect 253611 396747 253677 396748
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 363454 254414 398000
rect 254534 396813 254594 399470
rect 255822 396813 255882 399470
rect 256190 396813 256250 399470
rect 256926 399470 257060 399530
rect 258088 399530 258148 400106
rect 258496 399530 258556 400106
rect 258088 399470 258274 399530
rect 256926 396813 256986 399470
rect 254531 396812 254597 396813
rect 254531 396748 254532 396812
rect 254596 396748 254597 396812
rect 254531 396747 254597 396748
rect 255819 396812 255885 396813
rect 255819 396748 255820 396812
rect 255884 396748 255885 396812
rect 255819 396747 255885 396748
rect 256187 396812 256253 396813
rect 256187 396748 256188 396812
rect 256252 396748 256253 396812
rect 256187 396747 256253 396748
rect 256923 396812 256989 396813
rect 256923 396748 256924 396812
rect 256988 396748 256989 396812
rect 256923 396747 256989 396748
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 367174 258134 398000
rect 258214 396810 258274 399470
rect 258398 399470 258556 399530
rect 259448 399530 259508 400106
rect 260672 399530 260732 400106
rect 261080 399530 261140 400106
rect 259448 399470 259562 399530
rect 258398 396949 258458 399470
rect 259502 397357 259562 399470
rect 260606 399470 260732 399530
rect 260974 399470 261140 399530
rect 261760 399530 261820 400106
rect 262848 399530 262908 400106
rect 261760 399470 262138 399530
rect 259499 397356 259565 397357
rect 259499 397292 259500 397356
rect 259564 397292 259565 397356
rect 259499 397291 259565 397292
rect 258395 396948 258461 396949
rect 258395 396884 258396 396948
rect 258460 396884 258461 396948
rect 258395 396883 258461 396884
rect 260606 396813 260666 399470
rect 260974 397357 261034 399470
rect 260971 397356 261037 397357
rect 260971 397292 260972 397356
rect 261036 397292 261037 397356
rect 260971 397291 261037 397292
rect 258395 396812 258461 396813
rect 258395 396810 258396 396812
rect 258214 396750 258396 396810
rect 258395 396748 258396 396750
rect 258460 396748 258461 396812
rect 258395 396747 258461 396748
rect 260603 396812 260669 396813
rect 260603 396748 260604 396812
rect 260668 396748 260669 396812
rect 260603 396747 260669 396748
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 370894 261854 398000
rect 262078 397357 262138 399470
rect 262814 399470 262908 399530
rect 263528 399530 263588 400106
rect 263936 399530 263996 400106
rect 265296 399530 265356 400106
rect 265976 399530 266036 400106
rect 266384 399530 266444 400106
rect 267608 399530 267668 400106
rect 263528 399470 263610 399530
rect 262814 397357 262874 399470
rect 262075 397356 262141 397357
rect 262075 397292 262076 397356
rect 262140 397292 262141 397356
rect 262075 397291 262141 397292
rect 262811 397356 262877 397357
rect 262811 397292 262812 397356
rect 262876 397292 262877 397356
rect 262811 397291 262877 397292
rect 263550 396813 263610 399470
rect 263918 399470 263996 399530
rect 265206 399470 265356 399530
rect 265942 399470 266036 399530
rect 266310 399470 266444 399530
rect 267598 399470 267668 399530
rect 268288 399530 268348 400106
rect 268696 399530 268756 400106
rect 269784 399530 269844 400106
rect 271008 399530 271068 400106
rect 268288 399470 268394 399530
rect 268696 399470 268762 399530
rect 269784 399470 269866 399530
rect 263918 397357 263978 399470
rect 265206 398173 265266 399470
rect 265203 398172 265269 398173
rect 265203 398108 265204 398172
rect 265268 398108 265269 398172
rect 265203 398107 265269 398108
rect 263915 397356 263981 397357
rect 263915 397292 263916 397356
rect 263980 397292 263981 397356
rect 263915 397291 263981 397292
rect 263547 396812 263613 396813
rect 263547 396748 263548 396812
rect 263612 396748 263613 396812
rect 263547 396747 263613 396748
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 374614 265574 398000
rect 265942 396813 266002 399470
rect 266310 396813 266370 399470
rect 265939 396812 266005 396813
rect 265939 396748 265940 396812
rect 266004 396748 266005 396812
rect 265939 396747 266005 396748
rect 266307 396812 266373 396813
rect 266307 396748 266308 396812
rect 266372 396748 266373 396812
rect 266307 396747 266373 396748
rect 267598 396677 267658 399470
rect 268334 397357 268394 399470
rect 268702 397357 268762 399470
rect 268331 397356 268397 397357
rect 268331 397292 268332 397356
rect 268396 397292 268397 397356
rect 268331 397291 268397 397292
rect 268699 397356 268765 397357
rect 268699 397292 268700 397356
rect 268764 397292 268765 397356
rect 268699 397291 268765 397292
rect 269806 396813 269866 399470
rect 270910 399470 271068 399530
rect 271144 399530 271204 400106
rect 272232 399530 272292 400106
rect 273320 399530 273380 400106
rect 273592 399530 273652 400106
rect 274408 399530 274468 400106
rect 275768 399530 275828 400106
rect 271144 399470 271338 399530
rect 272232 399470 272626 399530
rect 270910 396813 270970 399470
rect 269803 396812 269869 396813
rect 269803 396748 269804 396812
rect 269868 396748 269869 396812
rect 269803 396747 269869 396748
rect 270907 396812 270973 396813
rect 270907 396748 270908 396812
rect 270972 396748 270973 396812
rect 270907 396747 270973 396748
rect 271278 396677 271338 399470
rect 267595 396676 267661 396677
rect 267595 396612 267596 396676
rect 267660 396612 267661 396676
rect 267595 396611 267661 396612
rect 271275 396676 271341 396677
rect 271275 396612 271276 396676
rect 271340 396612 271341 396676
rect 271275 396611 271341 396612
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 381454 272414 398000
rect 272566 397357 272626 399470
rect 273302 399470 273380 399530
rect 273486 399470 273652 399530
rect 274406 399470 274468 399530
rect 275326 399470 275828 399530
rect 276040 399530 276100 400106
rect 276992 399530 277052 400106
rect 276040 399470 276306 399530
rect 272563 397356 272629 397357
rect 272563 397292 272564 397356
rect 272628 397292 272629 397356
rect 272563 397291 272629 397292
rect 273302 396813 273362 399470
rect 273299 396812 273365 396813
rect 273299 396748 273300 396812
rect 273364 396748 273365 396812
rect 273299 396747 273365 396748
rect 273486 396677 273546 399470
rect 274406 396813 274466 399470
rect 275326 397357 275386 399470
rect 275323 397356 275389 397357
rect 275323 397292 275324 397356
rect 275388 397292 275389 397356
rect 275323 397291 275389 397292
rect 274403 396812 274469 396813
rect 274403 396748 274404 396812
rect 274468 396748 274469 396812
rect 274403 396747 274469 396748
rect 273483 396676 273549 396677
rect 273483 396612 273484 396676
rect 273548 396612 273549 396676
rect 273483 396611 273549 396612
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 385174 276134 398000
rect 276246 396813 276306 399470
rect 276982 399470 277052 399530
rect 278080 399530 278140 400106
rect 278488 399530 278548 400106
rect 279168 399530 279228 400106
rect 280936 399530 280996 400106
rect 278080 399470 278146 399530
rect 276243 396812 276309 396813
rect 276243 396748 276244 396812
rect 276308 396748 276309 396812
rect 276243 396747 276309 396748
rect 276982 396677 277042 399470
rect 278086 397357 278146 399470
rect 278454 399470 278548 399530
rect 279006 399470 279228 399530
rect 280846 399470 280996 399530
rect 283520 399530 283580 400106
rect 285968 399530 286028 400106
rect 288280 399530 288340 400106
rect 291000 399530 291060 400106
rect 293448 399530 293508 400106
rect 283520 399470 283850 399530
rect 285968 399470 286058 399530
rect 278083 397356 278149 397357
rect 278083 397292 278084 397356
rect 278148 397292 278149 397356
rect 278083 397291 278149 397292
rect 278454 396813 278514 399470
rect 279006 397357 279066 399470
rect 279003 397356 279069 397357
rect 279003 397292 279004 397356
rect 279068 397292 279069 397356
rect 279003 397291 279069 397292
rect 278451 396812 278517 396813
rect 278451 396748 278452 396812
rect 278516 396748 278517 396812
rect 278451 396747 278517 396748
rect 276979 396676 277045 396677
rect 276979 396612 276980 396676
rect 277044 396612 277045 396676
rect 276979 396611 277045 396612
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 388894 279854 398000
rect 280846 396813 280906 399470
rect 280843 396812 280909 396813
rect 280843 396748 280844 396812
rect 280908 396748 280909 396812
rect 280843 396747 280909 396748
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 392614 283574 398000
rect 283790 396813 283850 399470
rect 285998 396813 286058 399470
rect 288206 399470 288340 399530
rect 290966 399470 291060 399530
rect 293358 399470 293508 399530
rect 295896 399530 295956 400106
rect 298480 399530 298540 400106
rect 300928 399530 300988 400106
rect 303512 399530 303572 400106
rect 305960 399530 306020 400106
rect 295896 399470 295994 399530
rect 298480 399470 298570 399530
rect 288206 396813 288266 399470
rect 283787 396812 283853 396813
rect 283787 396748 283788 396812
rect 283852 396748 283853 396812
rect 283787 396747 283853 396748
rect 285995 396812 286061 396813
rect 285995 396748 285996 396812
rect 286060 396748 286061 396812
rect 285995 396747 286061 396748
rect 288203 396812 288269 396813
rect 288203 396748 288204 396812
rect 288268 396748 288269 396812
rect 288203 396747 288269 396748
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 363454 290414 398000
rect 290966 397357 291026 399470
rect 290963 397356 291029 397357
rect 290963 397292 290964 397356
rect 291028 397292 291029 397356
rect 290963 397291 291029 397292
rect 293358 396813 293418 399470
rect 293355 396812 293421 396813
rect 293355 396748 293356 396812
rect 293420 396748 293421 396812
rect 293355 396747 293421 396748
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 367174 294134 398000
rect 295934 396813 295994 399470
rect 295931 396812 295997 396813
rect 295931 396748 295932 396812
rect 295996 396748 295997 396812
rect 295931 396747 295997 396748
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 370894 297854 398000
rect 298510 397357 298570 399470
rect 300902 399470 300988 399530
rect 303478 399470 303572 399530
rect 305870 399470 306020 399530
rect 308544 399530 308604 400106
rect 310992 399530 311052 400106
rect 313440 399530 313500 400106
rect 315888 399530 315948 400106
rect 318472 399530 318532 400106
rect 308544 399470 308690 399530
rect 310992 399470 311082 399530
rect 300902 398173 300962 399470
rect 300899 398172 300965 398173
rect 300899 398108 300900 398172
rect 300964 398108 300965 398172
rect 300899 398107 300965 398108
rect 298507 397356 298573 397357
rect 298507 397292 298508 397356
rect 298572 397292 298573 397356
rect 298507 397291 298573 397292
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 374614 301574 398000
rect 303478 396813 303538 399470
rect 305870 396813 305930 399470
rect 303475 396812 303541 396813
rect 303475 396748 303476 396812
rect 303540 396748 303541 396812
rect 303475 396747 303541 396748
rect 305867 396812 305933 396813
rect 305867 396748 305868 396812
rect 305932 396748 305933 396812
rect 305867 396747 305933 396748
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 381454 308414 398000
rect 308630 397357 308690 399470
rect 308627 397356 308693 397357
rect 308627 397292 308628 397356
rect 308692 397292 308693 397356
rect 308627 397291 308693 397292
rect 311022 396813 311082 399470
rect 313414 399470 313500 399530
rect 315806 399470 315948 399530
rect 318382 399470 318532 399530
rect 320920 399530 320980 400106
rect 323368 399530 323428 400106
rect 325952 399530 326012 400106
rect 343224 399530 343284 400106
rect 320920 399470 321018 399530
rect 311019 396812 311085 396813
rect 311019 396748 311020 396812
rect 311084 396748 311085 396812
rect 311019 396747 311085 396748
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 385174 312134 398000
rect 313414 396813 313474 399470
rect 315806 398173 315866 399470
rect 315803 398172 315869 398173
rect 315803 398108 315804 398172
rect 315868 398108 315869 398172
rect 315803 398107 315869 398108
rect 313411 396812 313477 396813
rect 313411 396748 313412 396812
rect 313476 396748 313477 396812
rect 313411 396747 313477 396748
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 388894 315854 398000
rect 318382 396813 318442 399470
rect 318379 396812 318445 396813
rect 318379 396748 318380 396812
rect 318444 396748 318445 396812
rect 318379 396747 318445 396748
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 392614 319574 398000
rect 320958 396813 321018 399470
rect 323350 399470 323428 399530
rect 325926 399470 326012 399530
rect 343222 399470 343284 399530
rect 343360 399530 343420 400106
rect 343360 399470 343466 399530
rect 323350 396813 323410 399470
rect 325926 398173 325986 399470
rect 325923 398172 325989 398173
rect 325923 398108 325924 398172
rect 325988 398108 325989 398172
rect 325923 398107 325989 398108
rect 320955 396812 321021 396813
rect 320955 396748 320956 396812
rect 321020 396748 321021 396812
rect 320955 396747 321021 396748
rect 323347 396812 323413 396813
rect 323347 396748 323348 396812
rect 323412 396748 323413 396812
rect 323347 396747 323413 396748
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 363454 326414 398000
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 367174 330134 398000
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 370894 333854 398000
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 374614 337574 398000
rect 343222 397357 343282 399470
rect 343219 397356 343285 397357
rect 343219 397292 343220 397356
rect 343284 397292 343285 397356
rect 343219 397291 343285 397292
rect 343406 396813 343466 399470
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 343403 396812 343469 396813
rect 343403 396748 343404 396812
rect 343468 396748 343469 396812
rect 343403 396747 343469 396748
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 381454 344414 398000
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 385174 348134 398000
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 388894 351854 398000
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 392614 355574 398000
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 61008 471218 61244 471454
rect 61008 470898 61244 471134
rect 195376 471218 195612 471454
rect 195376 470898 195612 471134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 60328 453218 60564 453454
rect 60328 452898 60564 453134
rect 196056 453218 196292 453454
rect 196056 452898 196292 453134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 61008 435218 61244 435454
rect 61008 434898 61244 435134
rect 195376 435218 195612 435454
rect 195376 434898 195612 435134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 60328 417218 60564 417454
rect 60328 416898 60564 417134
rect 196056 417218 196292 417454
rect 196056 416898 196292 417134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 221008 471218 221244 471454
rect 221008 470898 221244 471134
rect 355376 471218 355612 471454
rect 355376 470898 355612 471134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 220328 453218 220564 453454
rect 220328 452898 220564 453134
rect 356056 453218 356292 453454
rect 356056 452898 356292 453134
rect 221008 435218 221244 435454
rect 221008 434898 221244 435134
rect 355376 435218 355612 435454
rect 355376 434898 355612 435134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 220328 417218 220564 417454
rect 220328 416898 220564 417134
rect 356056 417218 356292 417454
rect 356056 416898 356292 417134
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 64250 219218 64486 219454
rect 64250 218898 64486 219134
rect 94970 219218 95206 219454
rect 94970 218898 95206 219134
rect 125690 219218 125926 219454
rect 125690 218898 125926 219134
rect 156410 219218 156646 219454
rect 156410 218898 156646 219134
rect 187130 219218 187366 219454
rect 187130 218898 187366 219134
rect 217850 219218 218086 219454
rect 217850 218898 218086 219134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 79610 201218 79846 201454
rect 79610 200898 79846 201134
rect 110330 201218 110566 201454
rect 110330 200898 110566 201134
rect 141050 201218 141286 201454
rect 141050 200898 141286 201134
rect 171770 201218 172006 201454
rect 171770 200898 172006 201134
rect 202490 201218 202726 201454
rect 202490 200898 202726 201134
rect 64250 183218 64486 183454
rect 64250 182898 64486 183134
rect 94970 183218 95206 183454
rect 94970 182898 95206 183134
rect 125690 183218 125926 183454
rect 125690 182898 125926 183134
rect 156410 183218 156646 183454
rect 156410 182898 156646 183134
rect 187130 183218 187366 183454
rect 187130 182898 187366 183134
rect 217850 183218 218086 183454
rect 217850 182898 218086 183134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 79610 165218 79846 165454
rect 79610 164898 79846 165134
rect 110330 165218 110566 165454
rect 110330 164898 110566 165134
rect 141050 165218 141286 165454
rect 141050 164898 141286 165134
rect 171770 165218 172006 165454
rect 171770 164898 172006 165134
rect 202490 165218 202726 165454
rect 202490 164898 202726 165134
rect 64250 147218 64486 147454
rect 64250 146898 64486 147134
rect 94970 147218 95206 147454
rect 94970 146898 95206 147134
rect 125690 147218 125926 147454
rect 125690 146898 125926 147134
rect 156410 147218 156646 147454
rect 156410 146898 156646 147134
rect 187130 147218 187366 147454
rect 187130 146898 187366 147134
rect 217850 147218 218086 147454
rect 217850 146898 218086 147134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 79610 129218 79846 129454
rect 79610 128898 79846 129134
rect 110330 129218 110566 129454
rect 110330 128898 110566 129134
rect 141050 129218 141286 129454
rect 141050 128898 141286 129134
rect 171770 129218 172006 129454
rect 171770 128898 172006 129134
rect 202490 129218 202726 129454
rect 202490 128898 202726 129134
rect 64250 111218 64486 111454
rect 64250 110898 64486 111134
rect 94970 111218 95206 111454
rect 94970 110898 95206 111134
rect 125690 111218 125926 111454
rect 125690 110898 125926 111134
rect 156410 111218 156646 111454
rect 156410 110898 156646 111134
rect 187130 111218 187366 111454
rect 187130 110898 187366 111134
rect 217850 111218 218086 111454
rect 217850 110898 218086 111134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 79610 93218 79846 93454
rect 79610 92898 79846 93134
rect 110330 93218 110566 93454
rect 110330 92898 110566 93134
rect 141050 93218 141286 93454
rect 141050 92898 141286 93134
rect 171770 93218 172006 93454
rect 171770 92898 172006 93134
rect 202490 93218 202726 93454
rect 202490 92898 202726 93134
rect 64250 75218 64486 75454
rect 64250 74898 64486 75134
rect 94970 75218 95206 75454
rect 94970 74898 95206 75134
rect 125690 75218 125926 75454
rect 125690 74898 125926 75134
rect 156410 75218 156646 75454
rect 156410 74898 156646 75134
rect 187130 75218 187366 75454
rect 187130 74898 187366 75134
rect 217850 75218 218086 75454
rect 217850 74898 218086 75134
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 61008 471454
rect 61244 471218 195376 471454
rect 195612 471218 221008 471454
rect 221244 471218 355376 471454
rect 355612 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 61008 471134
rect 61244 470898 195376 471134
rect 195612 470898 221008 471134
rect 221244 470898 355376 471134
rect 355612 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 60328 453454
rect 60564 453218 196056 453454
rect 196292 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 220328 453454
rect 220564 453218 356056 453454
rect 356292 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 60328 453134
rect 60564 452898 196056 453134
rect 196292 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 220328 453134
rect 220564 452898 356056 453134
rect 356292 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 61008 435454
rect 61244 435218 195376 435454
rect 195612 435218 221008 435454
rect 221244 435218 355376 435454
rect 355612 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 61008 435134
rect 61244 434898 195376 435134
rect 195612 434898 221008 435134
rect 221244 434898 355376 435134
rect 355612 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 60328 417454
rect 60564 417218 196056 417454
rect 196292 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 220328 417454
rect 220564 417218 356056 417454
rect 356292 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 60328 417134
rect 60564 416898 196056 417134
rect 196292 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 220328 417134
rect 220564 416898 356056 417134
rect 356292 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 64250 219454
rect 64486 219218 94970 219454
rect 95206 219218 125690 219454
rect 125926 219218 156410 219454
rect 156646 219218 187130 219454
rect 187366 219218 217850 219454
rect 218086 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 64250 219134
rect 64486 218898 94970 219134
rect 95206 218898 125690 219134
rect 125926 218898 156410 219134
rect 156646 218898 187130 219134
rect 187366 218898 217850 219134
rect 218086 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 79610 201454
rect 79846 201218 110330 201454
rect 110566 201218 141050 201454
rect 141286 201218 171770 201454
rect 172006 201218 202490 201454
rect 202726 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 79610 201134
rect 79846 200898 110330 201134
rect 110566 200898 141050 201134
rect 141286 200898 171770 201134
rect 172006 200898 202490 201134
rect 202726 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 64250 183454
rect 64486 183218 94970 183454
rect 95206 183218 125690 183454
rect 125926 183218 156410 183454
rect 156646 183218 187130 183454
rect 187366 183218 217850 183454
rect 218086 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 64250 183134
rect 64486 182898 94970 183134
rect 95206 182898 125690 183134
rect 125926 182898 156410 183134
rect 156646 182898 187130 183134
rect 187366 182898 217850 183134
rect 218086 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 79610 165454
rect 79846 165218 110330 165454
rect 110566 165218 141050 165454
rect 141286 165218 171770 165454
rect 172006 165218 202490 165454
rect 202726 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 79610 165134
rect 79846 164898 110330 165134
rect 110566 164898 141050 165134
rect 141286 164898 171770 165134
rect 172006 164898 202490 165134
rect 202726 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 64250 147454
rect 64486 147218 94970 147454
rect 95206 147218 125690 147454
rect 125926 147218 156410 147454
rect 156646 147218 187130 147454
rect 187366 147218 217850 147454
rect 218086 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 64250 147134
rect 64486 146898 94970 147134
rect 95206 146898 125690 147134
rect 125926 146898 156410 147134
rect 156646 146898 187130 147134
rect 187366 146898 217850 147134
rect 218086 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 79610 129454
rect 79846 129218 110330 129454
rect 110566 129218 141050 129454
rect 141286 129218 171770 129454
rect 172006 129218 202490 129454
rect 202726 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 79610 129134
rect 79846 128898 110330 129134
rect 110566 128898 141050 129134
rect 141286 128898 171770 129134
rect 172006 128898 202490 129134
rect 202726 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 64250 111454
rect 64486 111218 94970 111454
rect 95206 111218 125690 111454
rect 125926 111218 156410 111454
rect 156646 111218 187130 111454
rect 187366 111218 217850 111454
rect 218086 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 64250 111134
rect 64486 110898 94970 111134
rect 95206 110898 125690 111134
rect 125926 110898 156410 111134
rect 156646 110898 187130 111134
rect 187366 110898 217850 111134
rect 218086 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 79610 93454
rect 79846 93218 110330 93454
rect 110566 93218 141050 93454
rect 141286 93218 171770 93454
rect 172006 93218 202490 93454
rect 202726 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 79610 93134
rect 79846 92898 110330 93134
rect 110566 92898 141050 93134
rect 141286 92898 171770 93134
rect 172006 92898 202490 93134
rect 202726 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 64250 75454
rect 64486 75218 94970 75454
rect 95206 75218 125690 75454
rect 125926 75218 156410 75454
rect 156646 75218 187130 75454
rect 187366 75218 217850 75454
rect 218086 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 64250 75134
rect 64486 74898 94970 75134
rect 95206 74898 125690 75134
rect 125926 74898 156410 75134
rect 156646 74898 187130 75134
rect 187366 74898 217850 75134
rect 218086 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  sram1
timestamp 1640332777
transform 1 0 220000 0 1 400000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  sram
timestamp 1640332777
transform 1 0 60000 0 1 400000
box 0 0 136620 83308
use user_proj  mprj
timestamp 1640332777
transform 1 0 60000 0 1 60000
box 0 0 164780 166924
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 228924 74414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 228924 110414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 228924 146414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 228924 182414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 228924 218414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 485308 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 485308 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 485308 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 485308 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 485308 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 485308 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 485308 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 485308 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 228924 78134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 228924 114134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 228924 150134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 228924 186134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 228924 222134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 485308 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 485308 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 485308 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 485308 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 485308 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 485308 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 485308 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 485308 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 228924 81854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 228924 117854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 228924 153854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 228924 189854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 228924 225854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 485308 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 485308 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 485308 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 485308 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 485308 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 485308 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 485308 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 485308 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 228924 85574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 228924 121574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 228924 157574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 228924 193574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 485308 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 485308 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 485308 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 485308 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 485308 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 485308 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 485308 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 485308 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 228924 63854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 228924 99854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 228924 135854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 228924 171854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 485308 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 485308 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 485308 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 485308 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 228924 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 485308 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 485308 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 485308 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 485308 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 228924 67574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 228924 103574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 228924 139574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 228924 175574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 485308 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 485308 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 485308 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 485308 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 228924 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 485308 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 485308 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 485308 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 485308 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 228924 92414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 228924 128414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 228924 164414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 485308 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 485308 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 485308 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 228924 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 485308 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 485308 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 485308 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 485308 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 228924 60134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 228924 96134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 228924 132134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 228924 168134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 485308 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 485308 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 485308 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 485308 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 228924 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 485308 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 485308 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 485308 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 485308 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
