VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO user_proj
  CLASS BLOCK ;
  FOREIGN user_proj ;
  ORIGIN 0.000 0.000 ;
  SIZE 823.065 BY 833.785 ;
  PIN i_dout0[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 32.000 823.065 32.600 ;
    END
  END i_dout0[0]
  PIN i_dout0[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 446.800 4.000 447.400 ;
    END
  END i_dout0[10]
  PIN i_dout0[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 396.480 823.065 397.080 ;
    END
  END i_dout0[11]
  PIN i_dout0[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 686.410 0.000 686.690 4.000 ;
    END
  END i_dout0[12]
  PIN i_dout0[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 461.760 4.000 462.360 ;
    END
  END i_dout0[13]
  PIN i_dout0[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 507.320 4.000 507.920 ;
    END
  END i_dout0[14]
  PIN i_dout0[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 552.880 4.000 553.480 ;
    END
  END i_dout0[15]
  PIN i_dout0[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 702.050 829.785 702.330 833.785 ;
    END
  END i_dout0[16]
  PIN i_dout0[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 710.330 0.000 710.610 4.000 ;
    END
  END i_dout0[17]
  PIN i_dout0[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 552.880 823.065 553.480 ;
    END
  END i_dout0[18]
  PIN i_dout0[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 613.400 4.000 614.000 ;
    END
  END i_dout0[19]
  PIN i_dout0[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END i_dout0[1]
  PIN i_dout0[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 644.000 4.000 644.600 ;
    END
  END i_dout0[20]
  PIN i_dout0[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 4.000 ;
    END
  END i_dout0[21]
  PIN i_dout0[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 592.320 823.065 592.920 ;
    END
  END i_dout0[22]
  PIN i_dout0[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 605.240 823.065 605.840 ;
    END
  END i_dout0[23]
  PIN i_dout0[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.550 829.785 782.830 833.785 ;
    END
  END i_dout0[24]
  PIN i_dout0[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 762.770 0.000 763.050 4.000 ;
    END
  END i_dout0[25]
  PIN i_dout0[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 709.280 823.065 709.880 ;
    END
  END i_dout0[26]
  PIN i_dout0[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 748.040 823.065 748.640 ;
    END
  END i_dout0[27]
  PIN i_dout0[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 774.560 823.065 775.160 ;
    END
  END i_dout0[28]
  PIN i_dout0[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 750.080 4.000 750.680 ;
    END
  END i_dout0[29]
  PIN i_dout0[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 0.000 567.090 4.000 ;
    END
  END i_dout0[2]
  PIN i_dout0[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 829.785 815.950 833.785 ;
    END
  END i_dout0[30]
  PIN i_dout0[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 825.560 4.000 826.160 ;
    END
  END i_dout0[31]
  PIN i_dout0[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 189.080 4.000 189.680 ;
    END
  END i_dout0[3]
  PIN i_dout0[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 188.400 823.065 189.000 ;
    END
  END i_dout0[4]
  PIN i_dout0[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 249.600 4.000 250.200 ;
    END
  END i_dout0[5]
  PIN i_dout0[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 624.310 0.000 624.590 4.000 ;
    END
  END i_dout0[6]
  PIN i_dout0[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 253.000 823.065 253.600 ;
    END
  END i_dout0[7]
  PIN i_dout0[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 648.230 0.000 648.510 4.000 ;
    END
  END i_dout0[8]
  PIN i_dout0[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 635.810 829.785 636.090 833.785 ;
    END
  END i_dout0[9]
  PIN i_dout0_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 44.920 823.065 45.520 ;
    END
  END i_dout0_1[0]
  PIN i_dout0_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 645.470 829.785 645.750 833.785 ;
    END
  END i_dout0_1[10]
  PIN i_dout0_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 659.730 829.785 660.010 833.785 ;
    END
  END i_dout0_1[11]
  PIN i_dout0_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 668.930 829.785 669.210 833.785 ;
    END
  END i_dout0_1[12]
  PIN i_dout0_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 678.590 829.785 678.870 833.785 ;
    END
  END i_dout0_1[13]
  PIN i_dout0_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 477.400 4.000 478.000 ;
    END
  END i_dout0_1[14]
  PIN i_dout0_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 448.840 823.065 449.440 ;
    END
  END i_dout0_1[15]
  PIN i_dout0_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 697.450 829.785 697.730 833.785 ;
    END
  END i_dout0_1[16]
  PIN i_dout0_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END i_dout0_1[17]
  PIN i_dout0_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 720.910 829.785 721.190 833.785 ;
    END
  END i_dout0_1[18]
  PIN i_dout0_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 730.570 829.785 730.850 833.785 ;
    END
  END i_dout0_1[19]
  PIN i_dout0_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 113.600 4.000 114.200 ;
    END
  END i_dout0_1[1]
  PIN i_dout0_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 628.360 4.000 628.960 ;
    END
  END i_dout0_1[20]
  PIN i_dout0_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 578.720 823.065 579.320 ;
    END
  END i_dout0_1[21]
  PIN i_dout0_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 673.920 4.000 674.520 ;
    END
  END i_dout0_1[22]
  PIN i_dout0_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 768.290 829.785 768.570 833.785 ;
    END
  END i_dout0_1[23]
  PIN i_dout0_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 631.080 823.065 631.680 ;
    END
  END i_dout0_1[24]
  PIN i_dout0_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 656.920 823.065 657.520 ;
    END
  END i_dout0_1[25]
  PIN i_dout0_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 767.830 0.000 768.110 4.000 ;
    END
  END i_dout0_1[26]
  PIN i_dout0_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.430 0.000 772.710 4.000 ;
    END
  END i_dout0_1[27]
  PIN i_dout0_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 829.785 806.290 833.785 ;
    END
  END i_dout0_1[28]
  PIN i_dout0_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.350 0.000 796.630 4.000 ;
    END
  END i_dout0_1[29]
  PIN i_dout0_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 83.680 823.065 84.280 ;
    END
  END i_dout0_1[2]
  PIN i_dout0_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 811.070 829.785 811.350 833.785 ;
    END
  END i_dout0_1[30]
  PIN i_dout0_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 810.610 0.000 810.890 4.000 ;
    END
  END i_dout0_1[31]
  PIN i_dout0_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 174.120 4.000 174.720 ;
    END
  END i_dout0_1[3]
  PIN i_dout0_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 585.670 0.000 585.950 4.000 ;
    END
  END i_dout0_1[4]
  PIN i_dout0_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 219.680 4.000 220.280 ;
    END
  END i_dout0_1[5]
  PIN i_dout0_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 619.250 0.000 619.530 4.000 ;
    END
  END i_dout0_1[6]
  PIN i_dout0_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 240.080 823.065 240.680 ;
    END
  END i_dout0_1[7]
  PIN i_dout0_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 305.360 823.065 305.960 ;
    END
  END i_dout0_1[8]
  PIN i_dout0_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 370.640 823.065 371.240 ;
    END
  END i_dout0_1[9]
  PIN i_dout1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 523.570 0.000 523.850 4.000 ;
    END
  END i_dout1[0]
  PIN i_dout1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 650.070 829.785 650.350 833.785 ;
    END
  END i_dout1[10]
  PIN i_dout1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 409.400 823.065 410.000 ;
    END
  END i_dout1[11]
  PIN i_dout1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 691.010 0.000 691.290 4.000 ;
    END
  END i_dout1[12]
  PIN i_dout1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 687.790 829.785 688.070 833.785 ;
    END
  END i_dout1[13]
  PIN i_dout1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 522.280 4.000 522.880 ;
    END
  END i_dout1[14]
  PIN i_dout1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 474.680 823.065 475.280 ;
    END
  END i_dout1[15]
  PIN i_dout1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 706.650 829.785 706.930 833.785 ;
    END
  END i_dout1[16]
  PIN i_dout1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 539.960 823.065 540.560 ;
    END
  END i_dout1[17]
  PIN i_dout1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 583.480 4.000 584.080 ;
    END
  END i_dout1[18]
  PIN i_dout1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 739.770 829.785 740.050 833.785 ;
    END
  END i_dout1[19]
  PIN i_dout1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 829.785 550.990 833.785 ;
    END
  END i_dout1[1]
  PIN i_dout1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 724.590 0.000 724.870 4.000 ;
    END
  END i_dout1[20]
  PIN i_dout1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 749.430 829.785 749.710 833.785 ;
    END
  END i_dout1[21]
  PIN i_dout1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 748.510 0.000 748.790 4.000 ;
    END
  END i_dout1[22]
  PIN i_dout1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.950 829.785 778.230 833.785 ;
    END
  END i_dout1[23]
  PIN i_dout1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 644.000 823.065 644.600 ;
    END
  END i_dout1[24]
  PIN i_dout1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 683.440 823.065 684.040 ;
    END
  END i_dout1[25]
  PIN i_dout1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 704.520 4.000 705.120 ;
    END
  END i_dout1[26]
  PIN i_dout1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 719.480 4.000 720.080 ;
    END
  END i_dout1[27]
  PIN i_dout1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 787.480 823.065 788.080 ;
    END
  END i_dout1[28]
  PIN i_dout1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 765.040 4.000 765.640 ;
    END
  END i_dout1[29]
  PIN i_dout1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 571.410 0.000 571.690 4.000 ;
    END
  END i_dout1[2]
  PIN i_dout1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 795.640 4.000 796.240 ;
    END
  END i_dout1[30]
  PIN i_dout1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.270 829.785 820.550 833.785 ;
    END
  END i_dout1[31]
  PIN i_dout1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 588.430 829.785 588.710 833.785 ;
    END
  END i_dout1[3]
  PIN i_dout1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 607.750 829.785 608.030 833.785 ;
    END
  END i_dout1[4]
  PIN i_dout1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 227.160 823.065 227.760 ;
    END
  END i_dout1[5]
  PIN i_dout1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 4.000 ;
    END
  END i_dout1[6]
  PIN i_dout1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 638.570 0.000 638.850 4.000 ;
    END
  END i_dout1[7]
  PIN i_dout1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 631.210 829.785 631.490 833.785 ;
    END
  END i_dout1[8]
  PIN i_dout1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 657.430 0.000 657.710 4.000 ;
    END
  END i_dout1[9]
  PIN i_dout1_1[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.510 829.785 541.790 833.785 ;
    END
  END i_dout1_1[0]
  PIN i_dout1_1[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END i_dout1_1[10]
  PIN i_dout1_1[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 672.150 0.000 672.430 4.000 ;
    END
  END i_dout1_1[11]
  PIN i_dout1_1[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 681.350 0.000 681.630 4.000 ;
    END
  END i_dout1_1[12]
  PIN i_dout1_1[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 683.190 829.785 683.470 833.785 ;
    END
  END i_dout1_1[13]
  PIN i_dout1_1[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 492.360 4.000 492.960 ;
    END
  END i_dout1_1[14]
  PIN i_dout1_1[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 461.760 823.065 462.360 ;
    END
  END i_dout1_1[15]
  PIN i_dout1_1[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 500.520 823.065 501.120 ;
    END
  END i_dout1_1[16]
  PIN i_dout1_1[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 527.040 823.065 527.640 ;
    END
  END i_dout1_1[17]
  PIN i_dout1_1[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 567.840 4.000 568.440 ;
    END
  END i_dout1_1[18]
  PIN i_dout1_1[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 735.170 829.785 735.450 833.785 ;
    END
  END i_dout1_1[19]
  PIN i_dout1_1[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 128.560 4.000 129.160 ;
    END
  END i_dout1_1[1]
  PIN i_dout1_1[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 719.990 0.000 720.270 4.000 ;
    END
  END i_dout1_1[20]
  PIN i_dout1_1[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 658.960 4.000 659.560 ;
    END
  END i_dout1_1[21]
  PIN i_dout1_1[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 759.090 829.785 759.370 833.785 ;
    END
  END i_dout1_1[22]
  PIN i_dout1_1[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 772.890 829.785 773.170 833.785 ;
    END
  END i_dout1_1[23]
  PIN i_dout1_1[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 689.560 4.000 690.160 ;
    END
  END i_dout1_1[24]
  PIN i_dout1_1[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 669.840 823.065 670.440 ;
    END
  END i_dout1_1[25]
  PIN i_dout1_1[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 801.410 829.785 801.690 833.785 ;
    END
  END i_dout1_1[26]
  PIN i_dout1_1[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 777.030 0.000 777.310 4.000 ;
    END
  END i_dout1_1[27]
  PIN i_dout1_1[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 734.440 4.000 735.040 ;
    END
  END i_dout1_1[28]
  PIN i_dout1_1[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 800.950 0.000 801.230 4.000 ;
    END
  END i_dout1_1[29]
  PIN i_dout1_1[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 97.280 823.065 97.880 ;
    END
  END i_dout1_1[2]
  PIN i_dout1_1[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 800.400 823.065 801.000 ;
    END
  END i_dout1_1[30]
  PIN i_dout1_1[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 815.670 0.000 815.950 4.000 ;
    END
  END i_dout1_1[31]
  PIN i_dout1_1[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END i_dout1_1[3]
  PIN i_dout1_1[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 175.480 823.065 176.080 ;
    END
  END i_dout1_1[4]
  PIN i_dout1_1[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 234.640 4.000 235.240 ;
    END
  END i_dout1_1[5]
  PIN i_dout1_1[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END i_dout1_1[6]
  PIN i_dout1_1[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 355.680 4.000 356.280 ;
    END
  END i_dout1_1[7]
  PIN i_dout1_1[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 318.280 823.065 318.880 ;
    END
  END i_dout1_1[8]
  PIN i_dout1_1[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 383.560 823.065 384.160 ;
    END
  END i_dout1_1[9]
  PIN io_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 829.785 2.670 833.785 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.070 829.785 144.350 833.785 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 158.330 829.785 158.610 833.785 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 172.590 829.785 172.870 833.785 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.390 829.785 186.670 833.785 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 829.785 200.930 833.785 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.910 829.785 215.190 833.785 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 229.170 829.785 229.450 833.785 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 243.430 829.785 243.710 833.785 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 829.785 257.970 833.785 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 829.785 272.230 833.785 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 829.785 16.470 833.785 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 829.785 286.030 833.785 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 300.010 829.785 300.290 833.785 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 314.270 829.785 314.550 833.785 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 328.530 829.785 328.810 833.785 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 342.790 829.785 343.070 833.785 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.050 829.785 357.330 833.785 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.850 829.785 371.130 833.785 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 829.785 385.390 833.785 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 829.785 399.650 833.785 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 829.785 413.910 833.785 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 829.785 30.730 833.785 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 829.785 428.170 833.785 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 829.785 442.430 833.785 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.410 829.785 456.690 833.785 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 829.785 470.490 833.785 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 484.470 829.785 484.750 833.785 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 498.730 829.785 499.010 833.785 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.990 829.785 513.270 833.785 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 527.250 829.785 527.530 833.785 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.710 829.785 44.990 833.785 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.970 829.785 59.250 833.785 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 73.230 829.785 73.510 833.785 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.490 829.785 87.770 833.785 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.290 829.785 101.570 833.785 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 829.785 115.830 833.785 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.810 829.785 130.090 833.785 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 829.785 7.270 833.785 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.670 829.785 148.950 833.785 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 162.930 829.785 163.210 833.785 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 829.785 177.470 833.785 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 829.785 191.730 833.785 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.710 829.785 205.990 833.785 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.510 829.785 219.790 833.785 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 233.770 829.785 234.050 833.785 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 829.785 248.310 833.785 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.290 829.785 262.570 833.785 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 829.785 276.830 833.785 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 829.785 21.530 833.785 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.810 829.785 291.090 833.785 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 305.070 829.785 305.350 833.785 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 829.785 319.150 833.785 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 333.130 829.785 333.410 833.785 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.390 829.785 347.670 833.785 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.650 829.785 361.930 833.785 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.910 829.785 376.190 833.785 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 390.170 829.785 390.450 833.785 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 829.785 404.250 833.785 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 829.785 418.510 833.785 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 829.785 35.330 833.785 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.490 829.785 432.770 833.785 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 446.750 829.785 447.030 833.785 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.010 829.785 461.290 833.785 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.270 829.785 475.550 833.785 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 829.785 489.810 833.785 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 503.330 829.785 503.610 833.785 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 517.590 829.785 517.870 833.785 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 531.850 829.785 532.130 833.785 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 49.310 829.785 49.590 833.785 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 63.570 829.785 63.850 833.785 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.830 829.785 78.110 833.785 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.090 829.785 92.370 833.785 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 829.785 106.630 833.785 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.610 829.785 120.890 833.785 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 134.410 829.785 134.690 833.785 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 829.785 11.870 833.785 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 153.730 829.785 154.010 833.785 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 829.785 167.810 833.785 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 181.790 829.785 182.070 833.785 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 829.785 196.330 833.785 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 210.310 829.785 210.590 833.785 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 224.570 829.785 224.850 833.785 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.830 829.785 239.110 833.785 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 252.630 829.785 252.910 833.785 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 266.890 829.785 267.170 833.785 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 829.785 281.430 833.785 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 829.785 26.130 833.785 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 295.410 829.785 295.690 833.785 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.670 829.785 309.950 833.785 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 323.930 829.785 324.210 833.785 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.730 829.785 338.010 833.785 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.990 829.785 352.270 833.785 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 366.250 829.785 366.530 833.785 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.510 829.785 380.790 833.785 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.770 829.785 395.050 833.785 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 829.785 409.310 833.785 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 829.785 423.570 833.785 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.110 829.785 40.390 833.785 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.090 829.785 437.370 833.785 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.350 829.785 451.630 833.785 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 465.610 829.785 465.890 833.785 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 829.785 480.150 833.785 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 494.130 829.785 494.410 833.785 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 508.390 829.785 508.670 833.785 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 522.190 829.785 522.470 833.785 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 536.450 829.785 536.730 833.785 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.370 829.785 54.650 833.785 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 68.170 829.785 68.450 833.785 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 82.430 829.785 82.710 833.785 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 96.690 829.785 96.970 833.785 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 829.785 111.230 833.785 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.210 829.785 125.490 833.785 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 139.470 829.785 139.750 833.785 ;
    END
  END io_out[9]
  PIN irq[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END irq[0]
  PIN irq[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 513.910 0.000 514.190 4.000 ;
    END
  END irq[1]
  PIN irq[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.970 0.000 519.250 4.000 ;
    END
  END irq[2]
  PIN o_addr1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.630 0.000 528.910 4.000 ;
    END
  END o_addr1[0]
  PIN o_addr1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 552.550 0.000 552.830 4.000 ;
    END
  END o_addr1[1]
  PIN o_addr1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 110.200 823.065 110.800 ;
    END
  END o_addr1[2]
  PIN o_addr1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 136.040 823.065 136.640 ;
    END
  END o_addr1[3]
  PIN o_addr1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 201.320 823.065 201.920 ;
    END
  END o_addr1[4]
  PIN o_addr1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 614.650 0.000 614.930 4.000 ;
    END
  END o_addr1[5]
  PIN o_addr1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.160 4.000 295.760 ;
    END
  END o_addr1[6]
  PIN o_addr1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 643.170 0.000 643.450 4.000 ;
    END
  END o_addr1[7]
  PIN o_addr1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 652.830 0.000 653.110 4.000 ;
    END
  END o_addr1[8]
  PIN o_addr1_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END o_addr1_1[0]
  PIN o_addr1_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 57.840 823.065 58.440 ;
    END
  END o_addr1_1[1]
  PIN o_addr1_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 564.970 829.785 565.250 833.785 ;
    END
  END o_addr1_1[2]
  PIN o_addr1_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 581.070 0.000 581.350 4.000 ;
    END
  END o_addr1_1[3]
  PIN o_addr1_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 590.730 0.000 591.010 4.000 ;
    END
  END o_addr1_1[4]
  PIN o_addr1_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 609.590 0.000 609.870 4.000 ;
    END
  END o_addr1_1[5]
  PIN o_addr1_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.200 4.000 280.800 ;
    END
  END o_addr1_1[6]
  PIN o_addr1_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 370.640 4.000 371.240 ;
    END
  END o_addr1_1[7]
  PIN o_addr1_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 401.240 4.000 401.840 ;
    END
  END o_addr1_1[8]
  PIN o_csb0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 7.520 4.000 8.120 ;
    END
  END o_csb0
  PIN o_csb0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END o_csb0_1
  PIN o_csb1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 37.440 4.000 38.040 ;
    END
  END o_csb1
  PIN o_csb1_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 52.400 4.000 53.000 ;
    END
  END o_csb1_1
  PIN o_din0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 533.230 0.000 533.510 4.000 ;
    END
  END o_din0[0]
  PIN o_din0[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 667.090 0.000 667.370 4.000 ;
    END
  END o_din0[10]
  PIN o_din0[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 664.330 829.785 664.610 833.785 ;
    END
  END o_din0[11]
  PIN o_din0[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 673.530 829.785 673.810 833.785 ;
    END
  END o_din0[12]
  PIN o_din0[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 435.920 823.065 436.520 ;
    END
  END o_din0[13]
  PIN o_din0[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 692.850 829.785 693.130 833.785 ;
    END
  END o_din0[14]
  PIN o_din0[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 700.670 0.000 700.950 4.000 ;
    END
  END o_din0[15]
  PIN o_din0[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 711.710 829.785 711.990 833.785 ;
    END
  END o_din0[16]
  PIN o_din0[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 714.930 0.000 715.210 4.000 ;
    END
  END o_din0[17]
  PIN o_din0[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 598.440 4.000 599.040 ;
    END
  END o_din0[18]
  PIN o_din0[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 744.830 829.785 745.110 833.785 ;
    END
  END o_din0[19]
  PIN o_din0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 555.310 829.785 555.590 833.785 ;
    END
  END o_din0[1]
  PIN o_din0[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 734.250 0.000 734.530 4.000 ;
    END
  END o_din0[20]
  PIN o_din0[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 743.910 0.000 744.190 4.000 ;
    END
  END o_din0[21]
  PIN o_din0[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 763.690 829.785 763.970 833.785 ;
    END
  END o_din0[22]
  PIN o_din0[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 758.170 0.000 758.450 4.000 ;
    END
  END o_din0[23]
  PIN o_din0[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 792.210 829.785 792.490 833.785 ;
    END
  END o_din0[24]
  PIN o_din0[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 696.360 823.065 696.960 ;
    END
  END o_din0[25]
  PIN o_din0[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 735.120 823.065 735.720 ;
    END
  END o_din0[26]
  PIN o_din0[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 761.640 823.065 762.240 ;
    END
  END o_din0[27]
  PIN o_din0[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 791.750 0.000 792.030 4.000 ;
    END
  END o_din0[28]
  PIN o_din0[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 780.000 4.000 780.600 ;
    END
  END o_din0[29]
  PIN o_din0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 574.630 829.785 574.910 833.785 ;
    END
  END o_din0[2]
  PIN o_din0[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 810.600 4.000 811.200 ;
    END
  END o_din0[30]
  PIN o_din0[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 820.270 0.000 820.550 4.000 ;
    END
  END o_din0[31]
  PIN o_din0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 204.040 4.000 204.640 ;
    END
  END o_din0[3]
  PIN o_din0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 600.390 0.000 600.670 4.000 ;
    END
  END o_din0[4]
  PIN o_din0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 616.950 829.785 617.230 833.785 ;
    END
  END o_din0[5]
  PIN o_din0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 325.760 4.000 326.360 ;
    END
  END o_din0[6]
  PIN o_din0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 279.520 823.065 280.120 ;
    END
  END o_din0[7]
  PIN o_din0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 344.800 823.065 345.400 ;
    END
  END o_din0[8]
  PIN o_din0[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 640.870 829.785 641.150 833.785 ;
    END
  END o_din0[9]
  PIN o_din0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 0.000 538.110 4.000 ;
    END
  END o_din0_1[0]
  PIN o_din0_1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 654.670 829.785 654.950 833.785 ;
    END
  END o_din0_1[10]
  PIN o_din0_1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 676.750 0.000 677.030 4.000 ;
    END
  END o_din0_1[11]
  PIN o_din0_1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 696.070 0.000 696.350 4.000 ;
    END
  END o_din0_1[12]
  PIN o_din0_1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 423.000 823.065 423.600 ;
    END
  END o_din0_1[13]
  PIN o_din0_1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 537.920 4.000 538.520 ;
    END
  END o_din0_1[14]
  PIN o_din0_1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 487.600 823.065 488.200 ;
    END
  END o_din0_1[15]
  PIN o_din0_1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 514.120 823.065 514.720 ;
    END
  END o_din0_1[16]
  PIN o_din0_1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 716.310 829.785 716.590 833.785 ;
    END
  END o_din0_1[17]
  PIN o_din0_1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 725.970 829.785 726.250 833.785 ;
    END
  END o_din0_1[18]
  PIN o_din0_1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 565.800 823.065 566.400 ;
    END
  END o_din0_1[19]
  PIN o_din0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END o_din0_1[1]
  PIN o_din0_1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 729.190 0.000 729.470 4.000 ;
    END
  END o_din0_1[20]
  PIN o_din0_1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 754.030 829.785 754.310 833.785 ;
    END
  END o_din0_1[21]
  PIN o_din0_1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 753.110 0.000 753.390 4.000 ;
    END
  END o_din0_1[22]
  PIN o_din0_1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 618.160 823.065 618.760 ;
    END
  END o_din0_1[23]
  PIN o_din0_1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 787.150 829.785 787.430 833.785 ;
    END
  END o_din0_1[24]
  PIN o_din0_1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 796.810 829.785 797.090 833.785 ;
    END
  END o_din0_1[25]
  PIN o_din0_1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 722.200 823.065 722.800 ;
    END
  END o_din0_1[26]
  PIN o_din0_1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 4.000 ;
    END
  END o_din0_1[27]
  PIN o_din0_1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 786.690 0.000 786.970 4.000 ;
    END
  END o_din0_1[28]
  PIN o_din0_1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 806.010 0.000 806.290 4.000 ;
    END
  END o_din0_1[29]
  PIN o_din0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 569.570 829.785 569.850 833.785 ;
    END
  END o_din0_1[2]
  PIN o_din0_1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 813.320 823.065 813.920 ;
    END
  END o_din0_1[30]
  PIN o_din0_1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 826.240 823.065 826.840 ;
    END
  END o_din0_1[31]
  PIN o_din0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 148.960 823.065 149.560 ;
    END
  END o_din0_1[3]
  PIN o_din0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END o_din0_1[4]
  PIN o_din0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 612.350 829.785 612.630 833.785 ;
    END
  END o_din0_1[5]
  PIN o_din0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 310.120 4.000 310.720 ;
    END
  END o_din0_1[6]
  PIN o_din0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 266.600 823.065 267.200 ;
    END
  END o_din0_1[7]
  PIN o_din0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 331.200 823.065 331.800 ;
    END
  END o_din0_1[8]
  PIN o_din0_1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 431.840 4.000 432.440 ;
    END
  END o_din0_1[9]
  PIN o_waddr0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 546.110 829.785 546.390 833.785 ;
    END
  END o_waddr0[0]
  PIN o_waddr0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 70.760 823.065 71.360 ;
    END
  END o_waddr0[1]
  PIN o_waddr0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 123.120 823.065 123.720 ;
    END
  END o_waddr0[2]
  PIN o_waddr0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 598.090 829.785 598.370 833.785 ;
    END
  END o_waddr0[3]
  PIN o_waddr0[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 604.990 0.000 605.270 4.000 ;
    END
  END o_waddr0[4]
  PIN o_waddr0[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 626.610 829.785 626.890 833.785 ;
    END
  END o_waddr0[5]
  PIN o_waddr0[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.720 4.000 341.320 ;
    END
  END o_waddr0[6]
  PIN o_waddr0[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 386.280 4.000 386.880 ;
    END
  END o_waddr0[7]
  PIN o_waddr0[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 416.200 4.000 416.800 ;
    END
  END o_waddr0[8]
  PIN o_waddr0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END o_waddr0_1[0]
  PIN o_waddr0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 829.785 560.650 833.785 ;
    END
  END o_waddr0_1[1]
  PIN o_waddr0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.230 829.785 579.510 833.785 ;
    END
  END o_waddr0_1[2]
  PIN o_waddr0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 593.490 829.785 593.770 833.785 ;
    END
  END o_waddr0_1[3]
  PIN o_waddr0_1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 214.240 823.065 214.840 ;
    END
  END o_waddr0_1[4]
  PIN o_waddr0_1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 621.550 829.785 621.830 833.785 ;
    END
  END o_waddr0_1[5]
  PIN o_waddr0_1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 633.510 0.000 633.790 4.000 ;
    END
  END o_waddr0_1[6]
  PIN o_waddr0_1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 292.440 823.065 293.040 ;
    END
  END o_waddr0_1[7]
  PIN o_waddr0_1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 357.720 823.065 358.320 ;
    END
  END o_waddr0_1[8]
  PIN o_web0
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 6.160 823.065 6.760 ;
    END
  END o_web0
  PIN o_web0_1
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 19.080 823.065 19.680 ;
    END
  END o_web0_1
  PIN o_wmask0[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 83.000 4.000 83.600 ;
    END
  END o_wmask0[0]
  PIN o_wmask0[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 561.750 0.000 562.030 4.000 ;
    END
  END o_wmask0[1]
  PIN o_wmask0[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 583.830 829.785 584.110 833.785 ;
    END
  END o_wmask0[2]
  PIN o_wmask0[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 819.065 161.880 823.065 162.480 ;
    END
  END o_wmask0[3]
  PIN o_wmask0_1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END o_wmask0_1[0]
  PIN o_wmask0_1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END o_wmask0_1[1]
  PIN o_wmask0_1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 158.480 4.000 159.080 ;
    END
  END o_wmask0_1[2]
  PIN o_wmask0_1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 602.690 829.785 602.970 833.785 ;
    END
  END o_wmask0_1[3]
  PIN vccd1
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 635.440 10.640 637.040 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 789.040 10.640 790.640 821.680 ;
    END
  END vccd1
  PIN vssd1
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 821.680 ;
    END
    PORT
      LAYER met4 ;
        RECT 712.240 10.640 713.840 821.680 ;
    END
  END vssd1
  PIN wb_clk_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 2.390 0.000 2.670 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.990 0.000 7.270 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 11.590 0.000 11.870 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.910 0.000 31.190 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 0.000 194.030 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 208.010 0.000 208.290 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 0.000 222.550 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 250.790 0.000 251.070 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.510 0.000 265.790 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.030 0.000 294.310 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 308.290 0.000 308.570 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 337.270 0.000 337.550 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 351.530 0.000 351.810 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 365.790 0.000 366.070 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 0.000 380.330 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 394.310 0.000 394.590 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 0.000 409.310 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 423.290 0.000 423.570 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 437.550 0.000 437.830 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 451.810 0.000 452.090 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.070 0.000 466.350 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.090 0.000 69.370 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 480.790 0.000 481.070 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.050 0.000 495.330 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 88.410 0.000 88.690 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 107.270 0.000 107.550 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 121.990 0.000 122.270 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 0.000 136.530 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.510 0.000 150.790 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.770 0.000 165.050 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.030 0.000 179.310 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 0.000 35.790 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 0.000 198.630 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 226.870 0.000 227.150 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 0.000 256.130 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.110 0.000 270.390 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 284.370 0.000 284.650 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 298.630 0.000 298.910 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 327.610 0.000 327.890 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.870 0.000 342.150 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 385.110 0.000 385.390 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 413.630 0.000 413.910 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 427.890 0.000 428.170 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 456.870 0.000 457.150 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 471.130 0.000 471.410 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 485.390 0.000 485.670 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.650 0.000 499.930 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.330 0.000 112.610 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 155.110 0.000 155.390 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.090 0.000 184.370 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 40.570 0.000 40.850 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 217.670 0.000 217.950 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 231.930 0.000 232.210 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 0.000 260.730 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.710 0.000 274.990 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.430 0.000 289.710 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 303.690 0.000 303.970 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 317.950 0.000 318.230 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 346.470 0.000 346.750 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 361.190 0.000 361.470 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 375.450 0.000 375.730 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 403.970 0.000 404.250 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 418.230 0.000 418.510 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.210 0.000 447.490 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 461.470 0.000 461.750 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 0.000 79.030 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.990 0.000 490.270 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 504.710 0.000 504.990 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 98.070 0.000 98.350 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.930 0.000 117.210 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.190 0.000 131.470 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.910 0.000 146.190 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 160.170 0.000 160.450 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 174.430 0.000 174.710 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 188.690 0.000 188.970 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 0.000 83.630 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 102.670 0.000 102.950 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 0.000 21.530 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 26.310 0.000 26.590 4.000 ;
    END
  END wbs_we_i
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 822.795 821.525 ;
      LAYER met1 ;
        RECT 0.070 3.440 822.870 821.680 ;
      LAYER met2 ;
        RECT 0.100 829.505 2.110 830.010 ;
        RECT 2.950 829.505 6.710 830.010 ;
        RECT 7.550 829.505 11.310 830.010 ;
        RECT 12.150 829.505 15.910 830.010 ;
        RECT 16.750 829.505 20.970 830.010 ;
        RECT 21.810 829.505 25.570 830.010 ;
        RECT 26.410 829.505 30.170 830.010 ;
        RECT 31.010 829.505 34.770 830.010 ;
        RECT 35.610 829.505 39.830 830.010 ;
        RECT 40.670 829.505 44.430 830.010 ;
        RECT 45.270 829.505 49.030 830.010 ;
        RECT 49.870 829.505 54.090 830.010 ;
        RECT 54.930 829.505 58.690 830.010 ;
        RECT 59.530 829.505 63.290 830.010 ;
        RECT 64.130 829.505 67.890 830.010 ;
        RECT 68.730 829.505 72.950 830.010 ;
        RECT 73.790 829.505 77.550 830.010 ;
        RECT 78.390 829.505 82.150 830.010 ;
        RECT 82.990 829.505 87.210 830.010 ;
        RECT 88.050 829.505 91.810 830.010 ;
        RECT 92.650 829.505 96.410 830.010 ;
        RECT 97.250 829.505 101.010 830.010 ;
        RECT 101.850 829.505 106.070 830.010 ;
        RECT 106.910 829.505 110.670 830.010 ;
        RECT 111.510 829.505 115.270 830.010 ;
        RECT 116.110 829.505 120.330 830.010 ;
        RECT 121.170 829.505 124.930 830.010 ;
        RECT 125.770 829.505 129.530 830.010 ;
        RECT 130.370 829.505 134.130 830.010 ;
        RECT 134.970 829.505 139.190 830.010 ;
        RECT 140.030 829.505 143.790 830.010 ;
        RECT 144.630 829.505 148.390 830.010 ;
        RECT 149.230 829.505 153.450 830.010 ;
        RECT 154.290 829.505 158.050 830.010 ;
        RECT 158.890 829.505 162.650 830.010 ;
        RECT 163.490 829.505 167.250 830.010 ;
        RECT 168.090 829.505 172.310 830.010 ;
        RECT 173.150 829.505 176.910 830.010 ;
        RECT 177.750 829.505 181.510 830.010 ;
        RECT 182.350 829.505 186.110 830.010 ;
        RECT 186.950 829.505 191.170 830.010 ;
        RECT 192.010 829.505 195.770 830.010 ;
        RECT 196.610 829.505 200.370 830.010 ;
        RECT 201.210 829.505 205.430 830.010 ;
        RECT 206.270 829.505 210.030 830.010 ;
        RECT 210.870 829.505 214.630 830.010 ;
        RECT 215.470 829.505 219.230 830.010 ;
        RECT 220.070 829.505 224.290 830.010 ;
        RECT 225.130 829.505 228.890 830.010 ;
        RECT 229.730 829.505 233.490 830.010 ;
        RECT 234.330 829.505 238.550 830.010 ;
        RECT 239.390 829.505 243.150 830.010 ;
        RECT 243.990 829.505 247.750 830.010 ;
        RECT 248.590 829.505 252.350 830.010 ;
        RECT 253.190 829.505 257.410 830.010 ;
        RECT 258.250 829.505 262.010 830.010 ;
        RECT 262.850 829.505 266.610 830.010 ;
        RECT 267.450 829.505 271.670 830.010 ;
        RECT 272.510 829.505 276.270 830.010 ;
        RECT 277.110 829.505 280.870 830.010 ;
        RECT 281.710 829.505 285.470 830.010 ;
        RECT 286.310 829.505 290.530 830.010 ;
        RECT 291.370 829.505 295.130 830.010 ;
        RECT 295.970 829.505 299.730 830.010 ;
        RECT 300.570 829.505 304.790 830.010 ;
        RECT 305.630 829.505 309.390 830.010 ;
        RECT 310.230 829.505 313.990 830.010 ;
        RECT 314.830 829.505 318.590 830.010 ;
        RECT 319.430 829.505 323.650 830.010 ;
        RECT 324.490 829.505 328.250 830.010 ;
        RECT 329.090 829.505 332.850 830.010 ;
        RECT 333.690 829.505 337.450 830.010 ;
        RECT 338.290 829.505 342.510 830.010 ;
        RECT 343.350 829.505 347.110 830.010 ;
        RECT 347.950 829.505 351.710 830.010 ;
        RECT 352.550 829.505 356.770 830.010 ;
        RECT 357.610 829.505 361.370 830.010 ;
        RECT 362.210 829.505 365.970 830.010 ;
        RECT 366.810 829.505 370.570 830.010 ;
        RECT 371.410 829.505 375.630 830.010 ;
        RECT 376.470 829.505 380.230 830.010 ;
        RECT 381.070 829.505 384.830 830.010 ;
        RECT 385.670 829.505 389.890 830.010 ;
        RECT 390.730 829.505 394.490 830.010 ;
        RECT 395.330 829.505 399.090 830.010 ;
        RECT 399.930 829.505 403.690 830.010 ;
        RECT 404.530 829.505 408.750 830.010 ;
        RECT 409.590 829.505 413.350 830.010 ;
        RECT 414.190 829.505 417.950 830.010 ;
        RECT 418.790 829.505 423.010 830.010 ;
        RECT 423.850 829.505 427.610 830.010 ;
        RECT 428.450 829.505 432.210 830.010 ;
        RECT 433.050 829.505 436.810 830.010 ;
        RECT 437.650 829.505 441.870 830.010 ;
        RECT 442.710 829.505 446.470 830.010 ;
        RECT 447.310 829.505 451.070 830.010 ;
        RECT 451.910 829.505 456.130 830.010 ;
        RECT 456.970 829.505 460.730 830.010 ;
        RECT 461.570 829.505 465.330 830.010 ;
        RECT 466.170 829.505 469.930 830.010 ;
        RECT 470.770 829.505 474.990 830.010 ;
        RECT 475.830 829.505 479.590 830.010 ;
        RECT 480.430 829.505 484.190 830.010 ;
        RECT 485.030 829.505 489.250 830.010 ;
        RECT 490.090 829.505 493.850 830.010 ;
        RECT 494.690 829.505 498.450 830.010 ;
        RECT 499.290 829.505 503.050 830.010 ;
        RECT 503.890 829.505 508.110 830.010 ;
        RECT 508.950 829.505 512.710 830.010 ;
        RECT 513.550 829.505 517.310 830.010 ;
        RECT 518.150 829.505 521.910 830.010 ;
        RECT 522.750 829.505 526.970 830.010 ;
        RECT 527.810 829.505 531.570 830.010 ;
        RECT 532.410 829.505 536.170 830.010 ;
        RECT 537.010 829.505 541.230 830.010 ;
        RECT 542.070 829.505 545.830 830.010 ;
        RECT 546.670 829.505 550.430 830.010 ;
        RECT 551.270 829.505 555.030 830.010 ;
        RECT 555.870 829.505 560.090 830.010 ;
        RECT 560.930 829.505 564.690 830.010 ;
        RECT 565.530 829.505 569.290 830.010 ;
        RECT 570.130 829.505 574.350 830.010 ;
        RECT 575.190 829.505 578.950 830.010 ;
        RECT 579.790 829.505 583.550 830.010 ;
        RECT 584.390 829.505 588.150 830.010 ;
        RECT 588.990 829.505 593.210 830.010 ;
        RECT 594.050 829.505 597.810 830.010 ;
        RECT 598.650 829.505 602.410 830.010 ;
        RECT 603.250 829.505 607.470 830.010 ;
        RECT 608.310 829.505 612.070 830.010 ;
        RECT 612.910 829.505 616.670 830.010 ;
        RECT 617.510 829.505 621.270 830.010 ;
        RECT 622.110 829.505 626.330 830.010 ;
        RECT 627.170 829.505 630.930 830.010 ;
        RECT 631.770 829.505 635.530 830.010 ;
        RECT 636.370 829.505 640.590 830.010 ;
        RECT 641.430 829.505 645.190 830.010 ;
        RECT 646.030 829.505 649.790 830.010 ;
        RECT 650.630 829.505 654.390 830.010 ;
        RECT 655.230 829.505 659.450 830.010 ;
        RECT 660.290 829.505 664.050 830.010 ;
        RECT 664.890 829.505 668.650 830.010 ;
        RECT 669.490 829.505 673.250 830.010 ;
        RECT 674.090 829.505 678.310 830.010 ;
        RECT 679.150 829.505 682.910 830.010 ;
        RECT 683.750 829.505 687.510 830.010 ;
        RECT 688.350 829.505 692.570 830.010 ;
        RECT 693.410 829.505 697.170 830.010 ;
        RECT 698.010 829.505 701.770 830.010 ;
        RECT 702.610 829.505 706.370 830.010 ;
        RECT 707.210 829.505 711.430 830.010 ;
        RECT 712.270 829.505 716.030 830.010 ;
        RECT 716.870 829.505 720.630 830.010 ;
        RECT 721.470 829.505 725.690 830.010 ;
        RECT 726.530 829.505 730.290 830.010 ;
        RECT 731.130 829.505 734.890 830.010 ;
        RECT 735.730 829.505 739.490 830.010 ;
        RECT 740.330 829.505 744.550 830.010 ;
        RECT 745.390 829.505 749.150 830.010 ;
        RECT 749.990 829.505 753.750 830.010 ;
        RECT 754.590 829.505 758.810 830.010 ;
        RECT 759.650 829.505 763.410 830.010 ;
        RECT 764.250 829.505 768.010 830.010 ;
        RECT 768.850 829.505 772.610 830.010 ;
        RECT 773.450 829.505 777.670 830.010 ;
        RECT 778.510 829.505 782.270 830.010 ;
        RECT 783.110 829.505 786.870 830.010 ;
        RECT 787.710 829.505 791.930 830.010 ;
        RECT 792.770 829.505 796.530 830.010 ;
        RECT 797.370 829.505 801.130 830.010 ;
        RECT 801.970 829.505 805.730 830.010 ;
        RECT 806.570 829.505 810.790 830.010 ;
        RECT 811.630 829.505 815.390 830.010 ;
        RECT 816.230 829.505 819.990 830.010 ;
        RECT 820.830 829.505 822.850 830.010 ;
        RECT 0.100 4.280 822.850 829.505 ;
        RECT 0.100 2.875 2.110 4.280 ;
        RECT 2.950 2.875 6.710 4.280 ;
        RECT 7.550 2.875 11.310 4.280 ;
        RECT 12.150 2.875 16.370 4.280 ;
        RECT 17.210 2.875 20.970 4.280 ;
        RECT 21.810 2.875 26.030 4.280 ;
        RECT 26.870 2.875 30.630 4.280 ;
        RECT 31.470 2.875 35.230 4.280 ;
        RECT 36.070 2.875 40.290 4.280 ;
        RECT 41.130 2.875 44.890 4.280 ;
        RECT 45.730 2.875 49.950 4.280 ;
        RECT 50.790 2.875 54.550 4.280 ;
        RECT 55.390 2.875 59.150 4.280 ;
        RECT 59.990 2.875 64.210 4.280 ;
        RECT 65.050 2.875 68.810 4.280 ;
        RECT 69.650 2.875 73.870 4.280 ;
        RECT 74.710 2.875 78.470 4.280 ;
        RECT 79.310 2.875 83.070 4.280 ;
        RECT 83.910 2.875 88.130 4.280 ;
        RECT 88.970 2.875 92.730 4.280 ;
        RECT 93.570 2.875 97.790 4.280 ;
        RECT 98.630 2.875 102.390 4.280 ;
        RECT 103.230 2.875 106.990 4.280 ;
        RECT 107.830 2.875 112.050 4.280 ;
        RECT 112.890 2.875 116.650 4.280 ;
        RECT 117.490 2.875 121.710 4.280 ;
        RECT 122.550 2.875 126.310 4.280 ;
        RECT 127.150 2.875 130.910 4.280 ;
        RECT 131.750 2.875 135.970 4.280 ;
        RECT 136.810 2.875 140.570 4.280 ;
        RECT 141.410 2.875 145.630 4.280 ;
        RECT 146.470 2.875 150.230 4.280 ;
        RECT 151.070 2.875 154.830 4.280 ;
        RECT 155.670 2.875 159.890 4.280 ;
        RECT 160.730 2.875 164.490 4.280 ;
        RECT 165.330 2.875 169.550 4.280 ;
        RECT 170.390 2.875 174.150 4.280 ;
        RECT 174.990 2.875 178.750 4.280 ;
        RECT 179.590 2.875 183.810 4.280 ;
        RECT 184.650 2.875 188.410 4.280 ;
        RECT 189.250 2.875 193.470 4.280 ;
        RECT 194.310 2.875 198.070 4.280 ;
        RECT 198.910 2.875 202.670 4.280 ;
        RECT 203.510 2.875 207.730 4.280 ;
        RECT 208.570 2.875 212.330 4.280 ;
        RECT 213.170 2.875 217.390 4.280 ;
        RECT 218.230 2.875 221.990 4.280 ;
        RECT 222.830 2.875 226.590 4.280 ;
        RECT 227.430 2.875 231.650 4.280 ;
        RECT 232.490 2.875 236.250 4.280 ;
        RECT 237.090 2.875 241.310 4.280 ;
        RECT 242.150 2.875 245.910 4.280 ;
        RECT 246.750 2.875 250.510 4.280 ;
        RECT 251.350 2.875 255.570 4.280 ;
        RECT 256.410 2.875 260.170 4.280 ;
        RECT 261.010 2.875 265.230 4.280 ;
        RECT 266.070 2.875 269.830 4.280 ;
        RECT 270.670 2.875 274.430 4.280 ;
        RECT 275.270 2.875 279.490 4.280 ;
        RECT 280.330 2.875 284.090 4.280 ;
        RECT 284.930 2.875 289.150 4.280 ;
        RECT 289.990 2.875 293.750 4.280 ;
        RECT 294.590 2.875 298.350 4.280 ;
        RECT 299.190 2.875 303.410 4.280 ;
        RECT 304.250 2.875 308.010 4.280 ;
        RECT 308.850 2.875 313.070 4.280 ;
        RECT 313.910 2.875 317.670 4.280 ;
        RECT 318.510 2.875 322.270 4.280 ;
        RECT 323.110 2.875 327.330 4.280 ;
        RECT 328.170 2.875 331.930 4.280 ;
        RECT 332.770 2.875 336.990 4.280 ;
        RECT 337.830 2.875 341.590 4.280 ;
        RECT 342.430 2.875 346.190 4.280 ;
        RECT 347.030 2.875 351.250 4.280 ;
        RECT 352.090 2.875 355.850 4.280 ;
        RECT 356.690 2.875 360.910 4.280 ;
        RECT 361.750 2.875 365.510 4.280 ;
        RECT 366.350 2.875 370.110 4.280 ;
        RECT 370.950 2.875 375.170 4.280 ;
        RECT 376.010 2.875 379.770 4.280 ;
        RECT 380.610 2.875 384.830 4.280 ;
        RECT 385.670 2.875 389.430 4.280 ;
        RECT 390.270 2.875 394.030 4.280 ;
        RECT 394.870 2.875 399.090 4.280 ;
        RECT 399.930 2.875 403.690 4.280 ;
        RECT 404.530 2.875 408.750 4.280 ;
        RECT 409.590 2.875 413.350 4.280 ;
        RECT 414.190 2.875 417.950 4.280 ;
        RECT 418.790 2.875 423.010 4.280 ;
        RECT 423.850 2.875 427.610 4.280 ;
        RECT 428.450 2.875 432.670 4.280 ;
        RECT 433.510 2.875 437.270 4.280 ;
        RECT 438.110 2.875 441.870 4.280 ;
        RECT 442.710 2.875 446.930 4.280 ;
        RECT 447.770 2.875 451.530 4.280 ;
        RECT 452.370 2.875 456.590 4.280 ;
        RECT 457.430 2.875 461.190 4.280 ;
        RECT 462.030 2.875 465.790 4.280 ;
        RECT 466.630 2.875 470.850 4.280 ;
        RECT 471.690 2.875 475.450 4.280 ;
        RECT 476.290 2.875 480.510 4.280 ;
        RECT 481.350 2.875 485.110 4.280 ;
        RECT 485.950 2.875 489.710 4.280 ;
        RECT 490.550 2.875 494.770 4.280 ;
        RECT 495.610 2.875 499.370 4.280 ;
        RECT 500.210 2.875 504.430 4.280 ;
        RECT 505.270 2.875 509.030 4.280 ;
        RECT 509.870 2.875 513.630 4.280 ;
        RECT 514.470 2.875 518.690 4.280 ;
        RECT 519.530 2.875 523.290 4.280 ;
        RECT 524.130 2.875 528.350 4.280 ;
        RECT 529.190 2.875 532.950 4.280 ;
        RECT 533.790 2.875 537.550 4.280 ;
        RECT 538.390 2.875 542.610 4.280 ;
        RECT 543.450 2.875 547.210 4.280 ;
        RECT 548.050 2.875 552.270 4.280 ;
        RECT 553.110 2.875 556.870 4.280 ;
        RECT 557.710 2.875 561.470 4.280 ;
        RECT 562.310 2.875 566.530 4.280 ;
        RECT 567.370 2.875 571.130 4.280 ;
        RECT 571.970 2.875 576.190 4.280 ;
        RECT 577.030 2.875 580.790 4.280 ;
        RECT 581.630 2.875 585.390 4.280 ;
        RECT 586.230 2.875 590.450 4.280 ;
        RECT 591.290 2.875 595.050 4.280 ;
        RECT 595.890 2.875 600.110 4.280 ;
        RECT 600.950 2.875 604.710 4.280 ;
        RECT 605.550 2.875 609.310 4.280 ;
        RECT 610.150 2.875 614.370 4.280 ;
        RECT 615.210 2.875 618.970 4.280 ;
        RECT 619.810 2.875 624.030 4.280 ;
        RECT 624.870 2.875 628.630 4.280 ;
        RECT 629.470 2.875 633.230 4.280 ;
        RECT 634.070 2.875 638.290 4.280 ;
        RECT 639.130 2.875 642.890 4.280 ;
        RECT 643.730 2.875 647.950 4.280 ;
        RECT 648.790 2.875 652.550 4.280 ;
        RECT 653.390 2.875 657.150 4.280 ;
        RECT 657.990 2.875 662.210 4.280 ;
        RECT 663.050 2.875 666.810 4.280 ;
        RECT 667.650 2.875 671.870 4.280 ;
        RECT 672.710 2.875 676.470 4.280 ;
        RECT 677.310 2.875 681.070 4.280 ;
        RECT 681.910 2.875 686.130 4.280 ;
        RECT 686.970 2.875 690.730 4.280 ;
        RECT 691.570 2.875 695.790 4.280 ;
        RECT 696.630 2.875 700.390 4.280 ;
        RECT 701.230 2.875 704.990 4.280 ;
        RECT 705.830 2.875 710.050 4.280 ;
        RECT 710.890 2.875 714.650 4.280 ;
        RECT 715.490 2.875 719.710 4.280 ;
        RECT 720.550 2.875 724.310 4.280 ;
        RECT 725.150 2.875 728.910 4.280 ;
        RECT 729.750 2.875 733.970 4.280 ;
        RECT 734.810 2.875 738.570 4.280 ;
        RECT 739.410 2.875 743.630 4.280 ;
        RECT 744.470 2.875 748.230 4.280 ;
        RECT 749.070 2.875 752.830 4.280 ;
        RECT 753.670 2.875 757.890 4.280 ;
        RECT 758.730 2.875 762.490 4.280 ;
        RECT 763.330 2.875 767.550 4.280 ;
        RECT 768.390 2.875 772.150 4.280 ;
        RECT 772.990 2.875 776.750 4.280 ;
        RECT 777.590 2.875 781.810 4.280 ;
        RECT 782.650 2.875 786.410 4.280 ;
        RECT 787.250 2.875 791.470 4.280 ;
        RECT 792.310 2.875 796.070 4.280 ;
        RECT 796.910 2.875 800.670 4.280 ;
        RECT 801.510 2.875 805.730 4.280 ;
        RECT 806.570 2.875 810.330 4.280 ;
        RECT 811.170 2.875 815.390 4.280 ;
        RECT 816.230 2.875 819.990 4.280 ;
        RECT 820.830 2.875 822.850 4.280 ;
      LAYER met3 ;
        RECT 4.000 826.560 818.665 826.705 ;
        RECT 4.400 825.840 818.665 826.560 ;
        RECT 4.400 825.160 822.900 825.840 ;
        RECT 4.000 814.320 822.900 825.160 ;
        RECT 4.000 812.920 818.665 814.320 ;
        RECT 4.000 811.600 822.900 812.920 ;
        RECT 4.400 810.200 822.900 811.600 ;
        RECT 4.000 801.400 822.900 810.200 ;
        RECT 4.000 800.000 818.665 801.400 ;
        RECT 4.000 796.640 822.900 800.000 ;
        RECT 4.400 795.240 822.900 796.640 ;
        RECT 4.000 788.480 822.900 795.240 ;
        RECT 4.000 787.080 818.665 788.480 ;
        RECT 4.000 781.000 822.900 787.080 ;
        RECT 4.400 779.600 822.900 781.000 ;
        RECT 4.000 775.560 822.900 779.600 ;
        RECT 4.000 774.160 818.665 775.560 ;
        RECT 4.000 766.040 822.900 774.160 ;
        RECT 4.400 764.640 822.900 766.040 ;
        RECT 4.000 762.640 822.900 764.640 ;
        RECT 4.000 761.240 818.665 762.640 ;
        RECT 4.000 751.080 822.900 761.240 ;
        RECT 4.400 749.680 822.900 751.080 ;
        RECT 4.000 749.040 822.900 749.680 ;
        RECT 4.000 747.640 818.665 749.040 ;
        RECT 4.000 736.120 822.900 747.640 ;
        RECT 4.000 735.440 818.665 736.120 ;
        RECT 4.400 734.720 818.665 735.440 ;
        RECT 4.400 734.040 822.900 734.720 ;
        RECT 4.000 723.200 822.900 734.040 ;
        RECT 4.000 721.800 818.665 723.200 ;
        RECT 4.000 720.480 822.900 721.800 ;
        RECT 4.400 719.080 822.900 720.480 ;
        RECT 4.000 710.280 822.900 719.080 ;
        RECT 4.000 708.880 818.665 710.280 ;
        RECT 4.000 705.520 822.900 708.880 ;
        RECT 4.400 704.120 822.900 705.520 ;
        RECT 4.000 697.360 822.900 704.120 ;
        RECT 4.000 695.960 818.665 697.360 ;
        RECT 4.000 690.560 822.900 695.960 ;
        RECT 4.400 689.160 822.900 690.560 ;
        RECT 4.000 684.440 822.900 689.160 ;
        RECT 4.000 683.040 818.665 684.440 ;
        RECT 4.000 674.920 822.900 683.040 ;
        RECT 4.400 673.520 822.900 674.920 ;
        RECT 4.000 670.840 822.900 673.520 ;
        RECT 4.000 669.440 818.665 670.840 ;
        RECT 4.000 659.960 822.900 669.440 ;
        RECT 4.400 658.560 822.900 659.960 ;
        RECT 4.000 657.920 822.900 658.560 ;
        RECT 4.000 656.520 818.665 657.920 ;
        RECT 4.000 645.000 822.900 656.520 ;
        RECT 4.400 643.600 818.665 645.000 ;
        RECT 4.000 632.080 822.900 643.600 ;
        RECT 4.000 630.680 818.665 632.080 ;
        RECT 4.000 629.360 822.900 630.680 ;
        RECT 4.400 627.960 822.900 629.360 ;
        RECT 4.000 619.160 822.900 627.960 ;
        RECT 4.000 617.760 818.665 619.160 ;
        RECT 4.000 614.400 822.900 617.760 ;
        RECT 4.400 613.000 822.900 614.400 ;
        RECT 4.000 606.240 822.900 613.000 ;
        RECT 4.000 604.840 818.665 606.240 ;
        RECT 4.000 599.440 822.900 604.840 ;
        RECT 4.400 598.040 822.900 599.440 ;
        RECT 4.000 593.320 822.900 598.040 ;
        RECT 4.000 591.920 818.665 593.320 ;
        RECT 4.000 584.480 822.900 591.920 ;
        RECT 4.400 583.080 822.900 584.480 ;
        RECT 4.000 579.720 822.900 583.080 ;
        RECT 4.000 578.320 818.665 579.720 ;
        RECT 4.000 568.840 822.900 578.320 ;
        RECT 4.400 567.440 822.900 568.840 ;
        RECT 4.000 566.800 822.900 567.440 ;
        RECT 4.000 565.400 818.665 566.800 ;
        RECT 4.000 553.880 822.900 565.400 ;
        RECT 4.400 552.480 818.665 553.880 ;
        RECT 4.000 540.960 822.900 552.480 ;
        RECT 4.000 539.560 818.665 540.960 ;
        RECT 4.000 538.920 822.900 539.560 ;
        RECT 4.400 537.520 822.900 538.920 ;
        RECT 4.000 528.040 822.900 537.520 ;
        RECT 4.000 526.640 818.665 528.040 ;
        RECT 4.000 523.280 822.900 526.640 ;
        RECT 4.400 521.880 822.900 523.280 ;
        RECT 4.000 515.120 822.900 521.880 ;
        RECT 4.000 513.720 818.665 515.120 ;
        RECT 4.000 508.320 822.900 513.720 ;
        RECT 4.400 506.920 822.900 508.320 ;
        RECT 4.000 501.520 822.900 506.920 ;
        RECT 4.000 500.120 818.665 501.520 ;
        RECT 4.000 493.360 822.900 500.120 ;
        RECT 4.400 491.960 822.900 493.360 ;
        RECT 4.000 488.600 822.900 491.960 ;
        RECT 4.000 487.200 818.665 488.600 ;
        RECT 4.000 478.400 822.900 487.200 ;
        RECT 4.400 477.000 822.900 478.400 ;
        RECT 4.000 475.680 822.900 477.000 ;
        RECT 4.000 474.280 818.665 475.680 ;
        RECT 4.000 462.760 822.900 474.280 ;
        RECT 4.400 461.360 818.665 462.760 ;
        RECT 4.000 449.840 822.900 461.360 ;
        RECT 4.000 448.440 818.665 449.840 ;
        RECT 4.000 447.800 822.900 448.440 ;
        RECT 4.400 446.400 822.900 447.800 ;
        RECT 4.000 436.920 822.900 446.400 ;
        RECT 4.000 435.520 818.665 436.920 ;
        RECT 4.000 432.840 822.900 435.520 ;
        RECT 4.400 431.440 822.900 432.840 ;
        RECT 4.000 424.000 822.900 431.440 ;
        RECT 4.000 422.600 818.665 424.000 ;
        RECT 4.000 417.200 822.900 422.600 ;
        RECT 4.400 415.800 822.900 417.200 ;
        RECT 4.000 410.400 822.900 415.800 ;
        RECT 4.000 409.000 818.665 410.400 ;
        RECT 4.000 402.240 822.900 409.000 ;
        RECT 4.400 400.840 822.900 402.240 ;
        RECT 4.000 397.480 822.900 400.840 ;
        RECT 4.000 396.080 818.665 397.480 ;
        RECT 4.000 387.280 822.900 396.080 ;
        RECT 4.400 385.880 822.900 387.280 ;
        RECT 4.000 384.560 822.900 385.880 ;
        RECT 4.000 383.160 818.665 384.560 ;
        RECT 4.000 371.640 822.900 383.160 ;
        RECT 4.400 370.240 818.665 371.640 ;
        RECT 4.000 358.720 822.900 370.240 ;
        RECT 4.000 357.320 818.665 358.720 ;
        RECT 4.000 356.680 822.900 357.320 ;
        RECT 4.400 355.280 822.900 356.680 ;
        RECT 4.000 345.800 822.900 355.280 ;
        RECT 4.000 344.400 818.665 345.800 ;
        RECT 4.000 341.720 822.900 344.400 ;
        RECT 4.400 340.320 822.900 341.720 ;
        RECT 4.000 332.200 822.900 340.320 ;
        RECT 4.000 330.800 818.665 332.200 ;
        RECT 4.000 326.760 822.900 330.800 ;
        RECT 4.400 325.360 822.900 326.760 ;
        RECT 4.000 319.280 822.900 325.360 ;
        RECT 4.000 317.880 818.665 319.280 ;
        RECT 4.000 311.120 822.900 317.880 ;
        RECT 4.400 309.720 822.900 311.120 ;
        RECT 4.000 306.360 822.900 309.720 ;
        RECT 4.000 304.960 818.665 306.360 ;
        RECT 4.000 296.160 822.900 304.960 ;
        RECT 4.400 294.760 822.900 296.160 ;
        RECT 4.000 293.440 822.900 294.760 ;
        RECT 4.000 292.040 818.665 293.440 ;
        RECT 4.000 281.200 822.900 292.040 ;
        RECT 4.400 280.520 822.900 281.200 ;
        RECT 4.400 279.800 818.665 280.520 ;
        RECT 4.000 279.120 818.665 279.800 ;
        RECT 4.000 267.600 822.900 279.120 ;
        RECT 4.000 266.200 818.665 267.600 ;
        RECT 4.000 265.560 822.900 266.200 ;
        RECT 4.400 264.160 822.900 265.560 ;
        RECT 4.000 254.000 822.900 264.160 ;
        RECT 4.000 252.600 818.665 254.000 ;
        RECT 4.000 250.600 822.900 252.600 ;
        RECT 4.400 249.200 822.900 250.600 ;
        RECT 4.000 241.080 822.900 249.200 ;
        RECT 4.000 239.680 818.665 241.080 ;
        RECT 4.000 235.640 822.900 239.680 ;
        RECT 4.400 234.240 822.900 235.640 ;
        RECT 4.000 228.160 822.900 234.240 ;
        RECT 4.000 226.760 818.665 228.160 ;
        RECT 4.000 220.680 822.900 226.760 ;
        RECT 4.400 219.280 822.900 220.680 ;
        RECT 4.000 215.240 822.900 219.280 ;
        RECT 4.000 213.840 818.665 215.240 ;
        RECT 4.000 205.040 822.900 213.840 ;
        RECT 4.400 203.640 822.900 205.040 ;
        RECT 4.000 202.320 822.900 203.640 ;
        RECT 4.000 200.920 818.665 202.320 ;
        RECT 4.000 190.080 822.900 200.920 ;
        RECT 4.400 189.400 822.900 190.080 ;
        RECT 4.400 188.680 818.665 189.400 ;
        RECT 4.000 188.000 818.665 188.680 ;
        RECT 4.000 176.480 822.900 188.000 ;
        RECT 4.000 175.120 818.665 176.480 ;
        RECT 4.400 175.080 818.665 175.120 ;
        RECT 4.400 173.720 822.900 175.080 ;
        RECT 4.000 162.880 822.900 173.720 ;
        RECT 4.000 161.480 818.665 162.880 ;
        RECT 4.000 159.480 822.900 161.480 ;
        RECT 4.400 158.080 822.900 159.480 ;
        RECT 4.000 149.960 822.900 158.080 ;
        RECT 4.000 148.560 818.665 149.960 ;
        RECT 4.000 144.520 822.900 148.560 ;
        RECT 4.400 143.120 822.900 144.520 ;
        RECT 4.000 137.040 822.900 143.120 ;
        RECT 4.000 135.640 818.665 137.040 ;
        RECT 4.000 129.560 822.900 135.640 ;
        RECT 4.400 128.160 822.900 129.560 ;
        RECT 4.000 124.120 822.900 128.160 ;
        RECT 4.000 122.720 818.665 124.120 ;
        RECT 4.000 114.600 822.900 122.720 ;
        RECT 4.400 113.200 822.900 114.600 ;
        RECT 4.000 111.200 822.900 113.200 ;
        RECT 4.000 109.800 818.665 111.200 ;
        RECT 4.000 98.960 822.900 109.800 ;
        RECT 4.400 98.280 822.900 98.960 ;
        RECT 4.400 97.560 818.665 98.280 ;
        RECT 4.000 96.880 818.665 97.560 ;
        RECT 4.000 84.680 822.900 96.880 ;
        RECT 4.000 84.000 818.665 84.680 ;
        RECT 4.400 83.280 818.665 84.000 ;
        RECT 4.400 82.600 822.900 83.280 ;
        RECT 4.000 71.760 822.900 82.600 ;
        RECT 4.000 70.360 818.665 71.760 ;
        RECT 4.000 69.040 822.900 70.360 ;
        RECT 4.400 67.640 822.900 69.040 ;
        RECT 4.000 58.840 822.900 67.640 ;
        RECT 4.000 57.440 818.665 58.840 ;
        RECT 4.000 53.400 822.900 57.440 ;
        RECT 4.400 52.000 822.900 53.400 ;
        RECT 4.000 45.920 822.900 52.000 ;
        RECT 4.000 44.520 818.665 45.920 ;
        RECT 4.000 38.440 822.900 44.520 ;
        RECT 4.400 37.040 822.900 38.440 ;
        RECT 4.000 33.000 822.900 37.040 ;
        RECT 4.000 31.600 818.665 33.000 ;
        RECT 4.000 23.480 822.900 31.600 ;
        RECT 4.400 22.080 822.900 23.480 ;
        RECT 4.000 20.080 822.900 22.080 ;
        RECT 4.000 18.680 818.665 20.080 ;
        RECT 4.000 8.520 822.900 18.680 ;
        RECT 4.400 7.160 822.900 8.520 ;
        RECT 4.400 7.120 818.665 7.160 ;
        RECT 4.000 5.760 818.665 7.120 ;
        RECT 4.000 2.895 822.900 5.760 ;
      LAYER met4 ;
        RECT 92.295 10.240 97.440 819.905 ;
        RECT 99.840 10.240 174.240 819.905 ;
        RECT 176.640 10.240 251.040 819.905 ;
        RECT 253.440 10.240 327.840 819.905 ;
        RECT 330.240 10.240 404.640 819.905 ;
        RECT 407.040 10.240 481.440 819.905 ;
        RECT 483.840 10.240 558.240 819.905 ;
        RECT 560.640 10.240 635.040 819.905 ;
        RECT 637.440 10.240 711.840 819.905 ;
        RECT 714.240 10.240 788.640 819.905 ;
        RECT 791.040 318.050 823.065 819.905 ;
        RECT 791.040 259.270 823.090 318.050 ;
        RECT 791.040 10.240 823.065 259.270 ;
        RECT 92.295 2.895 823.065 10.240 ;
  END
END user_proj
END LIBRARY

