magic
tech sky130A
magscale 1 2
timestamp 1640322195
<< metal1 >>
rect 201494 702992 201500 703044
rect 201552 703032 201558 703044
rect 202782 703032 202788 703044
rect 201552 703004 202788 703032
rect 201552 702992 201558 703004
rect 202782 702992 202788 703004
rect 202840 702992 202846 703044
rect 209130 700816 209136 700868
rect 209188 700856 209194 700868
rect 218974 700856 218980 700868
rect 209188 700828 218980 700856
rect 209188 700816 209194 700828
rect 218974 700816 218980 700828
rect 219032 700816 219038 700868
rect 197998 700748 198004 700800
rect 198056 700788 198062 700800
rect 235166 700788 235172 700800
rect 198056 700760 235172 700788
rect 198056 700748 198062 700760
rect 235166 700748 235172 700760
rect 235224 700748 235230 700800
rect 206278 700680 206284 700732
rect 206336 700720 206342 700732
rect 267642 700720 267648 700732
rect 206336 700692 267648 700720
rect 206336 700680 206342 700692
rect 267642 700680 267648 700692
rect 267700 700680 267706 700732
rect 200758 700612 200764 700664
rect 200816 700652 200822 700664
rect 283834 700652 283840 700664
rect 200816 700624 283840 700652
rect 200816 700612 200822 700624
rect 283834 700612 283840 700624
rect 283892 700612 283898 700664
rect 204898 700544 204904 700596
rect 204956 700584 204962 700596
rect 300118 700584 300124 700596
rect 204956 700556 300124 700584
rect 204956 700544 204962 700556
rect 300118 700544 300124 700556
rect 300176 700544 300182 700596
rect 385678 700544 385684 700596
rect 385736 700584 385742 700596
rect 462314 700584 462320 700596
rect 385736 700556 462320 700584
rect 385736 700544 385742 700556
rect 462314 700544 462320 700556
rect 462372 700544 462378 700596
rect 213178 700476 213184 700528
rect 213236 700516 213242 700528
rect 332502 700516 332508 700528
rect 213236 700488 332508 700516
rect 213236 700476 213242 700488
rect 332502 700476 332508 700488
rect 332560 700476 332566 700528
rect 388438 700476 388444 700528
rect 388496 700516 388502 700528
rect 397454 700516 397460 700528
rect 388496 700488 397460 700516
rect 388496 700476 388502 700488
rect 397454 700476 397460 700488
rect 397512 700476 397518 700528
rect 400858 700476 400864 700528
rect 400916 700516 400922 700528
rect 478506 700516 478512 700528
rect 400916 700488 478512 700516
rect 400916 700476 400922 700488
rect 478506 700476 478512 700488
rect 478564 700476 478570 700528
rect 215938 700408 215944 700460
rect 215996 700448 216002 700460
rect 348786 700448 348792 700460
rect 215996 700420 348792 700448
rect 215996 700408 216002 700420
rect 348786 700408 348792 700420
rect 348844 700408 348850 700460
rect 370498 700408 370504 700460
rect 370556 700448 370562 700460
rect 494790 700448 494796 700460
rect 370556 700420 494796 700448
rect 370556 700408 370562 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 40494 700340 40500 700392
rect 40552 700380 40558 700392
rect 41322 700380 41328 700392
rect 40552 700352 41328 700380
rect 40552 700340 40558 700352
rect 41322 700340 41328 700352
rect 41380 700340 41386 700392
rect 170306 700340 170312 700392
rect 170364 700380 170370 700392
rect 196526 700380 196532 700392
rect 170364 700352 196532 700380
rect 170364 700340 170370 700352
rect 196526 700340 196532 700352
rect 196584 700340 196590 700392
rect 214558 700340 214564 700392
rect 214616 700380 214622 700392
rect 364978 700380 364984 700392
rect 214616 700352 364984 700380
rect 214616 700340 214622 700352
rect 364978 700340 364984 700352
rect 365036 700340 365042 700392
rect 382918 700340 382924 700392
rect 382976 700380 382982 700392
rect 527174 700380 527180 700392
rect 382976 700352 527180 700380
rect 382976 700340 382982 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 33778 700312 33784 700324
rect 24360 700284 33784 700312
rect 24360 700272 24366 700284
rect 33778 700272 33784 700284
rect 33836 700272 33842 700324
rect 58802 700272 58808 700324
rect 58860 700312 58866 700324
rect 72970 700312 72976 700324
rect 58860 700284 72976 700312
rect 58860 700272 58866 700284
rect 72970 700272 72976 700284
rect 73028 700272 73034 700324
rect 137830 700272 137836 700324
rect 137888 700312 137894 700324
rect 146938 700312 146944 700324
rect 137888 700284 146944 700312
rect 137888 700272 137894 700284
rect 146938 700272 146944 700284
rect 146996 700272 147002 700324
rect 154114 700272 154120 700324
rect 154172 700312 154178 700324
rect 196618 700312 196624 700324
rect 154172 700284 196624 700312
rect 154172 700272 154178 700284
rect 196618 700272 196624 700284
rect 196676 700272 196682 700324
rect 209038 700272 209044 700324
rect 209096 700312 209102 700324
rect 559650 700312 559656 700324
rect 209096 700284 559656 700312
rect 209096 700272 209102 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 88334 699660 88340 699712
rect 88392 699700 88398 699712
rect 89162 699700 89168 699712
rect 88392 699672 89168 699700
rect 88392 699660 88398 699672
rect 89162 699660 89168 699672
rect 89220 699660 89226 699712
rect 104894 699660 104900 699712
rect 104952 699700 104958 699712
rect 105446 699700 105452 699712
rect 104952 699672 105452 699700
rect 104952 699660 104958 699672
rect 105446 699660 105452 699672
rect 105504 699660 105510 699712
rect 381538 696940 381544 696992
rect 381596 696980 381602 696992
rect 580166 696980 580172 696992
rect 381596 696952 580172 696980
rect 381596 696940 381602 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 2774 683680 2780 683732
rect 2832 683720 2838 683732
rect 4798 683720 4804 683732
rect 2832 683692 4804 683720
rect 2832 683680 2838 683692
rect 4798 683680 4804 683692
rect 4856 683680 4862 683732
rect 399478 683136 399484 683188
rect 399536 683176 399542 683188
rect 580166 683176 580172 683188
rect 399536 683148 580172 683176
rect 399536 683136 399542 683148
rect 580166 683136 580172 683148
rect 580224 683136 580230 683188
rect 146938 677492 146944 677544
rect 146996 677532 147002 677544
rect 153838 677532 153844 677544
rect 146996 677504 153844 677532
rect 146996 677492 147002 677504
rect 153838 677492 153844 677504
rect 153896 677492 153902 677544
rect 3510 670692 3516 670744
rect 3568 670732 3574 670744
rect 35158 670732 35164 670744
rect 3568 670704 35164 670732
rect 3568 670692 3574 670704
rect 35158 670692 35164 670704
rect 35216 670692 35222 670744
rect 206370 670692 206376 670744
rect 206428 670732 206434 670744
rect 580166 670732 580172 670744
rect 206428 670704 580172 670732
rect 206428 670692 206434 670704
rect 580166 670692 580172 670704
rect 580224 670692 580230 670744
rect 153838 661036 153844 661088
rect 153896 661076 153902 661088
rect 159358 661076 159364 661088
rect 153896 661048 159364 661076
rect 153896 661036 153902 661048
rect 159358 661036 159364 661048
rect 159416 661036 159422 661088
rect 3418 656888 3424 656940
rect 3476 656928 3482 656940
rect 15838 656928 15844 656940
rect 3476 656900 15844 656928
rect 3476 656888 3482 656900
rect 15838 656888 15844 656900
rect 15896 656888 15902 656940
rect 159358 652672 159364 652724
rect 159416 652712 159422 652724
rect 162762 652712 162768 652724
rect 159416 652684 162768 652712
rect 159416 652672 159422 652684
rect 162762 652672 162768 652684
rect 162820 652672 162826 652724
rect 162762 648864 162768 648916
rect 162820 648904 162826 648916
rect 166258 648904 166264 648916
rect 162820 648876 166264 648904
rect 162820 648864 162826 648876
rect 166258 648864 166264 648876
rect 166316 648864 166322 648916
rect 377398 643084 377404 643136
rect 377456 643124 377462 643136
rect 580166 643124 580172 643136
rect 377456 643096 580172 643124
rect 377456 643084 377462 643096
rect 580166 643084 580172 643096
rect 580224 643084 580230 643136
rect 166258 639548 166264 639600
rect 166316 639588 166322 639600
rect 175918 639588 175924 639600
rect 166316 639560 175924 639588
rect 166316 639548 166322 639560
rect 175918 639548 175924 639560
rect 175976 639548 175982 639600
rect 3418 632068 3424 632120
rect 3476 632108 3482 632120
rect 14458 632108 14464 632120
rect 3476 632080 14464 632108
rect 3476 632068 3482 632080
rect 14458 632068 14464 632080
rect 14516 632068 14522 632120
rect 396718 630640 396724 630692
rect 396776 630680 396782 630692
rect 580166 630680 580172 630692
rect 396776 630652 580172 630680
rect 396776 630640 396782 630652
rect 580166 630640 580172 630652
rect 580224 630640 580230 630692
rect 3142 618264 3148 618316
rect 3200 618304 3206 618316
rect 36538 618304 36544 618316
rect 3200 618276 36544 618304
rect 3200 618264 3206 618276
rect 36538 618264 36544 618276
rect 36596 618264 36602 618316
rect 175918 617516 175924 617568
rect 175976 617556 175982 617568
rect 186958 617556 186964 617568
rect 175976 617528 186964 617556
rect 175976 617516 175982 617528
rect 186958 617516 186964 617528
rect 187016 617516 187022 617568
rect 367738 616836 367744 616888
rect 367796 616876 367802 616888
rect 580166 616876 580172 616888
rect 367796 616848 580172 616876
rect 367796 616836 367802 616848
rect 580166 616836 580172 616848
rect 580224 616836 580230 616888
rect 3234 605820 3240 605872
rect 3292 605860 3298 605872
rect 22738 605860 22744 605872
rect 3292 605832 22744 605860
rect 3292 605820 3298 605832
rect 22738 605820 22744 605832
rect 22796 605820 22802 605872
rect 186958 597456 186964 597508
rect 187016 597496 187022 597508
rect 189718 597496 189724 597508
rect 187016 597468 189724 597496
rect 187016 597456 187022 597468
rect 189718 597456 189724 597468
rect 189776 597456 189782 597508
rect 376018 590656 376024 590708
rect 376076 590696 376082 590708
rect 579798 590696 579804 590708
rect 376076 590668 579804 590696
rect 376076 590656 376082 590668
rect 579798 590656 579804 590668
rect 579856 590656 579862 590708
rect 3326 579640 3332 579692
rect 3384 579680 3390 579692
rect 11698 579680 11704 579692
rect 3384 579652 11704 579680
rect 3384 579640 3390 579652
rect 11698 579640 11704 579652
rect 11756 579640 11762 579692
rect 395338 576852 395344 576904
rect 395396 576892 395402 576904
rect 580166 576892 580172 576904
rect 395396 576864 580172 576892
rect 395396 576852 395402 576864
rect 580166 576852 580172 576864
rect 580224 576852 580230 576904
rect 189718 566448 189724 566500
rect 189776 566488 189782 566500
rect 196894 566488 196900 566500
rect 189776 566460 196900 566488
rect 189776 566448 189782 566460
rect 196894 566448 196900 566460
rect 196952 566448 196958 566500
rect 3418 565836 3424 565888
rect 3476 565876 3482 565888
rect 39298 565876 39304 565888
rect 3476 565848 39304 565876
rect 3476 565836 3482 565848
rect 39298 565836 39304 565848
rect 39356 565836 39362 565888
rect 363598 563048 363604 563100
rect 363656 563088 363662 563100
rect 579798 563088 579804 563100
rect 363656 563060 579804 563088
rect 363656 563048 363662 563060
rect 579798 563048 579804 563060
rect 579856 563048 579862 563100
rect 3418 553392 3424 553444
rect 3476 553432 3482 553444
rect 25498 553432 25504 553444
rect 3476 553404 25504 553432
rect 3476 553392 3482 553404
rect 25498 553392 25504 553404
rect 25556 553392 25562 553444
rect 378778 536800 378784 536852
rect 378836 536840 378842 536852
rect 580166 536840 580172 536852
rect 378836 536812 580172 536840
rect 378836 536800 378842 536812
rect 580166 536800 580172 536812
rect 580224 536800 580230 536852
rect 3418 527144 3424 527196
rect 3476 527184 3482 527196
rect 17218 527184 17224 527196
rect 3476 527156 17224 527184
rect 3476 527144 3482 527156
rect 17218 527144 17224 527156
rect 17276 527144 17282 527196
rect 393958 524424 393964 524476
rect 394016 524464 394022 524476
rect 580166 524464 580172 524476
rect 394016 524436 580172 524464
rect 394016 524424 394022 524436
rect 580166 524424 580172 524436
rect 580224 524424 580230 524476
rect 3418 514768 3424 514820
rect 3476 514808 3482 514820
rect 43438 514808 43444 514820
rect 3476 514780 43444 514808
rect 3476 514768 3482 514780
rect 43438 514768 43444 514780
rect 43496 514768 43502 514820
rect 360838 510620 360844 510672
rect 360896 510660 360902 510672
rect 580166 510660 580172 510672
rect 360896 510632 580172 510660
rect 360896 510620 360902 510632
rect 580166 510620 580172 510632
rect 580224 510620 580230 510672
rect 3050 500964 3056 501016
rect 3108 501004 3114 501016
rect 29638 501004 29644 501016
rect 3108 500976 29644 501004
rect 3108 500964 3114 500976
rect 29638 500964 29644 500976
rect 29696 500964 29702 501016
rect 374638 484372 374644 484424
rect 374696 484412 374702 484424
rect 580166 484412 580172 484424
rect 374696 484384 580172 484412
rect 374696 484372 374702 484384
rect 580166 484372 580172 484384
rect 580224 484372 580230 484424
rect 3418 474716 3424 474768
rect 3476 474756 3482 474768
rect 18598 474756 18604 474768
rect 3476 474728 18604 474756
rect 3476 474716 3482 474728
rect 18598 474716 18604 474728
rect 18656 474716 18662 474768
rect 392578 470568 392584 470620
rect 392636 470608 392642 470620
rect 579982 470608 579988 470620
rect 392636 470580 579988 470608
rect 392636 470568 392642 470580
rect 579982 470568 579988 470580
rect 580040 470568 580046 470620
rect 3234 462340 3240 462392
rect 3292 462380 3298 462392
rect 47578 462380 47584 462392
rect 3292 462352 47584 462380
rect 3292 462340 3298 462352
rect 47578 462340 47584 462352
rect 47636 462340 47642 462392
rect 358078 456764 358084 456816
rect 358136 456804 358142 456816
rect 580166 456804 580172 456816
rect 358136 456776 580172 456804
rect 358136 456764 358142 456776
rect 580166 456764 580172 456776
rect 580224 456764 580230 456816
rect 3142 448536 3148 448588
rect 3200 448576 3206 448588
rect 32398 448576 32404 448588
rect 3200 448548 32404 448576
rect 3200 448536 3206 448548
rect 32398 448536 32404 448548
rect 32456 448536 32462 448588
rect 206462 434732 206468 434784
rect 206520 434772 206526 434784
rect 216674 434772 216680 434784
rect 206520 434744 216680 434772
rect 206520 434732 206526 434744
rect 216674 434732 216680 434744
rect 216732 434732 216738 434784
rect 202230 433304 202236 433356
rect 202288 433344 202294 433356
rect 216674 433344 216680 433356
rect 202288 433316 216680 433344
rect 202288 433304 202294 433316
rect 216674 433304 216680 433316
rect 216732 433304 216738 433356
rect 213270 432352 213276 432404
rect 213328 432392 213334 432404
rect 216674 432392 216680 432404
rect 213328 432364 216680 432392
rect 213328 432352 213334 432364
rect 216674 432352 216680 432364
rect 216732 432352 216738 432404
rect 389818 430584 389824 430636
rect 389876 430624 389882 430636
rect 580166 430624 580172 430636
rect 389876 430596 580172 430624
rect 389876 430584 389882 430596
rect 580166 430584 580172 430596
rect 580224 430584 580230 430636
rect 204990 429156 204996 429208
rect 205048 429196 205054 429208
rect 216674 429196 216680 429208
rect 205048 429168 216680 429196
rect 205048 429156 205054 429168
rect 216674 429156 216680 429168
rect 216732 429156 216738 429208
rect 3418 422288 3424 422340
rect 3476 422328 3482 422340
rect 21358 422328 21364 422340
rect 3476 422300 21364 422328
rect 3476 422288 3482 422300
rect 21358 422288 21364 422300
rect 21416 422288 21422 422340
rect 3142 409844 3148 409896
rect 3200 409884 3206 409896
rect 50338 409884 50344 409896
rect 3200 409856 50344 409884
rect 3200 409844 3206 409856
rect 50338 409844 50344 409856
rect 50396 409844 50402 409896
rect 211798 409844 211804 409896
rect 211856 409884 211862 409896
rect 216674 409884 216680 409896
rect 211856 409856 216680 409884
rect 211856 409844 211862 409856
rect 216674 409844 216680 409856
rect 216732 409844 216738 409896
rect 371878 404336 371884 404388
rect 371936 404376 371942 404388
rect 580166 404376 580172 404388
rect 371936 404348 580172 404376
rect 371936 404336 371942 404348
rect 580166 404336 580172 404348
rect 580224 404336 580230 404388
rect 219710 403044 219716 403096
rect 219768 403084 219774 403096
rect 219894 403084 219900 403096
rect 219768 403056 219900 403084
rect 219768 403044 219774 403056
rect 219894 403044 219900 403056
rect 219952 403044 219958 403096
rect 59354 400052 59360 400104
rect 59412 400092 59418 400104
rect 217318 400092 217324 400104
rect 59412 400064 217324 400092
rect 59412 400052 59418 400064
rect 217318 400052 217324 400064
rect 217376 400052 217382 400104
rect 122742 399984 122748 400036
rect 122800 400024 122806 400036
rect 209130 400024 209136 400036
rect 122800 399996 209136 400024
rect 122800 399984 122806 399996
rect 209130 399984 209136 399996
rect 209188 399984 209194 400036
rect 115750 399916 115756 399968
rect 115808 399956 115814 399968
rect 213178 399956 213184 399968
rect 115808 399928 213184 399956
rect 115808 399916 115814 399928
rect 213178 399916 213184 399928
rect 213236 399916 213242 399968
rect 218974 399916 218980 399968
rect 219032 399956 219038 399968
rect 227346 399956 227352 399968
rect 219032 399928 227352 399956
rect 219032 399916 219038 399928
rect 227346 399916 227352 399928
rect 227404 399916 227410 399968
rect 115658 399848 115664 399900
rect 115716 399888 115722 399900
rect 215938 399888 215944 399900
rect 115716 399860 215944 399888
rect 115716 399848 115722 399860
rect 215938 399848 215944 399860
rect 215996 399848 216002 399900
rect 218606 399848 218612 399900
rect 218664 399888 218670 399900
rect 226426 399888 226432 399900
rect 218664 399860 226432 399888
rect 218664 399848 218670 399860
rect 226426 399848 226432 399860
rect 226484 399848 226490 399900
rect 53466 399780 53472 399832
rect 53524 399820 53530 399832
rect 199010 399820 199016 399832
rect 53524 399792 199016 399820
rect 53524 399780 53530 399792
rect 199010 399780 199016 399792
rect 199068 399780 199074 399832
rect 218422 399780 218428 399832
rect 218480 399820 218486 399832
rect 226518 399820 226524 399832
rect 218480 399792 226524 399820
rect 218480 399780 218486 399792
rect 226518 399780 226524 399792
rect 226576 399780 226582 399832
rect 52270 399712 52276 399764
rect 52328 399752 52334 399764
rect 217226 399752 217232 399764
rect 52328 399724 217232 399752
rect 52328 399712 52334 399724
rect 217226 399712 217232 399724
rect 217284 399712 217290 399764
rect 217502 399712 217508 399764
rect 217560 399752 217566 399764
rect 233234 399752 233240 399764
rect 217560 399724 233240 399752
rect 217560 399712 217566 399724
rect 233234 399712 233240 399724
rect 233292 399712 233298 399764
rect 57790 399644 57796 399696
rect 57848 399684 57854 399696
rect 172514 399684 172520 399696
rect 57848 399656 172520 399684
rect 57848 399644 57854 399656
rect 172514 399644 172520 399656
rect 172572 399644 172578 399696
rect 187602 399644 187608 399696
rect 187660 399684 187666 399696
rect 357526 399684 357532 399696
rect 187660 399656 357532 399684
rect 187660 399644 187666 399656
rect 357526 399644 357532 399656
rect 357584 399644 357590 399696
rect 57882 399576 57888 399628
rect 57940 399616 57946 399628
rect 232038 399616 232044 399628
rect 57940 399588 232044 399616
rect 57940 399576 57946 399588
rect 232038 399576 232044 399588
rect 232096 399576 232102 399628
rect 57698 399508 57704 399560
rect 57756 399548 57762 399560
rect 233418 399548 233424 399560
rect 57756 399520 233424 399548
rect 57756 399508 57762 399520
rect 233418 399508 233424 399520
rect 233476 399508 233482 399560
rect 249150 399508 249156 399560
rect 249208 399548 249214 399560
rect 358998 399548 359004 399560
rect 249208 399520 359004 399548
rect 249208 399508 249214 399520
rect 358998 399508 359004 399520
rect 359056 399508 359062 399560
rect 57330 399440 57336 399492
rect 57388 399480 57394 399492
rect 233326 399480 233332 399492
rect 57388 399452 233332 399480
rect 57388 399440 57394 399452
rect 233326 399440 233332 399452
rect 233384 399440 233390 399492
rect 246298 399440 246304 399492
rect 246356 399480 246362 399492
rect 359090 399480 359096 399492
rect 246356 399452 359096 399480
rect 246356 399440 246362 399452
rect 359090 399440 359096 399452
rect 359148 399440 359154 399492
rect 58802 399372 58808 399424
rect 58860 399412 58866 399424
rect 125594 399412 125600 399424
rect 58860 399384 125600 399412
rect 58860 399372 58866 399384
rect 125594 399372 125600 399384
rect 125652 399372 125658 399424
rect 191742 399372 191748 399424
rect 191800 399412 191806 399424
rect 206462 399412 206468 399424
rect 191800 399384 206468 399412
rect 191800 399372 191806 399384
rect 206462 399372 206468 399384
rect 206520 399372 206526 399424
rect 188982 399304 188988 399356
rect 189040 399344 189046 399356
rect 202230 399344 202236 399356
rect 189040 399316 202236 399344
rect 189040 399304 189046 399316
rect 202230 399304 202236 399316
rect 202288 399304 202294 399356
rect 219526 398624 219532 398676
rect 219584 398664 219590 398676
rect 224954 398664 224960 398676
rect 219584 398636 224960 398664
rect 219584 398624 219590 398636
rect 224954 398624 224960 398636
rect 225012 398624 225018 398676
rect 219618 398556 219624 398608
rect 219676 398596 219682 398608
rect 224770 398596 224776 398608
rect 219676 398568 224776 398596
rect 219676 398556 219682 398568
rect 224770 398556 224776 398568
rect 224828 398556 224834 398608
rect 219434 398420 219440 398472
rect 219492 398460 219498 398472
rect 224862 398460 224868 398472
rect 219492 398432 224868 398460
rect 219492 398420 219498 398432
rect 224862 398420 224868 398432
rect 224920 398420 224926 398472
rect 227898 398324 227904 398336
rect 219406 398296 227904 398324
rect 175182 398216 175188 398268
rect 175240 398256 175246 398268
rect 211798 398256 211804 398268
rect 175240 398228 211804 398256
rect 175240 398216 175246 398228
rect 211798 398216 211804 398228
rect 211856 398216 211862 398268
rect 217686 398216 217692 398268
rect 217744 398256 217750 398268
rect 219406 398256 219434 398296
rect 227898 398284 227904 398296
rect 227956 398284 227962 398336
rect 227990 398256 227996 398268
rect 217744 398228 219434 398256
rect 219636 398228 227996 398256
rect 217744 398216 217750 398228
rect 125502 398148 125508 398200
rect 125560 398188 125566 398200
rect 196618 398188 196624 398200
rect 125560 398160 196624 398188
rect 125560 398148 125566 398160
rect 196618 398148 196624 398160
rect 196676 398148 196682 398200
rect 217594 398148 217600 398200
rect 217652 398188 217658 398200
rect 219636 398188 219664 398228
rect 227990 398216 227996 398228
rect 228048 398216 228054 398268
rect 217652 398160 219664 398188
rect 217652 398148 217658 398160
rect 219710 398148 219716 398200
rect 219768 398188 219774 398200
rect 227806 398188 227812 398200
rect 219768 398160 227812 398188
rect 219768 398148 219774 398160
rect 227806 398148 227812 398160
rect 227864 398148 227870 398200
rect 119982 398080 119988 398132
rect 120040 398120 120046 398132
rect 197998 398120 198004 398132
rect 120040 398092 198004 398120
rect 120040 398080 120046 398092
rect 197998 398080 198004 398092
rect 198056 398080 198062 398132
rect 217778 398080 217784 398132
rect 217836 398120 217842 398132
rect 217836 398092 219434 398120
rect 217836 398080 217842 398092
rect 219406 397984 219434 398092
rect 220078 398080 220084 398132
rect 220136 398120 220142 398132
rect 228082 398120 228088 398132
rect 220136 398092 228088 398120
rect 220136 398080 220142 398092
rect 228082 398080 228088 398092
rect 228140 398080 228146 398132
rect 228174 397984 228180 397996
rect 219406 397956 228180 397984
rect 228174 397944 228180 397956
rect 228232 397944 228238 397996
rect 3418 397468 3424 397520
rect 3476 397508 3482 397520
rect 146294 397508 146300 397520
rect 3476 397480 146300 397508
rect 3476 397468 3482 397480
rect 146294 397468 146300 397480
rect 146352 397468 146358 397520
rect 87690 397332 87696 397384
rect 87748 397372 87754 397384
rect 229094 397372 229100 397384
rect 87748 397344 229100 397372
rect 87748 397332 87754 397344
rect 229094 397332 229100 397344
rect 229152 397332 229158 397384
rect 61470 397264 61476 397316
rect 61528 397304 61534 397316
rect 265158 397304 265164 397316
rect 61528 397276 265164 397304
rect 61528 397264 61534 397276
rect 265158 397264 265164 397276
rect 265216 397264 265222 397316
rect 300118 397264 300124 397316
rect 300176 397304 300182 397316
rect 308582 397304 308588 397316
rect 300176 397276 308588 397304
rect 300176 397264 300182 397276
rect 308582 397264 308588 397276
rect 308640 397264 308646 397316
rect 83274 397196 83280 397248
rect 83332 397236 83338 397248
rect 225046 397236 225052 397248
rect 83332 397208 225052 397236
rect 83332 397196 83338 397208
rect 225046 397196 225052 397208
rect 225104 397196 225110 397248
rect 238018 397196 238024 397248
rect 238076 397236 238082 397248
rect 239214 397236 239220 397248
rect 238076 397208 239220 397236
rect 238076 397196 238082 397208
rect 239214 397196 239220 397208
rect 239272 397196 239278 397248
rect 61746 397128 61752 397180
rect 61804 397168 61810 397180
rect 273254 397168 273260 397180
rect 61804 397140 273260 397168
rect 61804 397128 61810 397140
rect 273254 397128 273260 397140
rect 273312 397128 273318 397180
rect 62758 397060 62764 397112
rect 62816 397100 62822 397112
rect 278038 397100 278044 397112
rect 62816 397072 278044 397100
rect 62816 397060 62822 397072
rect 278038 397060 278044 397072
rect 278096 397060 278102 397112
rect 58434 396992 58440 397044
rect 58492 397032 58498 397044
rect 113174 397032 113180 397044
rect 58492 397004 113180 397032
rect 58492 396992 58498 397004
rect 113174 396992 113180 397004
rect 113232 396992 113238 397044
rect 114462 396992 114468 397044
rect 114520 397032 114526 397044
rect 137278 397032 137284 397044
rect 114520 397004 137284 397032
rect 114520 396992 114526 397004
rect 137278 396992 137284 397004
rect 137336 396992 137342 397044
rect 78306 396924 78312 396976
rect 78364 396964 78370 396976
rect 170398 396964 170404 396976
rect 78364 396936 170404 396964
rect 78364 396924 78370 396936
rect 170398 396924 170404 396936
rect 170456 396924 170462 396976
rect 183462 396924 183468 396976
rect 183520 396964 183526 396976
rect 228266 396964 228272 396976
rect 183520 396936 228272 396964
rect 183520 396924 183526 396936
rect 228266 396924 228272 396936
rect 228324 396924 228330 396976
rect 92290 396856 92296 396908
rect 92348 396896 92354 396908
rect 189074 396896 189080 396908
rect 92348 396868 189080 396896
rect 92348 396856 92354 396868
rect 189074 396856 189080 396868
rect 189132 396856 189138 396908
rect 191098 396856 191104 396908
rect 191156 396896 191162 396908
rect 236178 396896 236184 396908
rect 191156 396868 236184 396896
rect 191156 396856 191162 396868
rect 236178 396856 236184 396868
rect 236236 396856 236242 396908
rect 93486 396788 93492 396840
rect 93544 396828 93550 396840
rect 193214 396828 193220 396840
rect 93544 396800 193220 396828
rect 93544 396788 93550 396800
rect 193214 396788 193220 396800
rect 193272 396788 193278 396840
rect 196618 396788 196624 396840
rect 196676 396828 196682 396840
rect 241606 396828 241612 396840
rect 196676 396800 241612 396828
rect 196676 396788 196682 396800
rect 241606 396788 241612 396800
rect 241664 396788 241670 396840
rect 109770 396720 109776 396772
rect 109828 396760 109834 396772
rect 231946 396760 231952 396772
rect 109828 396732 231952 396760
rect 109828 396720 109834 396732
rect 231946 396720 231952 396732
rect 232004 396720 232010 396772
rect 244918 396720 244924 396772
rect 244976 396760 244982 396772
rect 247126 396760 247132 396772
rect 244976 396732 247132 396760
rect 244976 396720 244982 396732
rect 247126 396720 247132 396732
rect 247184 396720 247190 396772
rect 264238 396720 264244 396772
rect 264296 396760 264302 396772
rect 265250 396760 265256 396772
rect 264296 396732 265256 396760
rect 264296 396720 264302 396732
rect 265250 396720 265256 396732
rect 265308 396720 265314 396772
rect 269758 396720 269764 396772
rect 269816 396760 269822 396772
rect 272518 396760 272524 396772
rect 269816 396732 272524 396760
rect 269816 396720 269822 396732
rect 272518 396720 272524 396732
rect 272576 396720 272582 396772
rect 282178 396720 282184 396772
rect 282236 396760 282242 396772
rect 283558 396760 283564 396772
rect 282236 396732 283564 396760
rect 282236 396720 282242 396732
rect 283558 396720 283564 396732
rect 283616 396720 283622 396772
rect 58526 396652 58532 396704
rect 58584 396692 58590 396704
rect 103698 396692 103704 396704
rect 58584 396664 103704 396692
rect 58584 396652 58590 396664
rect 103698 396652 103704 396664
rect 103756 396652 103762 396704
rect 105906 396652 105912 396704
rect 105964 396692 105970 396704
rect 231854 396692 231860 396704
rect 105964 396664 231860 396692
rect 105964 396652 105970 396664
rect 231854 396652 231860 396664
rect 231912 396652 231918 396704
rect 242250 396652 242256 396704
rect 242308 396692 242314 396704
rect 242308 396664 248414 396692
rect 242308 396652 242314 396664
rect 101858 396584 101864 396636
rect 101916 396624 101922 396636
rect 230566 396624 230572 396636
rect 101916 396596 230572 396624
rect 101916 396584 101922 396596
rect 230566 396584 230572 396596
rect 230624 396584 230630 396636
rect 242158 396584 242164 396636
rect 242216 396624 242222 396636
rect 247678 396624 247684 396636
rect 242216 396596 247684 396624
rect 242216 396584 242222 396596
rect 247678 396584 247684 396596
rect 247736 396584 247742 396636
rect 248386 396624 248414 396664
rect 253198 396652 253204 396704
rect 253256 396692 253262 396704
rect 254486 396692 254492 396704
rect 253256 396664 254492 396692
rect 253256 396652 253262 396664
rect 254486 396652 254492 396664
rect 254544 396652 254550 396704
rect 262858 396652 262864 396704
rect 262916 396692 262922 396704
rect 263870 396692 263876 396704
rect 262916 396664 263876 396692
rect 262916 396652 262922 396664
rect 263870 396652 263876 396664
rect 263928 396652 263934 396704
rect 284938 396652 284944 396704
rect 284996 396692 285002 396704
rect 285950 396692 285956 396704
rect 284996 396664 285956 396692
rect 284996 396652 285002 396664
rect 285950 396652 285956 396664
rect 286008 396652 286014 396704
rect 307018 396652 307024 396704
rect 307076 396692 307082 396704
rect 315758 396692 315764 396704
rect 307076 396664 315764 396692
rect 307076 396652 307082 396664
rect 315758 396652 315764 396664
rect 315816 396652 315822 396704
rect 274726 396624 274732 396636
rect 248386 396596 274732 396624
rect 274726 396584 274732 396596
rect 274784 396584 274790 396636
rect 79962 396516 79968 396568
rect 80020 396556 80026 396568
rect 98638 396556 98644 396568
rect 80020 396528 98644 396556
rect 80020 396516 80026 396528
rect 98638 396516 98644 396528
rect 98696 396516 98702 396568
rect 100110 396516 100116 396568
rect 100168 396556 100174 396568
rect 230474 396556 230480 396568
rect 100168 396528 230480 396556
rect 100168 396516 100174 396528
rect 230474 396516 230480 396528
rect 230532 396516 230538 396568
rect 238110 396516 238116 396568
rect 238168 396556 238174 396568
rect 273622 396556 273628 396568
rect 238168 396528 273628 396556
rect 238168 396516 238174 396528
rect 273622 396516 273628 396528
rect 273680 396516 273686 396568
rect 61654 396448 61660 396500
rect 61712 396488 61718 396500
rect 88702 396488 88708 396500
rect 61712 396460 88708 396488
rect 61712 396448 61718 396460
rect 88702 396448 88708 396460
rect 88760 396448 88766 396500
rect 98914 396448 98920 396500
rect 98972 396488 98978 396500
rect 229186 396488 229192 396500
rect 98972 396460 229192 396488
rect 98972 396448 98978 396460
rect 229186 396448 229192 396460
rect 229244 396448 229250 396500
rect 233970 396448 233976 396500
rect 234028 396488 234034 396500
rect 271138 396488 271144 396500
rect 234028 396460 271144 396488
rect 234028 396448 234034 396460
rect 271138 396448 271144 396460
rect 271196 396448 271202 396500
rect 58802 396380 58808 396432
rect 58860 396420 58866 396432
rect 86494 396420 86500 396432
rect 58860 396392 86500 396420
rect 58860 396380 58866 396392
rect 86494 396380 86500 396392
rect 86552 396380 86558 396432
rect 226978 396380 226984 396432
rect 227036 396420 227042 396432
rect 263594 396420 263600 396432
rect 227036 396392 263600 396420
rect 227036 396380 227042 396392
rect 263594 396380 263600 396392
rect 263652 396380 263658 396432
rect 59906 396312 59912 396364
rect 59964 396352 59970 396364
rect 80422 396352 80428 396364
rect 59964 396324 80428 396352
rect 59964 396312 59970 396324
rect 80422 396312 80428 396324
rect 80480 396312 80486 396364
rect 101582 396312 101588 396364
rect 101640 396352 101646 396364
rect 112438 396352 112444 396364
rect 101640 396324 112444 396352
rect 101640 396312 101646 396324
rect 112438 396312 112444 396324
rect 112496 396312 112502 396364
rect 220078 396312 220084 396364
rect 220136 396352 220142 396364
rect 310974 396352 310980 396364
rect 220136 396324 310980 396352
rect 220136 396312 220142 396324
rect 310974 396312 310980 396324
rect 311032 396312 311038 396364
rect 59538 396244 59544 396296
rect 59596 396284 59602 396296
rect 252646 396284 252652 396296
rect 59596 396256 252652 396284
rect 59596 396244 59602 396256
rect 252646 396244 252652 396256
rect 252704 396244 252710 396296
rect 258718 396244 258724 396296
rect 258776 396284 258782 396296
rect 342254 396284 342260 396296
rect 258776 396256 342260 396284
rect 258776 396244 258782 396256
rect 342254 396244 342260 396256
rect 342312 396244 342318 396296
rect 102870 396176 102876 396228
rect 102928 396216 102934 396228
rect 107010 396216 107016 396228
rect 102928 396188 107016 396216
rect 102928 396176 102934 396188
rect 107010 396176 107016 396188
rect 107068 396176 107074 396228
rect 263594 396176 263600 396228
rect 263652 396216 263658 396228
rect 276382 396216 276388 396228
rect 263652 396188 276388 396216
rect 263652 396176 263658 396188
rect 276382 396176 276388 396188
rect 276440 396176 276446 396228
rect 276658 396176 276664 396228
rect 276716 396216 276722 396228
rect 298462 396216 298468 396228
rect 276716 396188 298468 396216
rect 276716 396176 276722 396188
rect 298462 396176 298468 396188
rect 298520 396176 298526 396228
rect 111610 396108 111616 396160
rect 111668 396148 111674 396160
rect 119338 396148 119344 396160
rect 111668 396120 119344 396148
rect 111668 396108 111674 396120
rect 119338 396108 119344 396120
rect 119396 396108 119402 396160
rect 249058 396108 249064 396160
rect 249116 396148 249122 396160
rect 262030 396148 262036 396160
rect 249116 396120 262036 396148
rect 249116 396108 249122 396120
rect 262030 396108 262036 396120
rect 262088 396108 262094 396160
rect 291838 396108 291844 396160
rect 291896 396148 291902 396160
rect 300854 396148 300860 396160
rect 291896 396120 300860 396148
rect 291896 396108 291902 396120
rect 300854 396108 300860 396120
rect 300912 396108 300918 396160
rect 96522 396040 96528 396092
rect 96580 396080 96586 396092
rect 106918 396080 106924 396092
rect 96580 396052 106924 396080
rect 96580 396040 96586 396052
rect 106918 396040 106924 396052
rect 106976 396040 106982 396092
rect 107194 396040 107200 396092
rect 107252 396080 107258 396092
rect 116578 396080 116584 396092
rect 107252 396052 116584 396080
rect 107252 396040 107258 396052
rect 116578 396040 116584 396052
rect 116636 396040 116642 396092
rect 304258 396040 304264 396092
rect 304316 396080 304322 396092
rect 313366 396080 313372 396092
rect 304316 396052 313372 396080
rect 304316 396040 304322 396052
rect 313366 396040 313372 396052
rect 313424 396040 313430 396092
rect 183186 395972 183192 396024
rect 183244 396012 183250 396024
rect 187694 396012 187700 396024
rect 183244 395984 187700 396012
rect 183244 395972 183250 395984
rect 187694 395972 187700 395984
rect 187752 395972 187758 396024
rect 232498 395972 232504 396024
rect 232556 396012 232562 396024
rect 250070 396012 250076 396024
rect 232556 395984 250076 396012
rect 232556 395972 232562 395984
rect 250070 395972 250076 395984
rect 250128 395972 250134 396024
rect 179322 395904 179328 395956
rect 179380 395944 179386 395956
rect 244458 395944 244464 395956
rect 179380 395916 244464 395944
rect 179380 395904 179386 395916
rect 244458 395904 244464 395916
rect 244516 395904 244522 395956
rect 113634 395836 113640 395888
rect 113692 395876 113698 395888
rect 194594 395876 194600 395888
rect 113692 395848 194600 395876
rect 113692 395836 113698 395848
rect 194594 395836 194600 395848
rect 194652 395836 194658 395888
rect 233878 395836 233884 395888
rect 233936 395876 233942 395888
rect 256142 395876 256148 395888
rect 233936 395848 256148 395876
rect 233936 395836 233942 395848
rect 256142 395836 256148 395848
rect 256200 395836 256206 395888
rect 138474 395768 138480 395820
rect 138532 395808 138538 395820
rect 228542 395808 228548 395820
rect 138532 395780 228548 395808
rect 138532 395768 138538 395780
rect 228542 395768 228548 395780
rect 228600 395768 228606 395820
rect 231118 395768 231124 395820
rect 231176 395808 231182 395820
rect 260926 395808 260932 395820
rect 231176 395780 260932 395808
rect 231176 395768 231182 395780
rect 260926 395768 260932 395780
rect 260984 395768 260990 395820
rect 56318 395700 56324 395752
rect 56376 395740 56382 395752
rect 118142 395740 118148 395752
rect 56376 395712 118148 395740
rect 56376 395700 56382 395712
rect 118142 395700 118148 395712
rect 118200 395700 118206 395752
rect 136450 395700 136456 395752
rect 136508 395740 136514 395752
rect 228450 395740 228456 395752
rect 136508 395712 228456 395740
rect 136508 395700 136514 395712
rect 228450 395700 228456 395712
rect 228508 395700 228514 395752
rect 235258 395700 235264 395752
rect 235316 395740 235322 395752
rect 273438 395740 273444 395752
rect 235316 395712 273444 395740
rect 235316 395700 235322 395712
rect 273438 395700 273444 395712
rect 273496 395700 273502 395752
rect 54662 395632 54668 395684
rect 54720 395672 54726 395684
rect 150710 395672 150716 395684
rect 54720 395644 150716 395672
rect 54720 395632 54726 395644
rect 150710 395632 150716 395644
rect 150768 395632 150774 395684
rect 177942 395632 177948 395684
rect 178000 395672 178006 395684
rect 253566 395672 253572 395684
rect 178000 395644 253572 395672
rect 178000 395632 178006 395644
rect 253566 395632 253572 395644
rect 253624 395632 253630 395684
rect 54846 395564 54852 395616
rect 54904 395604 54910 395616
rect 98454 395604 98460 395616
rect 54904 395576 98460 395604
rect 54904 395564 54910 395576
rect 98454 395564 98460 395576
rect 98512 395564 98518 395616
rect 115842 395564 115848 395616
rect 115900 395604 115906 395616
rect 222194 395604 222200 395616
rect 115900 395576 222200 395604
rect 115900 395564 115906 395576
rect 222194 395564 222200 395576
rect 222252 395564 222258 395616
rect 224678 395564 224684 395616
rect 224736 395604 224742 395616
rect 263594 395604 263600 395616
rect 224736 395576 263600 395604
rect 224736 395564 224742 395576
rect 263594 395564 263600 395576
rect 263652 395564 263658 395616
rect 96430 395496 96436 395548
rect 96488 395536 96494 395548
rect 229278 395536 229284 395548
rect 96488 395508 229284 395536
rect 96488 395496 96494 395508
rect 229278 395496 229284 395508
rect 229336 395496 229342 395548
rect 231210 395496 231216 395548
rect 231268 395536 231274 395548
rect 293310 395536 293316 395548
rect 231268 395508 293316 395536
rect 231268 395496 231274 395508
rect 293310 395496 293316 395508
rect 293368 395496 293374 395548
rect 52362 395428 52368 395480
rect 52420 395468 52426 395480
rect 242894 395468 242900 395480
rect 52420 395440 242900 395468
rect 52420 395428 52426 395440
rect 242894 395428 242900 395440
rect 242952 395428 242958 395480
rect 52178 395360 52184 395412
rect 52236 395400 52242 395412
rect 248598 395400 248604 395412
rect 52236 395372 248604 395400
rect 52236 395360 52242 395372
rect 248598 395360 248604 395372
rect 248656 395360 248662 395412
rect 54754 395292 54760 395344
rect 54812 395332 54818 395344
rect 290182 395332 290188 395344
rect 54812 395304 290188 395332
rect 54812 395292 54818 395304
rect 290182 395292 290188 395304
rect 290240 395292 290246 395344
rect 196894 393360 196900 393372
rect 194704 393332 196900 393360
rect 193306 393252 193312 393304
rect 193364 393292 193370 393304
rect 194704 393292 194732 393332
rect 196894 393320 196900 393332
rect 196952 393320 196958 393372
rect 193364 393264 194732 393292
rect 193364 393252 193370 393264
rect 219066 392912 219072 392964
rect 219124 392952 219130 392964
rect 219342 392952 219348 392964
rect 219124 392924 219348 392952
rect 219124 392912 219130 392924
rect 219342 392912 219348 392924
rect 219400 392912 219406 392964
rect 191374 390328 191380 390380
rect 191432 390368 191438 390380
rect 193306 390368 193312 390380
rect 191432 390340 193312 390368
rect 191432 390328 191438 390340
rect 193306 390328 193312 390340
rect 193364 390328 193370 390380
rect 186314 387812 186320 387864
rect 186372 387852 186378 387864
rect 191374 387852 191380 387864
rect 186372 387824 191380 387852
rect 186372 387812 186378 387824
rect 191374 387812 191380 387824
rect 191432 387812 191438 387864
rect 185670 385636 185676 385688
rect 185728 385676 185734 385688
rect 186314 385676 186320 385688
rect 185728 385648 186320 385676
rect 185728 385636 185734 385648
rect 186314 385636 186320 385648
rect 186372 385636 186378 385688
rect 219066 383732 219072 383784
rect 219124 383772 219130 383784
rect 219124 383744 219388 383772
rect 219124 383732 219130 383744
rect 219360 383716 219388 383744
rect 219342 383664 219348 383716
rect 219400 383664 219406 383716
rect 183554 379516 183560 379568
rect 183612 379556 183618 379568
rect 185670 379556 185676 379568
rect 183612 379528 185676 379556
rect 183612 379516 183618 379528
rect 185670 379516 185676 379528
rect 185728 379516 185734 379568
rect 85390 378768 85396 378820
rect 85448 378808 85454 378820
rect 232130 378808 232136 378820
rect 85448 378780 232136 378808
rect 85448 378768 85454 378780
rect 232130 378768 232136 378780
rect 232188 378768 232194 378820
rect 85390 378156 85396 378208
rect 85448 378196 85454 378208
rect 580166 378196 580172 378208
rect 85448 378168 580172 378196
rect 85448 378156 85454 378168
rect 580166 378156 580172 378168
rect 580224 378156 580230 378208
rect 177298 374620 177304 374672
rect 177356 374660 177362 374672
rect 183554 374660 183560 374672
rect 177356 374632 183560 374660
rect 177356 374620 177362 374632
rect 183554 374620 183560 374632
rect 183612 374620 183618 374672
rect 3418 371220 3424 371272
rect 3476 371260 3482 371272
rect 149054 371260 149060 371272
rect 3476 371232 149060 371260
rect 3476 371220 3482 371232
rect 149054 371220 149060 371232
rect 149112 371220 149118 371272
rect 86862 364352 86868 364404
rect 86920 364392 86926 364404
rect 579614 364392 579620 364404
rect 86920 364364 579620 364392
rect 86920 364352 86926 364364
rect 579614 364352 579620 364364
rect 579672 364352 579678 364404
rect 177298 360244 177304 360256
rect 173912 360216 177304 360244
rect 173434 360136 173440 360188
rect 173492 360176 173498 360188
rect 173912 360176 173940 360216
rect 177298 360204 177304 360216
rect 177356 360204 177362 360256
rect 173492 360148 173940 360176
rect 173492 360136 173498 360148
rect 171778 358504 171784 358556
rect 171836 358544 171842 358556
rect 173434 358544 173440 358556
rect 171836 358516 173440 358544
rect 171836 358504 171842 358516
rect 173434 358504 173440 358516
rect 173492 358504 173498 358556
rect 119890 358028 119896 358080
rect 119948 358068 119954 358080
rect 223574 358068 223580 358080
rect 119948 358040 223580 358068
rect 119948 358028 119954 358040
rect 223574 358028 223580 358040
rect 223632 358028 223638 358080
rect 3142 357416 3148 357468
rect 3200 357456 3206 357468
rect 150434 357456 150440 357468
rect 3200 357428 150440 357456
rect 3200 357416 3206 357428
rect 150434 357416 150440 357428
rect 150492 357416 150498 357468
rect 170490 352044 170496 352096
rect 170548 352084 170554 352096
rect 171778 352084 171784 352096
rect 170548 352056 171784 352084
rect 170548 352044 170554 352056
rect 171778 352044 171784 352056
rect 171836 352044 171842 352096
rect 84102 351908 84108 351960
rect 84160 351948 84166 351960
rect 580166 351948 580172 351960
rect 84160 351920 580172 351948
rect 84160 351908 84166 351920
rect 580166 351908 580172 351920
rect 580224 351908 580230 351960
rect 3326 345040 3332 345092
rect 3384 345080 3390 345092
rect 149146 345080 149152 345092
rect 3384 345052 149152 345080
rect 3384 345040 3390 345052
rect 149146 345040 149152 345052
rect 149204 345040 149210 345092
rect 166718 340892 166724 340944
rect 166776 340932 166782 340944
rect 170490 340932 170496 340944
rect 166776 340904 170496 340932
rect 166776 340892 166782 340904
rect 170490 340892 170496 340904
rect 170548 340892 170554 340944
rect 166718 338144 166724 338156
rect 164252 338116 166724 338144
rect 162854 338036 162860 338088
rect 162912 338076 162918 338088
rect 164252 338076 164280 338116
rect 166718 338104 166724 338116
rect 166776 338104 166782 338156
rect 162912 338048 164280 338076
rect 162912 338036 162918 338048
rect 219066 335112 219072 335164
rect 219124 335152 219130 335164
rect 219342 335152 219348 335164
rect 219124 335124 219348 335152
rect 219124 335112 219130 335124
rect 219342 335112 219348 335124
rect 219400 335112 219406 335164
rect 162854 331276 162860 331288
rect 158732 331248 162860 331276
rect 156598 331168 156604 331220
rect 156656 331208 156662 331220
rect 158732 331208 158760 331248
rect 162854 331236 162860 331248
rect 162912 331236 162918 331288
rect 156656 331180 158760 331208
rect 156656 331168 156662 331180
rect 219066 325796 219072 325848
rect 219124 325836 219130 325848
rect 219342 325836 219348 325848
rect 219124 325808 219348 325836
rect 219124 325796 219130 325808
rect 219342 325796 219348 325808
rect 219400 325796 219406 325848
rect 82630 324300 82636 324352
rect 82688 324340 82694 324352
rect 580166 324340 580172 324352
rect 82688 324312 580172 324340
rect 82688 324300 82694 324312
rect 580166 324300 580172 324312
rect 580224 324300 580230 324352
rect 155218 320424 155224 320476
rect 155276 320464 155282 320476
rect 156598 320464 156604 320476
rect 155276 320436 156604 320464
rect 155276 320424 155282 320436
rect 156598 320424 156604 320436
rect 156656 320424 156662 320476
rect 131022 319404 131028 319456
rect 131080 319444 131086 319456
rect 228726 319444 228732 319456
rect 131080 319416 228732 319444
rect 131080 319404 131086 319416
rect 228726 319404 228732 319416
rect 228784 319404 228790 319456
rect 3418 318792 3424 318844
rect 3476 318832 3482 318844
rect 151814 318832 151820 318844
rect 3476 318804 151820 318832
rect 3476 318792 3482 318804
rect 151814 318792 151820 318804
rect 151872 318792 151878 318844
rect 84010 311856 84016 311908
rect 84068 311896 84074 311908
rect 579982 311896 579988 311908
rect 84068 311868 579988 311896
rect 84068 311856 84074 311868
rect 579982 311856 579988 311868
rect 580040 311856 580046 311908
rect 154482 305600 154488 305652
rect 154540 305640 154546 305652
rect 228358 305640 228364 305652
rect 154540 305612 228364 305640
rect 154540 305600 154546 305612
rect 228358 305600 228364 305612
rect 228416 305600 228422 305652
rect 3234 304988 3240 305040
rect 3292 305028 3298 305040
rect 153194 305028 153200 305040
rect 3292 305000 153200 305028
rect 3292 304988 3298 305000
rect 153194 304988 153200 305000
rect 153252 304988 153258 305040
rect 153838 301520 153844 301572
rect 153896 301560 153902 301572
rect 155218 301560 155224 301572
rect 153896 301532 155224 301560
rect 153896 301520 153902 301532
rect 155218 301520 155224 301532
rect 155276 301520 155282 301572
rect 191650 301452 191656 301504
rect 191708 301492 191714 301504
rect 342346 301492 342352 301504
rect 191708 301464 342352 301492
rect 191708 301452 191714 301464
rect 342346 301452 342352 301464
rect 342404 301452 342410 301504
rect 97810 300092 97816 300144
rect 97868 300132 97874 300144
rect 376018 300132 376024 300144
rect 97868 300104 376024 300132
rect 97868 300092 97874 300104
rect 376018 300092 376024 300104
rect 376076 300092 376082 300144
rect 95050 298732 95056 298784
rect 95108 298772 95114 298784
rect 378778 298772 378784 298784
rect 95108 298744 378784 298772
rect 95108 298732 95114 298744
rect 378778 298732 378784 298744
rect 378836 298732 378842 298784
rect 81342 298120 81348 298172
rect 81400 298160 81406 298172
rect 580166 298160 580172 298172
rect 81400 298132 580172 298160
rect 81400 298120 81406 298132
rect 580166 298120 580172 298132
rect 580224 298120 580230 298172
rect 18598 297372 18604 297424
rect 18656 297412 18662 297424
rect 142154 297412 142160 297424
rect 18656 297384 142160 297412
rect 18656 297372 18662 297384
rect 142154 297372 142160 297384
rect 142212 297372 142218 297424
rect 112990 294652 112996 294704
rect 113048 294692 113054 294704
rect 412634 294692 412640 294704
rect 113048 294664 412640 294692
rect 113048 294652 113054 294664
rect 412634 294652 412640 294664
rect 412692 294652 412698 294704
rect 107470 294584 107476 294636
rect 107528 294624 107534 294636
rect 542354 294624 542360 294636
rect 107528 294596 542360 294624
rect 107528 294584 107534 294596
rect 542354 294584 542360 294596
rect 542412 294584 542418 294636
rect 3418 292544 3424 292596
rect 3476 292584 3482 292596
rect 153286 292584 153292 292596
rect 3476 292556 153292 292584
rect 3476 292544 3482 292556
rect 153286 292544 153292 292556
rect 153344 292544 153350 292596
rect 14458 290436 14464 290488
rect 14516 290476 14522 290488
rect 133874 290476 133880 290488
rect 14516 290448 133880 290476
rect 14516 290436 14522 290448
rect 133874 290436 133880 290448
rect 133932 290436 133938 290488
rect 111610 284928 111616 284980
rect 111668 284968 111674 284980
rect 429194 284968 429200 284980
rect 111668 284940 429200 284968
rect 111668 284928 111674 284940
rect 429194 284928 429200 284940
rect 429252 284928 429258 284980
rect 152826 276020 152832 276072
rect 152884 276060 152890 276072
rect 153838 276060 153844 276072
rect 152884 276032 153844 276060
rect 152884 276020 152890 276032
rect 153838 276020 153844 276032
rect 153896 276020 153902 276072
rect 79962 271872 79968 271924
rect 80020 271912 80026 271924
rect 580166 271912 580172 271924
rect 80020 271884 580172 271912
rect 80020 271872 80026 271884
rect 580166 271872 580172 271884
rect 580224 271872 580230 271924
rect 144822 269764 144828 269816
rect 144880 269804 144886 269816
rect 213914 269804 213920 269816
rect 144880 269776 213920 269804
rect 144880 269764 144886 269776
rect 213914 269764 213920 269776
rect 213972 269764 213978 269816
rect 150526 269084 150532 269136
rect 150584 269124 150590 269136
rect 152826 269124 152832 269136
rect 150584 269096 152832 269124
rect 150584 269084 150590 269096
rect 152826 269084 152832 269096
rect 152884 269084 152890 269136
rect 52086 268336 52092 268388
rect 52144 268376 52150 268388
rect 258166 268376 258172 268388
rect 52144 268348 258172 268376
rect 52144 268336 52150 268348
rect 258166 268336 258172 268348
rect 258224 268336 258230 268388
rect 176562 267044 176568 267096
rect 176620 267084 176626 267096
rect 191098 267084 191104 267096
rect 176620 267056 191104 267084
rect 176620 267044 176626 267056
rect 191098 267044 191104 267056
rect 191156 267044 191162 267096
rect 98638 266976 98644 267028
rect 98696 267016 98702 267028
rect 176654 267016 176660 267028
rect 98696 266988 176660 267016
rect 98696 266976 98702 266988
rect 176654 266976 176660 266988
rect 176712 266976 176718 267028
rect 182082 266976 182088 267028
rect 182140 267016 182146 267028
rect 204990 267016 204996 267028
rect 182140 266988 204996 267016
rect 182140 266976 182146 266988
rect 204990 266976 204996 266988
rect 205048 266976 205054 267028
rect 213178 266976 213184 267028
rect 213236 267016 213242 267028
rect 266446 267016 266452 267028
rect 213236 266988 266452 267016
rect 213236 266976 213242 266988
rect 266446 266976 266452 266988
rect 266504 266976 266510 267028
rect 3050 266364 3056 266416
rect 3108 266404 3114 266416
rect 154574 266404 154580 266416
rect 3108 266376 154580 266404
rect 3108 266364 3114 266376
rect 154574 266364 154580 266376
rect 154632 266364 154638 266416
rect 112438 266296 112444 266348
rect 112496 266336 112502 266348
rect 204254 266336 204260 266348
rect 112496 266308 204260 266336
rect 112496 266296 112502 266308
rect 204254 266296 204260 266308
rect 204312 266296 204318 266348
rect 116578 266228 116584 266280
rect 116636 266268 116642 266280
rect 211154 266268 211160 266280
rect 116636 266240 211160 266268
rect 116636 266228 116642 266240
rect 211154 266228 211160 266240
rect 211212 266228 211218 266280
rect 107010 266160 107016 266212
rect 107068 266200 107074 266212
rect 207014 266200 207020 266212
rect 107068 266172 207020 266200
rect 107068 266160 107074 266172
rect 207014 266160 207020 266172
rect 207072 266160 207078 266212
rect 101950 266092 101956 266144
rect 102008 266132 102014 266144
rect 225138 266132 225144 266144
rect 102008 266104 225144 266132
rect 102008 266092 102014 266104
rect 225138 266092 225144 266104
rect 225196 266092 225202 266144
rect 107378 266024 107384 266076
rect 107436 266064 107442 266076
rect 232406 266064 232412 266076
rect 107436 266036 232412 266064
rect 107436 266024 107442 266036
rect 232406 266024 232412 266036
rect 232464 266024 232470 266076
rect 82722 265956 82728 266008
rect 82780 265996 82786 266008
rect 233510 265996 233516 266008
rect 82780 265968 233516 265996
rect 82780 265956 82786 265968
rect 233510 265956 233516 265968
rect 233568 265956 233574 266008
rect 77202 265888 77208 265940
rect 77260 265928 77266 265940
rect 232222 265928 232228 265940
rect 77260 265900 232228 265928
rect 77260 265888 77266 265900
rect 232222 265888 232228 265900
rect 232280 265888 232286 265940
rect 57146 265820 57152 265872
rect 57204 265860 57210 265872
rect 213270 265860 213276 265872
rect 57204 265832 213276 265860
rect 57204 265820 57210 265832
rect 213270 265820 213276 265832
rect 213328 265820 213334 265872
rect 51994 265752 52000 265804
rect 52052 265792 52058 265804
rect 259546 265792 259552 265804
rect 52052 265764 259552 265792
rect 52052 265752 52058 265764
rect 259546 265752 259552 265764
rect 259604 265752 259610 265804
rect 61562 265684 61568 265736
rect 61620 265724 61626 265736
rect 278774 265724 278780 265736
rect 61620 265696 278780 265724
rect 61620 265684 61626 265696
rect 278774 265684 278780 265696
rect 278832 265684 278838 265736
rect 56226 265616 56232 265668
rect 56284 265656 56290 265668
rect 325694 265656 325700 265668
rect 56284 265628 325700 265656
rect 56284 265616 56290 265628
rect 325694 265616 325700 265628
rect 325752 265616 325758 265668
rect 137278 265548 137284 265600
rect 137336 265588 137342 265600
rect 219434 265588 219440 265600
rect 137336 265560 219440 265588
rect 137336 265548 137342 265560
rect 219434 265548 219440 265560
rect 219492 265548 219498 265600
rect 111518 265480 111524 265532
rect 111576 265520 111582 265532
rect 191834 265520 191840 265532
rect 111576 265492 191840 265520
rect 111576 265480 111582 265492
rect 191834 265480 191840 265492
rect 191892 265480 191898 265532
rect 197262 265480 197268 265532
rect 197320 265520 197326 265532
rect 276106 265520 276112 265532
rect 197320 265492 276112 265520
rect 197320 265480 197326 265492
rect 276106 265480 276112 265492
rect 276164 265480 276170 265532
rect 195882 265412 195888 265464
rect 195940 265452 195946 265464
rect 253198 265452 253204 265464
rect 195940 265424 253204 265452
rect 195940 265412 195946 265424
rect 253198 265412 253204 265424
rect 253256 265412 253262 265464
rect 50338 264868 50344 264920
rect 50396 264908 50402 264920
rect 147766 264908 147772 264920
rect 50396 264880 147772 264908
rect 50396 264868 50402 264880
rect 147766 264868 147772 264880
rect 147824 264868 147830 264920
rect 47578 264800 47584 264852
rect 47636 264840 47642 264852
rect 144914 264840 144920 264852
rect 47636 264812 144920 264840
rect 47636 264800 47642 264812
rect 144914 264800 144920 264812
rect 144972 264800 144978 264852
rect 43438 264732 43444 264784
rect 43496 264772 43502 264784
rect 142246 264772 142252 264784
rect 43496 264744 142252 264772
rect 43496 264732 43502 264744
rect 142246 264732 142252 264744
rect 142304 264732 142310 264784
rect 164142 264732 164148 264784
rect 164200 264772 164206 264784
rect 229370 264772 229376 264784
rect 164200 264744 229376 264772
rect 164200 264732 164206 264744
rect 229370 264732 229376 264744
rect 229428 264732 229434 264784
rect 97902 264664 97908 264716
rect 97960 264704 97966 264716
rect 197538 264704 197544 264716
rect 97960 264676 197544 264704
rect 97960 264664 97966 264676
rect 197538 264664 197544 264676
rect 197596 264664 197602 264716
rect 209682 264664 209688 264716
rect 209740 264704 209746 264716
rect 262858 264704 262864 264716
rect 209740 264676 262864 264704
rect 209740 264664 209746 264676
rect 262858 264664 262864 264676
rect 262916 264664 262922 264716
rect 93762 264596 93768 264648
rect 93820 264636 93826 264648
rect 228634 264636 228640 264648
rect 93820 264608 228640 264636
rect 93820 264596 93826 264608
rect 228634 264596 228640 264608
rect 228692 264596 228698 264648
rect 95142 264528 95148 264580
rect 95200 264568 95206 264580
rect 230658 264568 230664 264580
rect 95200 264540 230664 264568
rect 95200 264528 95206 264540
rect 230658 264528 230664 264540
rect 230716 264528 230722 264580
rect 91002 264460 91008 264512
rect 91060 264500 91066 264512
rect 232314 264500 232320 264512
rect 91060 264472 232320 264500
rect 91060 264460 91066 264472
rect 232314 264460 232320 264472
rect 232372 264460 232378 264512
rect 234062 264460 234068 264512
rect 234120 264500 234126 264512
rect 256694 264500 256700 264512
rect 234120 264472 256700 264500
rect 234120 264460 234126 264472
rect 256694 264460 256700 264472
rect 256752 264460 256758 264512
rect 54478 264392 54484 264444
rect 54536 264432 54542 264444
rect 280154 264432 280160 264444
rect 54536 264404 280160 264432
rect 54536 264392 54542 264404
rect 280154 264392 280160 264404
rect 280212 264392 280218 264444
rect 54386 264324 54392 264376
rect 54444 264364 54450 264376
rect 295334 264364 295340 264376
rect 54444 264336 295340 264364
rect 54444 264324 54450 264336
rect 295334 264324 295340 264336
rect 295392 264324 295398 264376
rect 54294 264256 54300 264308
rect 54352 264296 54358 264308
rect 304994 264296 305000 264308
rect 54352 264268 305000 264296
rect 54352 264256 54358 264268
rect 304994 264256 305000 264268
rect 305052 264256 305058 264308
rect 89530 264188 89536 264240
rect 89588 264228 89594 264240
rect 580258 264228 580264 264240
rect 89588 264200 580264 264228
rect 89588 264188 89594 264200
rect 580258 264188 580264 264200
rect 580316 264188 580322 264240
rect 35158 264120 35164 264172
rect 35216 264160 35222 264172
rect 132494 264160 132500 264172
rect 35216 264132 132500 264160
rect 35216 264120 35222 264132
rect 132494 264120 132500 264132
rect 132552 264120 132558 264172
rect 133782 264120 133788 264172
rect 133840 264160 133846 264172
rect 208394 264160 208400 264172
rect 133840 264132 208400 264160
rect 133840 264120 133846 264132
rect 208394 264120 208400 264132
rect 208452 264120 208458 264172
rect 119338 264052 119344 264104
rect 119396 264092 119402 264104
rect 215294 264092 215300 264104
rect 119396 264064 215300 264092
rect 119396 264052 119402 264064
rect 215294 264052 215300 264064
rect 215352 264052 215358 264104
rect 106918 263984 106924 264036
rect 106976 264024 106982 264036
rect 197446 264024 197452 264036
rect 106976 263996 197452 264024
rect 106976 263984 106982 263996
rect 197446 263984 197452 263996
rect 197504 263984 197510 264036
rect 56042 263916 56048 263968
rect 56100 263956 56106 263968
rect 140774 263956 140780 263968
rect 56100 263928 140780 263956
rect 56100 263916 56106 263928
rect 140774 263916 140780 263928
rect 140832 263916 140838 263968
rect 126882 263848 126888 263900
rect 126940 263888 126946 263900
rect 201678 263888 201684 263900
rect 126940 263860 201684 263888
rect 126940 263848 126946 263860
rect 201678 263848 201684 263860
rect 201736 263848 201742 263900
rect 149238 263576 149244 263628
rect 149296 263616 149302 263628
rect 150526 263616 150532 263628
rect 149296 263588 150532 263616
rect 149296 263576 149302 263588
rect 150526 263576 150532 263588
rect 150584 263576 150590 263628
rect 29638 263508 29644 263560
rect 29696 263548 29702 263560
rect 140774 263548 140780 263560
rect 29696 263520 140780 263548
rect 29696 263508 29702 263520
rect 140774 263508 140780 263520
rect 140832 263508 140838 263560
rect 213822 263508 213828 263560
rect 213880 263548 213886 263560
rect 291838 263548 291844 263560
rect 213880 263520 291844 263548
rect 213880 263508 213886 263520
rect 291838 263508 291844 263520
rect 291896 263508 291902 263560
rect 8202 263440 8208 263492
rect 8260 263480 8266 263492
rect 128354 263480 128360 263492
rect 8260 263452 128360 263480
rect 8260 263440 8266 263452
rect 128354 263440 128360 263452
rect 128412 263440 128418 263492
rect 181990 263440 181996 263492
rect 182048 263480 182054 263492
rect 196618 263480 196624 263492
rect 182048 263452 196624 263480
rect 182048 263440 182054 263452
rect 196618 263440 196624 263452
rect 196676 263440 196682 263492
rect 205542 263440 205548 263492
rect 205600 263480 205606 263492
rect 287054 263480 287060 263492
rect 205600 263452 287060 263480
rect 205600 263440 205606 263452
rect 287054 263440 287060 263452
rect 287112 263440 287118 263492
rect 108850 263372 108856 263424
rect 108908 263412 108914 263424
rect 230842 263412 230848 263424
rect 108908 263384 230848 263412
rect 108908 263372 108914 263384
rect 230842 263372 230848 263384
rect 230900 263372 230906 263424
rect 235350 263372 235356 263424
rect 235408 263412 235414 263424
rect 358814 263412 358820 263424
rect 235408 263384 358820 263412
rect 235408 263372 235414 263384
rect 358814 263372 358820 263384
rect 358872 263372 358878 263424
rect 111702 263304 111708 263356
rect 111760 263344 111766 263356
rect 388438 263344 388444 263356
rect 111760 263316 388444 263344
rect 111760 263304 111766 263316
rect 388438 263304 388444 263316
rect 388496 263304 388502 263356
rect 108850 263236 108856 263288
rect 108908 263276 108914 263288
rect 385678 263276 385684 263288
rect 108908 263248 385684 263276
rect 108908 263236 108914 263248
rect 385678 263236 385684 263248
rect 385736 263236 385742 263288
rect 102042 263168 102048 263220
rect 102100 263208 102106 263220
rect 396718 263208 396724 263220
rect 102100 263180 396724 263208
rect 102100 263168 102106 263180
rect 396718 263168 396724 263180
rect 396776 263168 396782 263220
rect 104710 263100 104716 263152
rect 104768 263140 104774 263152
rect 399478 263140 399484 263152
rect 104768 263112 399484 263140
rect 104768 263100 104774 263112
rect 399478 263100 399484 263112
rect 399536 263100 399542 263152
rect 97902 263032 97908 263084
rect 97960 263072 97966 263084
rect 395338 263072 395344 263084
rect 97960 263044 395344 263072
rect 97960 263032 97966 263044
rect 395338 263032 395344 263044
rect 395396 263032 395402 263084
rect 95142 262964 95148 263016
rect 95200 263004 95206 263016
rect 393958 263004 393964 263016
rect 95200 262976 393964 263004
rect 95200 262964 95206 262976
rect 393958 262964 393964 262976
rect 394016 262964 394022 263016
rect 92382 262896 92388 262948
rect 92440 262936 92446 262948
rect 392578 262936 392584 262948
rect 92440 262908 392584 262936
rect 92440 262896 92446 262908
rect 392578 262896 392584 262908
rect 392636 262896 392642 262948
rect 88242 262828 88248 262880
rect 88300 262868 88306 262880
rect 389818 262868 389824 262880
rect 88300 262840 389824 262868
rect 88300 262828 88306 262840
rect 389818 262828 389824 262840
rect 389876 262828 389882 262880
rect 32398 262760 32404 262812
rect 32456 262800 32462 262812
rect 143534 262800 143540 262812
rect 32456 262772 143540 262800
rect 32456 262760 32462 262772
rect 143534 262760 143540 262772
rect 143592 262760 143598 262812
rect 201402 262760 201408 262812
rect 201460 262800 201466 262812
rect 259454 262800 259460 262812
rect 201460 262772 259460 262800
rect 201460 262760 201466 262772
rect 259454 262760 259460 262772
rect 259512 262760 259518 262812
rect 39298 262692 39304 262744
rect 39356 262732 39362 262744
rect 138014 262732 138020 262744
rect 39356 262704 138020 262732
rect 39356 262692 39362 262704
rect 138014 262692 138020 262704
rect 138072 262692 138078 262744
rect 36538 262624 36544 262676
rect 36596 262664 36602 262676
rect 135254 262664 135260 262676
rect 36596 262636 135260 262664
rect 36596 262624 36602 262636
rect 135254 262624 135260 262636
rect 135312 262624 135318 262676
rect 33778 262556 33784 262608
rect 33836 262596 33842 262608
rect 129734 262596 129740 262608
rect 33836 262568 129740 262596
rect 33836 262556 33842 262568
rect 129734 262556 129740 262568
rect 129792 262556 129798 262608
rect 55950 262488 55956 262540
rect 56008 262528 56014 262540
rect 147674 262528 147680 262540
rect 56008 262500 147680 262528
rect 56008 262488 56014 262500
rect 147674 262488 147680 262500
rect 147732 262488 147738 262540
rect 118510 262420 118516 262472
rect 118568 262460 118574 262472
rect 200758 262460 200764 262472
rect 118568 262432 200764 262460
rect 118568 262420 118574 262432
rect 200758 262420 200764 262432
rect 200816 262420 200822 262472
rect 129642 262352 129648 262404
rect 129700 262392 129706 262404
rect 205634 262392 205640 262404
rect 129700 262364 205640 262392
rect 129700 262352 129706 262364
rect 205634 262352 205640 262364
rect 205692 262352 205698 262404
rect 11698 262148 11704 262200
rect 11756 262188 11762 262200
rect 136634 262188 136640 262200
rect 11756 262160 136640 262188
rect 11756 262148 11762 262160
rect 136634 262148 136640 262160
rect 136692 262148 136698 262200
rect 146938 262148 146944 262200
rect 146996 262188 147002 262200
rect 149238 262188 149244 262200
rect 146996 262160 149244 262188
rect 146996 262148 147002 262160
rect 149238 262148 149244 262160
rect 149296 262148 149302 262200
rect 202782 262148 202788 262200
rect 202840 262188 202846 262200
rect 284938 262188 284944 262200
rect 202840 262160 284944 262188
rect 202840 262148 202846 262160
rect 284938 262148 284944 262160
rect 284996 262148 285002 262200
rect 21358 262080 21364 262132
rect 21416 262120 21422 262132
rect 146386 262120 146392 262132
rect 21416 262092 146392 262120
rect 21416 262080 21422 262092
rect 146386 262080 146392 262092
rect 146444 262080 146450 262132
rect 170398 262080 170404 262132
rect 170456 262120 170462 262132
rect 173894 262120 173900 262132
rect 170456 262092 173900 262120
rect 170456 262080 170462 262092
rect 173894 262080 173900 262092
rect 173952 262080 173958 262132
rect 218974 262080 218980 262132
rect 219032 262120 219038 262132
rect 307018 262120 307024 262132
rect 219032 262092 307024 262120
rect 219032 262080 219038 262092
rect 307018 262080 307024 262092
rect 307076 262080 307082 262132
rect 53190 262012 53196 262064
rect 53248 262052 53254 262064
rect 198918 262052 198924 262064
rect 53248 262024 198924 262052
rect 53248 262012 53254 262024
rect 198918 262012 198924 262024
rect 198976 262012 198982 262064
rect 222102 262012 222108 262064
rect 222160 262052 222166 262064
rect 317414 262052 317420 262064
rect 222160 262024 317420 262052
rect 222160 262012 222166 262024
rect 317414 262012 317420 262024
rect 317472 262012 317478 262064
rect 108758 261944 108764 261996
rect 108816 261984 108822 261996
rect 370498 261984 370504 261996
rect 108816 261956 370504 261984
rect 108816 261944 108822 261956
rect 370498 261944 370504 261956
rect 370556 261944 370562 261996
rect 99282 261876 99288 261928
rect 99340 261916 99346 261928
rect 367738 261916 367744 261928
rect 99340 261888 367744 261916
rect 99340 261876 99346 261888
rect 367738 261876 367744 261888
rect 367796 261876 367802 261928
rect 100662 261808 100668 261860
rect 100720 261848 100726 261860
rect 377398 261848 377404 261860
rect 100720 261820 377404 261848
rect 100720 261808 100726 261820
rect 377398 261808 377404 261820
rect 377456 261808 377462 261860
rect 106090 261740 106096 261792
rect 106148 261780 106154 261792
rect 382918 261780 382924 261792
rect 106148 261752 382924 261780
rect 106148 261740 106154 261752
rect 382918 261740 382924 261752
rect 382976 261740 382982 261792
rect 103422 261672 103428 261724
rect 103480 261712 103486 261724
rect 381538 261712 381544 261724
rect 103480 261684 381544 261712
rect 103480 261672 103486 261684
rect 381538 261672 381544 261684
rect 381596 261672 381602 261724
rect 91002 261604 91008 261656
rect 91060 261644 91066 261656
rect 374638 261644 374644 261656
rect 91060 261616 374644 261644
rect 91060 261604 91066 261616
rect 374638 261604 374644 261616
rect 374696 261604 374702 261656
rect 88150 261536 88156 261588
rect 88208 261576 88214 261588
rect 371878 261576 371884 261588
rect 88208 261548 371884 261576
rect 88208 261536 88214 261548
rect 371878 261536 371884 261548
rect 371936 261536 371942 261588
rect 110322 261468 110328 261520
rect 110380 261508 110386 261520
rect 400858 261508 400864 261520
rect 110380 261480 400864 261508
rect 110380 261468 110386 261480
rect 400858 261468 400864 261480
rect 400916 261468 400922 261520
rect 17218 261400 17224 261452
rect 17276 261440 17282 261452
rect 139394 261440 139400 261452
rect 17276 261412 139400 261440
rect 17276 261400 17282 261412
rect 139394 261400 139400 261412
rect 139452 261400 139458 261452
rect 161382 261400 161388 261452
rect 161440 261440 161446 261452
rect 228818 261440 228824 261452
rect 161440 261412 228824 261440
rect 161440 261400 161446 261412
rect 228818 261400 228824 261412
rect 228876 261400 228882 261452
rect 238202 261400 238208 261452
rect 238260 261440 238266 261452
rect 270586 261440 270592 261452
rect 238260 261412 270592 261440
rect 238260 261400 238266 261412
rect 270586 261400 270592 261412
rect 270644 261400 270650 261452
rect 22738 261332 22744 261384
rect 22796 261372 22802 261384
rect 135346 261372 135352 261384
rect 22796 261344 135352 261372
rect 22796 261332 22802 261344
rect 135346 261332 135352 261344
rect 135404 261332 135410 261384
rect 186222 261332 186228 261384
rect 186280 261372 186286 261384
rect 226978 261372 226984 261384
rect 186280 261344 226984 261372
rect 186280 261332 186286 261344
rect 226978 261332 226984 261344
rect 227036 261332 227042 261384
rect 240870 261332 240876 261384
rect 240928 261372 240934 261384
rect 266354 261372 266360 261384
rect 240928 261344 266360 261372
rect 240928 261332 240934 261344
rect 266354 261332 266360 261344
rect 266412 261332 266418 261384
rect 117130 261264 117136 261316
rect 117188 261304 117194 261316
rect 226058 261304 226064 261316
rect 117188 261276 226064 261304
rect 117188 261264 117194 261276
rect 226058 261264 226064 261276
rect 226116 261264 226122 261316
rect 104618 261196 104624 261248
rect 104676 261236 104682 261248
rect 209038 261236 209044 261248
rect 104676 261208 209044 261236
rect 104676 261196 104682 261208
rect 209038 261196 209044 261208
rect 209096 261196 209102 261248
rect 55858 261128 55864 261180
rect 55916 261168 55922 261180
rect 155954 261168 155960 261180
rect 55916 261140 155960 261168
rect 55916 261128 55922 261140
rect 155954 261128 155960 261140
rect 156012 261128 156018 261180
rect 117130 261060 117136 261112
rect 117188 261100 117194 261112
rect 204898 261100 204904 261112
rect 117188 261072 204904 261100
rect 117188 261060 117194 261072
rect 204898 261060 204904 261072
rect 204956 261060 204962 261112
rect 41322 260992 41328 261044
rect 41380 261032 41386 261044
rect 128446 261032 128452 261044
rect 41380 261004 128452 261032
rect 41380 260992 41386 261004
rect 128446 260992 128452 261004
rect 128504 260992 128510 261044
rect 121270 260924 121276 260976
rect 121328 260964 121334 260976
rect 201494 260964 201500 260976
rect 121328 260936 201500 260964
rect 121328 260924 121334 260936
rect 201494 260924 201500 260936
rect 201552 260924 201558 260976
rect 114462 260788 114468 260840
rect 114520 260828 114526 260840
rect 214558 260828 214564 260840
rect 114520 260800 214564 260828
rect 114520 260788 114526 260800
rect 214558 260788 214564 260800
rect 214616 260788 214622 260840
rect 101950 260720 101956 260772
rect 102008 260760 102014 260772
rect 206370 260760 206376 260772
rect 102008 260732 206376 260760
rect 102008 260720 102014 260732
rect 206370 260720 206376 260732
rect 206428 260720 206434 260772
rect 121362 260652 121368 260704
rect 121420 260692 121426 260704
rect 226150 260692 226156 260704
rect 121420 260664 226156 260692
rect 121420 260652 121426 260664
rect 226150 260652 226156 260664
rect 226208 260652 226214 260704
rect 25498 260584 25504 260636
rect 25556 260624 25562 260636
rect 138106 260624 138112 260636
rect 25556 260596 138112 260624
rect 25556 260584 25562 260596
rect 138106 260584 138112 260596
rect 138164 260584 138170 260636
rect 166902 260584 166908 260636
rect 166960 260624 166966 260636
rect 228910 260624 228916 260636
rect 166960 260596 228916 260624
rect 166960 260584 166966 260596
rect 228910 260584 228916 260596
rect 228968 260584 228974 260636
rect 15838 260516 15844 260568
rect 15896 260556 15902 260568
rect 131114 260556 131120 260568
rect 15896 260528 131120 260556
rect 15896 260516 15902 260528
rect 131114 260516 131120 260528
rect 131172 260516 131178 260568
rect 200022 260516 200028 260568
rect 200080 260556 200086 260568
rect 282178 260556 282184 260568
rect 200080 260528 282184 260556
rect 200080 260516 200086 260528
rect 282178 260516 282184 260528
rect 282236 260516 282242 260568
rect 4798 260448 4804 260500
rect 4856 260488 4862 260500
rect 131206 260488 131212 260500
rect 4856 260460 131212 260488
rect 4856 260448 4862 260460
rect 131206 260448 131212 260460
rect 131264 260448 131270 260500
rect 218606 260448 218612 260500
rect 218664 260488 218670 260500
rect 304258 260488 304264 260500
rect 218664 260460 304264 260488
rect 218664 260448 218670 260460
rect 304258 260448 304264 260460
rect 304316 260448 304322 260500
rect 89622 260380 89628 260432
rect 89680 260420 89686 260432
rect 225230 260420 225236 260432
rect 89680 260392 225236 260420
rect 89680 260380 89686 260392
rect 225230 260380 225236 260392
rect 225288 260380 225294 260432
rect 231302 260380 231308 260432
rect 231360 260420 231366 260432
rect 320174 260420 320180 260432
rect 231360 260392 320180 260420
rect 231360 260380 231366 260392
rect 320174 260380 320180 260392
rect 320232 260380 320238 260432
rect 93762 260312 93768 260364
rect 93820 260352 93826 260364
rect 360838 260352 360844 260364
rect 93820 260324 360844 260352
rect 93820 260312 93826 260324
rect 360838 260312 360844 260324
rect 360896 260312 360902 260364
rect 96522 260244 96528 260296
rect 96580 260284 96586 260296
rect 363598 260284 363604 260296
rect 96580 260256 363604 260284
rect 96580 260244 96586 260256
rect 363598 260244 363604 260256
rect 363656 260244 363662 260296
rect 56134 260176 56140 260228
rect 56192 260216 56198 260228
rect 89714 260216 89720 260228
rect 56192 260188 89720 260216
rect 56192 260176 56198 260188
rect 89714 260176 89720 260188
rect 89772 260176 89778 260228
rect 90910 260176 90916 260228
rect 90968 260216 90974 260228
rect 358078 260216 358084 260228
rect 90968 260188 358084 260216
rect 90968 260176 90974 260188
rect 358078 260176 358084 260188
rect 358136 260176 358142 260228
rect 53282 260108 53288 260160
rect 53340 260148 53346 260160
rect 358906 260148 358912 260160
rect 53340 260120 358912 260148
rect 53340 260108 53346 260120
rect 358906 260108 358912 260120
rect 358964 260108 358970 260160
rect 118418 260040 118424 260092
rect 118476 260080 118482 260092
rect 206278 260080 206284 260092
rect 118476 260052 206284 260080
rect 118476 260040 118482 260052
rect 206278 260040 206284 260052
rect 206336 260040 206342 260092
rect 281994 245556 282000 245608
rect 282052 245596 282058 245608
rect 580166 245596 580172 245608
rect 282052 245568 580172 245596
rect 282052 245556 282058 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 54570 225360 54576 225412
rect 54628 225400 54634 225412
rect 57238 225400 57244 225412
rect 54628 225372 57244 225400
rect 54628 225360 54634 225372
rect 57238 225360 57244 225372
rect 57296 225360 57302 225412
rect 2774 215228 2780 215280
rect 2832 215268 2838 215280
rect 4798 215268 4804 215280
rect 2832 215240 4804 215268
rect 2832 215228 2838 215240
rect 4798 215228 4804 215240
rect 4856 215228 4862 215280
rect 54662 195916 54668 195968
rect 54720 195956 54726 195968
rect 57514 195956 57520 195968
rect 54720 195928 57520 195956
rect 54720 195916 54726 195928
rect 57514 195916 57520 195928
rect 57572 195916 57578 195968
rect 53374 192652 53380 192704
rect 53432 192692 53438 192704
rect 57514 192692 57520 192704
rect 53432 192664 57520 192692
rect 53432 192652 53438 192664
rect 57514 192652 57520 192664
rect 57572 192652 57578 192704
rect 3142 188980 3148 189032
rect 3200 189020 3206 189032
rect 17218 189020 17224 189032
rect 3200 188992 17224 189020
rect 3200 188980 3206 188992
rect 17218 188980 17224 188992
rect 17276 188980 17282 189032
rect 54938 187620 54944 187672
rect 54996 187660 55002 187672
rect 57238 187660 57244 187672
rect 54996 187632 57244 187660
rect 54996 187620 55002 187632
rect 57238 187620 57244 187632
rect 57296 187620 57302 187672
rect 54294 182792 54300 182844
rect 54352 182832 54358 182844
rect 57514 182832 57520 182844
rect 54352 182804 57520 182832
rect 54352 182792 54358 182804
rect 57514 182792 57520 182804
rect 57572 182792 57578 182844
rect 57514 175584 57520 175636
rect 57572 175624 57578 175636
rect 59814 175624 59820 175636
rect 57572 175596 59820 175624
rect 57572 175584 57578 175596
rect 59814 175584 59820 175596
rect 59872 175584 59878 175636
rect 57422 175176 57428 175228
rect 57480 175216 57486 175228
rect 58894 175216 58900 175228
rect 57480 175188 58900 175216
rect 57480 175176 57486 175188
rect 58894 175176 58900 175188
rect 58952 175176 58958 175228
rect 54386 169668 54392 169720
rect 54444 169708 54450 169720
rect 57790 169708 57796 169720
rect 54444 169680 57796 169708
rect 54444 169668 54450 169680
rect 57790 169668 57796 169680
rect 57848 169668 57854 169720
rect 3326 162936 3332 162988
rect 3384 162976 3390 162988
rect 7558 162976 7564 162988
rect 3384 162948 7564 162976
rect 3384 162936 3390 162948
rect 7558 162936 7564 162948
rect 7616 162936 7622 162988
rect 55030 162800 55036 162852
rect 55088 162840 55094 162852
rect 57422 162840 57428 162852
rect 55088 162812 57428 162840
rect 55088 162800 55094 162812
rect 57422 162800 57428 162812
rect 57480 162800 57486 162852
rect 54754 160012 54760 160064
rect 54812 160052 54818 160064
rect 57790 160052 57796 160064
rect 54812 160024 57796 160052
rect 54812 160012 54818 160024
rect 57790 160012 57796 160024
rect 57848 160012 57854 160064
rect 51994 157292 52000 157344
rect 52052 157332 52058 157344
rect 57422 157332 57428 157344
rect 52052 157304 57428 157332
rect 52052 157292 52058 157304
rect 57422 157292 57428 157304
rect 57480 157292 57486 157344
rect 52086 153824 52092 153876
rect 52144 153864 52150 153876
rect 57422 153864 57428 153876
rect 52144 153836 57428 153864
rect 52144 153824 52150 153836
rect 57422 153824 57428 153836
rect 57480 153824 57486 153876
rect 396718 153144 396724 153196
rect 396776 153184 396782 153196
rect 579614 153184 579620 153196
rect 396776 153156 579620 153184
rect 396776 153144 396782 153156
rect 579614 153144 579620 153156
rect 579672 153144 579678 153196
rect 54478 151716 54484 151768
rect 54536 151756 54542 151768
rect 57422 151756 57428 151768
rect 54536 151728 57428 151756
rect 54536 151716 54542 151728
rect 57422 151716 57428 151728
rect 57480 151716 57486 151768
rect 53558 144576 53564 144628
rect 53616 144616 53622 144628
rect 57422 144616 57428 144628
rect 53616 144588 57428 144616
rect 53616 144576 53622 144588
rect 57422 144576 57428 144588
rect 57480 144576 57486 144628
rect 53650 142060 53656 142112
rect 53708 142100 53714 142112
rect 57790 142100 57796 142112
rect 53708 142072 57796 142100
rect 53708 142060 53714 142072
rect 57790 142060 57796 142072
rect 57848 142060 57854 142112
rect 3326 137912 3332 137964
rect 3384 137952 3390 137964
rect 18598 137952 18604 137964
rect 3384 137924 18604 137952
rect 3384 137912 3390 137924
rect 18598 137912 18604 137924
rect 18656 137912 18662 137964
rect 57606 137436 57612 137488
rect 57664 137476 57670 137488
rect 57790 137476 57796 137488
rect 57664 137448 57796 137476
rect 57664 137436 57670 137448
rect 57790 137436 57796 137448
rect 57848 137436 57854 137488
rect 53742 136552 53748 136604
rect 53800 136592 53806 136604
rect 57606 136592 57612 136604
rect 53800 136564 57612 136592
rect 53800 136552 53806 136564
rect 57606 136552 57612 136564
rect 57664 136552 57670 136604
rect 55122 126896 55128 126948
rect 55180 126936 55186 126948
rect 57606 126936 57612 126948
rect 55180 126908 57612 126936
rect 55180 126896 55186 126908
rect 57606 126896 57612 126908
rect 57664 126896 57670 126948
rect 260098 126896 260104 126948
rect 260156 126936 260162 126948
rect 580166 126936 580172 126948
rect 260156 126908 580172 126936
rect 260156 126896 260162 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 53190 121388 53196 121440
rect 53248 121428 53254 121440
rect 57606 121428 57612 121440
rect 53248 121400 57612 121428
rect 53248 121388 53254 121400
rect 57606 121388 57612 121400
rect 57664 121388 57670 121440
rect 52178 113092 52184 113144
rect 52236 113132 52242 113144
rect 57606 113132 57612 113144
rect 52236 113104 57612 113132
rect 52236 113092 52242 113104
rect 57606 113092 57612 113104
rect 57664 113092 57670 113144
rect 3142 111732 3148 111784
rect 3200 111772 3206 111784
rect 11698 111772 11704 111784
rect 3200 111744 11704 111772
rect 3200 111732 3206 111744
rect 11698 111732 11704 111744
rect 11756 111732 11762 111784
rect 56502 108332 56508 108384
rect 56560 108372 56566 108384
rect 57238 108372 57244 108384
rect 56560 108344 57244 108372
rect 56560 108332 56566 108344
rect 57238 108332 57244 108344
rect 57296 108332 57302 108384
rect 53466 105544 53472 105596
rect 53524 105584 53530 105596
rect 57606 105584 57612 105596
rect 53524 105556 57612 105584
rect 53524 105544 53530 105556
rect 57606 105544 57612 105556
rect 57664 105544 57670 105596
rect 54846 103436 54852 103488
rect 54904 103476 54910 103488
rect 57606 103476 57612 103488
rect 54904 103448 57612 103476
rect 54904 103436 54910 103448
rect 57606 103436 57612 103448
rect 57664 103436 57670 103488
rect 54570 100648 54576 100700
rect 54628 100688 54634 100700
rect 57606 100688 57612 100700
rect 54628 100660 57612 100688
rect 54628 100648 54634 100660
rect 57606 100648 57612 100660
rect 57664 100648 57670 100700
rect 3234 97928 3240 97980
rect 3292 97968 3298 97980
rect 25498 97968 25504 97980
rect 3292 97940 25504 97968
rect 3292 97928 3298 97940
rect 25498 97928 25504 97940
rect 25556 97928 25562 97980
rect 52270 88272 52276 88324
rect 52328 88312 52334 88324
rect 57606 88312 57612 88324
rect 52328 88284 57612 88312
rect 52328 88272 52334 88284
rect 57606 88272 57612 88284
rect 57664 88272 57670 88324
rect 3326 85484 3332 85536
rect 3384 85524 3390 85536
rect 21358 85524 21364 85536
rect 3384 85496 21364 85524
rect 3384 85484 3390 85496
rect 21358 85484 21364 85496
rect 21416 85484 21422 85536
rect 53282 82764 53288 82816
rect 53340 82804 53346 82816
rect 57238 82804 57244 82816
rect 53340 82776 57244 82804
rect 53340 82764 53346 82776
rect 57238 82764 57244 82776
rect 57296 82764 57302 82816
rect 3326 71680 3332 71732
rect 3384 71720 3390 71732
rect 14458 71720 14464 71732
rect 3384 71692 14464 71720
rect 3384 71680 3390 71692
rect 14458 71680 14464 71692
rect 14516 71680 14522 71732
rect 52362 70320 52368 70372
rect 52420 70360 52426 70372
rect 57606 70360 57612 70372
rect 52420 70332 57612 70360
rect 52420 70320 52426 70332
rect 57606 70320 57612 70332
rect 57664 70320 57670 70372
rect 580166 59956 580172 59968
rect 209746 59928 239444 59956
rect 208118 59848 208124 59900
rect 208176 59888 208182 59900
rect 209746 59888 209774 59928
rect 208176 59860 209774 59888
rect 208176 59848 208182 59860
rect 223850 59848 223856 59900
rect 223908 59888 223914 59900
rect 225414 59888 225420 59900
rect 223908 59860 225420 59888
rect 223908 59848 223914 59860
rect 225414 59848 225420 59860
rect 225472 59848 225478 59900
rect 226058 59848 226064 59900
rect 226116 59888 226122 59900
rect 239416 59888 239444 59928
rect 240704 59928 580172 59956
rect 240704 59900 240732 59928
rect 580166 59916 580172 59928
rect 580224 59916 580230 59968
rect 240134 59888 240140 59900
rect 226116 59860 238892 59888
rect 239416 59860 240140 59888
rect 226116 59848 226122 59860
rect 214558 59780 214564 59832
rect 214616 59820 214622 59832
rect 214616 59792 238800 59820
rect 214616 59780 214622 59792
rect 218054 59712 218060 59764
rect 218112 59752 218118 59764
rect 218112 59724 238156 59752
rect 218112 59712 218118 59724
rect 212442 59644 212448 59696
rect 212500 59684 212506 59696
rect 212500 59656 233188 59684
rect 212500 59644 212506 59656
rect 213822 59576 213828 59628
rect 213880 59616 213886 59628
rect 232222 59616 232228 59628
rect 213880 59588 232228 59616
rect 213880 59576 213886 59588
rect 232222 59576 232228 59588
rect 232280 59576 232286 59628
rect 224126 59508 224132 59560
rect 224184 59548 224190 59560
rect 226058 59548 226064 59560
rect 224184 59520 226064 59548
rect 224184 59508 224190 59520
rect 226058 59508 226064 59520
rect 226116 59508 226122 59560
rect 233160 59548 233188 59656
rect 233326 59576 233332 59628
rect 233384 59616 233390 59628
rect 238018 59616 238024 59628
rect 233384 59588 238024 59616
rect 233384 59576 233390 59588
rect 238018 59576 238024 59588
rect 238076 59576 238082 59628
rect 238128 59616 238156 59724
rect 238772 59684 238800 59792
rect 238864 59752 238892 59860
rect 240134 59848 240140 59860
rect 240192 59848 240198 59900
rect 240686 59848 240692 59900
rect 240744 59848 240750 59900
rect 267826 59888 267832 59900
rect 241072 59860 267832 59888
rect 241072 59752 241100 59860
rect 267826 59848 267832 59860
rect 267884 59848 267890 59900
rect 251174 59820 251180 59832
rect 238864 59724 241100 59752
rect 248386 59792 251180 59820
rect 248386 59684 248414 59792
rect 251174 59780 251180 59792
rect 251232 59780 251238 59832
rect 238772 59656 248414 59684
rect 245654 59616 245660 59628
rect 238128 59588 245660 59616
rect 245654 59576 245660 59588
rect 245712 59576 245718 59628
rect 237374 59548 237380 59560
rect 233160 59520 237380 59548
rect 237374 59508 237380 59520
rect 237432 59508 237438 59560
rect 207290 59440 207296 59492
rect 207348 59480 207354 59492
rect 207348 59452 232360 59480
rect 207348 59440 207354 59452
rect 205542 59372 205548 59424
rect 205600 59412 205606 59424
rect 212442 59412 212448 59424
rect 205600 59384 212448 59412
rect 205600 59372 205606 59384
rect 212442 59372 212448 59384
rect 212500 59372 212506 59424
rect 223942 59372 223948 59424
rect 224000 59412 224006 59424
rect 232222 59412 232228 59424
rect 224000 59384 232228 59412
rect 224000 59372 224006 59384
rect 232222 59372 232228 59384
rect 232280 59372 232286 59424
rect 56686 59304 56692 59356
rect 56744 59344 56750 59356
rect 212902 59344 212908 59356
rect 56744 59316 212908 59344
rect 56744 59304 56750 59316
rect 212902 59304 212908 59316
rect 212960 59304 212966 59356
rect 216950 59304 216956 59356
rect 217008 59344 217014 59356
rect 224770 59344 224776 59356
rect 217008 59316 224776 59344
rect 217008 59304 217014 59316
rect 224770 59304 224776 59316
rect 224828 59304 224834 59356
rect 232332 59344 232360 59452
rect 232406 59440 232412 59492
rect 232464 59480 232470 59492
rect 235994 59480 236000 59492
rect 232464 59452 236000 59480
rect 232464 59440 232470 59452
rect 235994 59440 236000 59452
rect 236052 59440 236058 59492
rect 232498 59372 232504 59424
rect 232556 59412 232562 59424
rect 322934 59412 322940 59424
rect 232556 59384 322940 59412
rect 232556 59372 232562 59384
rect 322934 59372 322940 59384
rect 322992 59372 322998 59424
rect 233326 59344 233332 59356
rect 232332 59316 233332 59344
rect 233326 59304 233332 59316
rect 233384 59304 233390 59356
rect 56594 59236 56600 59288
rect 56652 59276 56658 59288
rect 203794 59276 203800 59288
rect 56652 59248 203800 59276
rect 56652 59236 56658 59248
rect 203794 59236 203800 59248
rect 203852 59236 203858 59288
rect 215754 59236 215760 59288
rect 215812 59276 215818 59288
rect 215812 59248 220952 59276
rect 215812 59236 215818 59248
rect 218422 59168 218428 59220
rect 218480 59208 218486 59220
rect 220924 59208 220952 59248
rect 220998 59236 221004 59288
rect 221056 59276 221062 59288
rect 267734 59276 267740 59288
rect 221056 59248 267740 59276
rect 221056 59236 221062 59248
rect 267734 59236 267740 59248
rect 267792 59236 267798 59288
rect 224954 59208 224960 59220
rect 218480 59180 219434 59208
rect 220924 59180 224960 59208
rect 218480 59168 218486 59180
rect 219406 59140 219434 59180
rect 224954 59168 224960 59180
rect 225012 59168 225018 59220
rect 262214 59140 262220 59152
rect 219406 59112 262220 59140
rect 262214 59100 262220 59112
rect 262272 59100 262278 59152
rect 223390 59032 223396 59084
rect 223448 59072 223454 59084
rect 225230 59072 225236 59084
rect 223448 59044 225236 59072
rect 223448 59032 223454 59044
rect 225230 59032 225236 59044
rect 225288 59032 225294 59084
rect 207566 58964 207572 59016
rect 207624 59004 207630 59016
rect 227990 59004 227996 59016
rect 207624 58976 227996 59004
rect 207624 58964 207630 58976
rect 227990 58964 227996 58976
rect 228048 58964 228054 59016
rect 208210 58896 208216 58948
rect 208268 58936 208274 58948
rect 227898 58936 227904 58948
rect 208268 58908 227904 58936
rect 208268 58896 208274 58908
rect 227898 58896 227904 58908
rect 227956 58896 227962 58948
rect 209314 58828 209320 58880
rect 209372 58868 209378 58880
rect 222470 58868 222476 58880
rect 209372 58840 222476 58868
rect 209372 58828 209378 58840
rect 222470 58828 222476 58840
rect 222528 58828 222534 58880
rect 223758 58828 223764 58880
rect 223816 58868 223822 58880
rect 228082 58868 228088 58880
rect 223816 58840 228088 58868
rect 223816 58828 223822 58840
rect 228082 58828 228088 58840
rect 228140 58828 228146 58880
rect 216398 58760 216404 58812
rect 216456 58800 216462 58812
rect 229186 58800 229192 58812
rect 216456 58772 229192 58800
rect 216456 58760 216462 58772
rect 229186 58760 229192 58772
rect 229244 58760 229250 58812
rect 216674 58692 216680 58744
rect 216732 58732 216738 58744
rect 224218 58732 224224 58744
rect 216732 58704 224224 58732
rect 216732 58692 216738 58704
rect 224218 58692 224224 58704
rect 224276 58692 224282 58744
rect 224402 58692 224408 58744
rect 224460 58732 224466 58744
rect 228266 58732 228272 58744
rect 224460 58704 228272 58732
rect 224460 58692 224466 58704
rect 228266 58692 228272 58704
rect 228324 58692 228330 58744
rect 211982 58624 211988 58676
rect 212040 58664 212046 58676
rect 264238 58664 264244 58676
rect 212040 58636 264244 58664
rect 212040 58624 212046 58636
rect 264238 58624 264244 58636
rect 264296 58624 264302 58676
rect 214926 58556 214932 58608
rect 214984 58596 214990 58608
rect 214984 58568 219572 58596
rect 214984 58556 214990 58568
rect 140222 58488 140228 58540
rect 140280 58528 140286 58540
rect 140682 58528 140688 58540
rect 140280 58500 140688 58528
rect 140280 58488 140286 58500
rect 140682 58488 140688 58500
rect 140740 58488 140746 58540
rect 217778 58488 217784 58540
rect 217836 58528 217842 58540
rect 219434 58528 219440 58540
rect 217836 58500 219440 58528
rect 217836 58488 217842 58500
rect 219434 58488 219440 58500
rect 219492 58488 219498 58540
rect 219544 58528 219572 58568
rect 222286 58556 222292 58608
rect 222344 58596 222350 58608
rect 258718 58596 258724 58608
rect 222344 58568 258724 58596
rect 222344 58556 222350 58568
rect 258718 58556 258724 58568
rect 258776 58556 258782 58608
rect 224862 58528 224868 58540
rect 219544 58500 224868 58528
rect 224862 58488 224868 58500
rect 224920 58488 224926 58540
rect 210786 58420 210792 58472
rect 210844 58460 210850 58472
rect 222378 58460 222384 58472
rect 210844 58432 222384 58460
rect 210844 58420 210850 58432
rect 222378 58420 222384 58432
rect 222436 58420 222442 58472
rect 222470 58420 222476 58472
rect 222528 58460 222534 58472
rect 229094 58460 229100 58472
rect 222528 58432 229100 58460
rect 222528 58420 222534 58432
rect 229094 58420 229100 58432
rect 229152 58420 229158 58472
rect 217502 58352 217508 58404
rect 217560 58392 217566 58404
rect 249058 58392 249064 58404
rect 217560 58364 249064 58392
rect 217560 58352 217566 58364
rect 249058 58352 249064 58364
rect 249116 58352 249122 58404
rect 212534 58284 212540 58336
rect 212592 58324 212598 58336
rect 222286 58324 222292 58336
rect 212592 58296 222292 58324
rect 212592 58284 212598 58296
rect 222286 58284 222292 58296
rect 222344 58284 222350 58336
rect 222378 58284 222384 58336
rect 222436 58324 222442 58336
rect 228174 58324 228180 58336
rect 222436 58296 228180 58324
rect 222436 58284 222442 58296
rect 228174 58284 228180 58296
rect 228232 58284 228238 58336
rect 205818 58216 205824 58268
rect 205876 58256 205882 58268
rect 223758 58256 223764 58268
rect 205876 58228 223764 58256
rect 205876 58216 205882 58228
rect 223758 58216 223764 58228
rect 223816 58216 223822 58268
rect 224218 58216 224224 58268
rect 224276 58256 224282 58268
rect 230474 58256 230480 58268
rect 224276 58228 230480 58256
rect 224276 58216 224282 58228
rect 230474 58216 230480 58228
rect 230532 58216 230538 58268
rect 214006 58148 214012 58200
rect 214064 58188 214070 58200
rect 221826 58188 221832 58200
rect 214064 58160 221832 58188
rect 214064 58148 214070 58160
rect 221826 58148 221832 58160
rect 221884 58148 221890 58200
rect 221918 58148 221924 58200
rect 221976 58188 221982 58200
rect 231946 58188 231952 58200
rect 221976 58160 231952 58188
rect 221976 58148 221982 58160
rect 231946 58148 231952 58160
rect 232004 58148 232010 58200
rect 162210 58120 162216 58132
rect 159836 58092 162216 58120
rect 64616 58024 65196 58052
rect 59262 57944 59268 57996
rect 59320 57984 59326 57996
rect 61286 57984 61292 57996
rect 59320 57956 61292 57984
rect 59320 57944 59326 57956
rect 61286 57944 61292 57956
rect 61344 57944 61350 57996
rect 45462 57876 45468 57928
rect 45520 57916 45526 57928
rect 64616 57916 64644 58024
rect 64690 57944 64696 57996
rect 64748 57984 64754 57996
rect 64748 57956 65104 57984
rect 64748 57944 64754 57956
rect 45520 57888 64644 57916
rect 45520 57876 45526 57888
rect 41322 57808 41328 57860
rect 41380 57848 41386 57860
rect 64874 57848 64880 57860
rect 41380 57820 64880 57848
rect 41380 57808 41386 57820
rect 64874 57808 64880 57820
rect 64932 57808 64938 57860
rect 65076 57848 65104 57956
rect 65168 57916 65196 58024
rect 143166 58012 143172 58064
rect 143224 58052 143230 58064
rect 149422 58052 149428 58064
rect 143224 58024 149428 58052
rect 143224 58012 143230 58024
rect 149422 58012 149428 58024
rect 149480 58012 149486 58064
rect 102134 57984 102140 57996
rect 100496 57956 102140 57984
rect 65168 57888 70394 57916
rect 65076 57820 68600 57848
rect 35802 57740 35808 57792
rect 35860 57780 35866 57792
rect 68462 57780 68468 57792
rect 35860 57752 68468 57780
rect 35860 57740 35866 57752
rect 68462 57740 68468 57752
rect 68520 57740 68526 57792
rect 39942 57672 39948 57724
rect 40000 57712 40006 57724
rect 61930 57712 61936 57724
rect 40000 57684 61936 57712
rect 40000 57672 40006 57684
rect 61930 57672 61936 57684
rect 61988 57672 61994 57724
rect 67910 57712 67916 57724
rect 62132 57684 67916 57712
rect 34422 57604 34428 57656
rect 34480 57644 34486 57656
rect 62022 57644 62028 57656
rect 34480 57616 62028 57644
rect 34480 57604 34486 57616
rect 62022 57604 62028 57616
rect 62080 57604 62086 57656
rect 33042 57536 33048 57588
rect 33100 57576 33106 57588
rect 62132 57576 62160 57684
rect 67910 57672 67916 57684
rect 67968 57672 67974 57724
rect 68572 57712 68600 57820
rect 70366 57780 70394 57888
rect 84562 57876 84568 57928
rect 84620 57916 84626 57928
rect 92842 57916 92848 57928
rect 84620 57888 92848 57916
rect 84620 57876 84626 57888
rect 92842 57876 92848 57888
rect 92900 57876 92906 57928
rect 95050 57876 95056 57928
rect 95108 57916 95114 57928
rect 100496 57916 100524 57956
rect 102134 57944 102140 57956
rect 102192 57944 102198 57996
rect 120350 57944 120356 57996
rect 120408 57984 120414 57996
rect 128170 57984 128176 57996
rect 120408 57956 128176 57984
rect 120408 57944 120414 57956
rect 128170 57944 128176 57956
rect 128228 57944 128234 57996
rect 132862 57944 132868 57996
rect 132920 57984 132926 57996
rect 140958 57984 140964 57996
rect 132920 57956 140964 57984
rect 132920 57944 132926 57956
rect 140958 57944 140964 57956
rect 141016 57944 141022 57996
rect 143258 57944 143264 57996
rect 143316 57984 143322 57996
rect 143442 57984 143448 57996
rect 143316 57956 143448 57984
rect 143316 57944 143322 57956
rect 143442 57944 143448 57956
rect 143500 57944 143506 57996
rect 159836 57984 159864 58092
rect 162210 58080 162216 58092
rect 162268 58080 162274 58132
rect 172146 58080 172152 58132
rect 172204 58120 172210 58132
rect 179230 58120 179236 58132
rect 172204 58092 179236 58120
rect 172204 58080 172210 58092
rect 179230 58080 179236 58092
rect 179288 58080 179294 58132
rect 204990 58080 204996 58132
rect 205048 58120 205054 58132
rect 205048 58092 219434 58120
rect 205048 58080 205054 58092
rect 175292 58024 175596 58052
rect 159744 57956 159864 57984
rect 168484 57956 169984 57984
rect 95108 57888 100524 57916
rect 95108 57876 95114 57888
rect 100570 57876 100576 57928
rect 100628 57916 100634 57928
rect 159744 57916 159772 57956
rect 100628 57888 159772 57916
rect 100628 57876 100634 57888
rect 159818 57876 159824 57928
rect 159876 57916 159882 57928
rect 165798 57916 165804 57928
rect 159876 57888 165804 57916
rect 159876 57876 159882 57888
rect 165798 57876 165804 57888
rect 165856 57876 165862 57928
rect 165890 57876 165896 57928
rect 165948 57916 165954 57928
rect 168484 57916 168512 57956
rect 165948 57888 168512 57916
rect 165948 57876 165954 57888
rect 168558 57876 168564 57928
rect 168616 57916 168622 57928
rect 169956 57916 169984 57956
rect 175292 57916 175320 58024
rect 168616 57888 169892 57916
rect 169956 57888 175320 57916
rect 175568 57916 175596 58024
rect 219406 57984 219434 58092
rect 219526 58080 219532 58132
rect 219584 58120 219590 58132
rect 230566 58120 230572 58132
rect 219584 58092 230572 58120
rect 219584 58080 219590 58092
rect 230566 58080 230572 58092
rect 230624 58080 230630 58132
rect 219802 58012 219808 58064
rect 219860 58052 219866 58064
rect 231854 58052 231860 58064
rect 219860 58024 231860 58052
rect 219860 58012 219866 58024
rect 231854 58012 231860 58024
rect 231912 58012 231918 58064
rect 225046 57984 225052 57996
rect 219406 57956 225052 57984
rect 225046 57944 225052 57956
rect 225104 57944 225110 57996
rect 213178 57916 213184 57928
rect 175568 57888 213184 57916
rect 168616 57876 168622 57888
rect 85390 57808 85396 57860
rect 85448 57848 85454 57860
rect 85448 57820 93854 57848
rect 85448 57808 85454 57820
rect 70854 57780 70860 57792
rect 70366 57752 70860 57780
rect 70854 57740 70860 57752
rect 70912 57740 70918 57792
rect 80422 57740 80428 57792
rect 80480 57780 80486 57792
rect 82998 57780 83004 57792
rect 80480 57752 83004 57780
rect 80480 57740 80486 57752
rect 82998 57740 83004 57752
rect 83056 57740 83062 57792
rect 83734 57740 83740 57792
rect 83792 57780 83798 57792
rect 83918 57780 83924 57792
rect 83792 57752 83924 57780
rect 83792 57740 83798 57752
rect 83918 57740 83924 57752
rect 83976 57740 83982 57792
rect 86310 57740 86316 57792
rect 86368 57780 86374 57792
rect 86368 57752 92704 57780
rect 86368 57740 86374 57752
rect 68572 57684 70394 57712
rect 62206 57604 62212 57656
rect 62264 57644 62270 57656
rect 68186 57644 68192 57656
rect 62264 57616 68192 57644
rect 62264 57604 62270 57616
rect 68186 57604 68192 57616
rect 68244 57604 68250 57656
rect 70366 57644 70394 57684
rect 73062 57672 73068 57724
rect 73120 57712 73126 57724
rect 77846 57712 77852 57724
rect 73120 57684 77852 57712
rect 73120 57672 73126 57684
rect 77846 57672 77852 57684
rect 77904 57672 77910 57724
rect 81894 57672 81900 57724
rect 81952 57712 81958 57724
rect 87598 57712 87604 57724
rect 81952 57684 87604 57712
rect 81952 57672 81958 57684
rect 87598 57672 87604 57684
rect 87656 57672 87662 57724
rect 73706 57644 73712 57656
rect 70366 57616 73712 57644
rect 73706 57604 73712 57616
rect 73764 57604 73770 57656
rect 74718 57604 74724 57656
rect 74776 57644 74782 57656
rect 75270 57644 75276 57656
rect 74776 57616 75276 57644
rect 74776 57604 74782 57616
rect 75270 57604 75276 57616
rect 75328 57604 75334 57656
rect 76650 57604 76656 57656
rect 76708 57644 76714 57656
rect 78398 57644 78404 57656
rect 76708 57616 78404 57644
rect 76708 57604 76714 57616
rect 78398 57604 78404 57616
rect 78456 57604 78462 57656
rect 81066 57604 81072 57656
rect 81124 57644 81130 57656
rect 81342 57644 81348 57656
rect 81124 57616 81348 57644
rect 81124 57604 81130 57616
rect 81342 57604 81348 57616
rect 81400 57604 81406 57656
rect 86586 57604 86592 57656
rect 86644 57644 86650 57656
rect 86862 57644 86868 57656
rect 86644 57616 86868 57644
rect 86644 57604 86650 57616
rect 86862 57604 86868 57616
rect 86920 57604 86926 57656
rect 87414 57604 87420 57656
rect 87472 57644 87478 57656
rect 88150 57644 88156 57656
rect 87472 57616 88156 57644
rect 87472 57604 87478 57616
rect 88150 57604 88156 57616
rect 88208 57604 88214 57656
rect 88610 57604 88616 57656
rect 88668 57644 88674 57656
rect 89346 57644 89352 57656
rect 88668 57616 89352 57644
rect 88668 57604 88674 57616
rect 89346 57604 89352 57616
rect 89404 57604 89410 57656
rect 91278 57604 91284 57656
rect 91336 57644 91342 57656
rect 92290 57644 92296 57656
rect 91336 57616 92296 57644
rect 91336 57604 91342 57616
rect 92290 57604 92296 57616
rect 92348 57604 92354 57656
rect 66714 57576 66720 57588
rect 33100 57548 62160 57576
rect 62224 57548 66720 57576
rect 33100 57536 33106 57548
rect 28902 57468 28908 57520
rect 28960 57508 28966 57520
rect 62224 57508 62252 57548
rect 66714 57536 66720 57548
rect 66772 57536 66778 57588
rect 66898 57536 66904 57588
rect 66956 57576 66962 57588
rect 70210 57576 70216 57588
rect 66956 57548 70216 57576
rect 66956 57536 66962 57548
rect 70210 57536 70216 57548
rect 70268 57536 70274 57588
rect 71682 57536 71688 57588
rect 71740 57576 71746 57588
rect 77570 57576 77576 57588
rect 71740 57548 77576 57576
rect 71740 57536 71746 57548
rect 77570 57536 77576 57548
rect 77628 57536 77634 57588
rect 80146 57536 80152 57588
rect 80204 57576 80210 57588
rect 81250 57576 81256 57588
rect 80204 57548 81256 57576
rect 80204 57536 80210 57548
rect 81250 57536 81256 57548
rect 81308 57536 81314 57588
rect 83366 57536 83372 57588
rect 83424 57576 83430 57588
rect 84102 57576 84108 57588
rect 83424 57548 84108 57576
rect 83424 57536 83430 57548
rect 84102 57536 84108 57548
rect 84160 57536 84166 57588
rect 86034 57536 86040 57588
rect 86092 57576 86098 57588
rect 86678 57576 86684 57588
rect 86092 57548 86684 57576
rect 86092 57536 86098 57548
rect 86678 57536 86684 57548
rect 86736 57536 86742 57588
rect 88334 57536 88340 57588
rect 88392 57576 88398 57588
rect 89622 57576 89628 57588
rect 88392 57548 89628 57576
rect 88392 57536 88398 57548
rect 89622 57536 89628 57548
rect 89680 57536 89686 57588
rect 28960 57480 62252 57508
rect 28960 57468 28966 57480
rect 64874 57468 64880 57520
rect 64932 57508 64938 57520
rect 64932 57480 66116 57508
rect 64932 57468 64938 57480
rect 26142 57400 26148 57452
rect 26200 57440 26206 57452
rect 65978 57440 65984 57452
rect 26200 57412 65984 57440
rect 26200 57400 26206 57412
rect 65978 57400 65984 57412
rect 66036 57400 66042 57452
rect 66088 57440 66116 57480
rect 66162 57468 66168 57520
rect 66220 57508 66226 57520
rect 76098 57508 76104 57520
rect 66220 57480 76104 57508
rect 66220 57468 66226 57480
rect 76098 57468 76104 57480
rect 76156 57468 76162 57520
rect 77294 57508 77300 57520
rect 76208 57480 77300 57508
rect 69934 57440 69940 57452
rect 66088 57412 69940 57440
rect 69934 57400 69940 57412
rect 69992 57400 69998 57452
rect 70210 57400 70216 57452
rect 70268 57440 70274 57452
rect 76208 57440 76236 57480
rect 77294 57468 77300 57480
rect 77352 57468 77358 57520
rect 80790 57468 80796 57520
rect 80848 57508 80854 57520
rect 81342 57508 81348 57520
rect 80848 57480 81348 57508
rect 80848 57468 80854 57480
rect 81342 57468 81348 57480
rect 81400 57468 81406 57520
rect 82814 57468 82820 57520
rect 82872 57508 82878 57520
rect 83918 57508 83924 57520
rect 82872 57480 83924 57508
rect 82872 57468 82878 57480
rect 83918 57468 83924 57480
rect 83976 57468 83982 57520
rect 84286 57468 84292 57520
rect 84344 57508 84350 57520
rect 85390 57508 85396 57520
rect 84344 57480 85396 57508
rect 84344 57468 84350 57480
rect 85390 57468 85396 57480
rect 85448 57468 85454 57520
rect 85666 57468 85672 57520
rect 85724 57508 85730 57520
rect 86586 57508 86592 57520
rect 85724 57480 86592 57508
rect 85724 57468 85730 57480
rect 86586 57468 86592 57480
rect 86644 57468 86650 57520
rect 92676 57508 92704 57752
rect 92750 57604 92756 57656
rect 92808 57644 92814 57656
rect 93670 57644 93676 57656
rect 92808 57616 93676 57644
rect 92808 57604 92814 57616
rect 93670 57604 93676 57616
rect 93728 57604 93734 57656
rect 93826 57644 93854 57820
rect 94130 57808 94136 57860
rect 94188 57848 94194 57860
rect 96706 57848 96712 57860
rect 94188 57820 96712 57848
rect 94188 57808 94194 57820
rect 96706 57808 96712 57820
rect 96764 57808 96770 57860
rect 96798 57808 96804 57860
rect 96856 57848 96862 57860
rect 143166 57848 143172 57860
rect 96856 57820 143172 57848
rect 96856 57808 96862 57820
rect 143166 57808 143172 57820
rect 143224 57808 143230 57860
rect 143258 57808 143264 57860
rect 143316 57848 143322 57860
rect 148318 57848 148324 57860
rect 143316 57820 148324 57848
rect 143316 57808 143322 57820
rect 148318 57808 148324 57820
rect 148376 57808 148382 57860
rect 149238 57808 149244 57860
rect 149296 57848 149302 57860
rect 156782 57848 156788 57860
rect 149296 57820 156788 57848
rect 149296 57808 149302 57820
rect 156782 57808 156788 57820
rect 156840 57808 156846 57860
rect 156874 57808 156880 57860
rect 156932 57848 156938 57860
rect 157150 57848 157156 57860
rect 156932 57820 157156 57848
rect 156932 57808 156938 57820
rect 157150 57808 157156 57820
rect 157208 57808 157214 57860
rect 159174 57808 159180 57860
rect 159232 57848 159238 57860
rect 166810 57848 166816 57860
rect 159232 57820 166816 57848
rect 159232 57808 159238 57820
rect 166810 57808 166816 57820
rect 166868 57808 166874 57860
rect 166994 57808 167000 57860
rect 167052 57848 167058 57860
rect 168282 57848 168288 57860
rect 167052 57820 168288 57848
rect 167052 57808 167058 57820
rect 168282 57808 168288 57820
rect 168340 57808 168346 57860
rect 168834 57808 168840 57860
rect 168892 57848 168898 57860
rect 169570 57848 169576 57860
rect 168892 57820 169576 57848
rect 168892 57808 168898 57820
rect 169570 57808 169576 57820
rect 169628 57808 169634 57860
rect 169864 57848 169892 57888
rect 213178 57876 213184 57888
rect 213236 57876 213242 57928
rect 216030 57876 216036 57928
rect 216088 57916 216094 57928
rect 216088 57888 221228 57916
rect 216088 57876 216094 57888
rect 173710 57848 173716 57860
rect 169864 57820 173716 57848
rect 173710 57808 173716 57820
rect 173768 57808 173774 57860
rect 175550 57808 175556 57860
rect 175608 57848 175614 57860
rect 183002 57848 183008 57860
rect 175608 57820 183008 57848
rect 175608 57808 175614 57820
rect 183002 57808 183008 57820
rect 183060 57808 183066 57860
rect 183094 57808 183100 57860
rect 183152 57848 183158 57860
rect 183370 57848 183376 57860
rect 183152 57820 183376 57848
rect 183152 57808 183158 57820
rect 183370 57808 183376 57820
rect 183428 57808 183434 57860
rect 185118 57808 185124 57860
rect 185176 57848 185182 57860
rect 186038 57848 186044 57860
rect 185176 57820 186044 57848
rect 185176 57808 185182 57820
rect 186038 57808 186044 57820
rect 186096 57808 186102 57860
rect 186774 57808 186780 57860
rect 186832 57848 186838 57860
rect 187510 57848 187516 57860
rect 186832 57820 187516 57848
rect 186832 57808 186838 57820
rect 187510 57808 187516 57820
rect 187568 57808 187574 57860
rect 188062 57808 188068 57860
rect 188120 57848 188126 57860
rect 188890 57848 188896 57860
rect 188120 57820 188896 57848
rect 188120 57808 188126 57820
rect 188890 57808 188896 57820
rect 188948 57808 188954 57860
rect 189534 57808 189540 57860
rect 189592 57848 189598 57860
rect 190270 57848 190276 57860
rect 189592 57820 190276 57848
rect 189592 57808 189598 57820
rect 190270 57808 190276 57820
rect 190328 57808 190334 57860
rect 191282 57808 191288 57860
rect 191340 57848 191346 57860
rect 191558 57848 191564 57860
rect 191340 57820 191564 57848
rect 191340 57808 191346 57820
rect 191558 57808 191564 57820
rect 191616 57808 191622 57860
rect 192202 57808 192208 57860
rect 192260 57848 192266 57860
rect 193030 57848 193036 57860
rect 192260 57820 193036 57848
rect 192260 57808 192266 57820
rect 193030 57808 193036 57820
rect 193088 57808 193094 57860
rect 193214 57808 193220 57860
rect 193272 57848 193278 57860
rect 193858 57848 193864 57860
rect 193272 57820 193864 57848
rect 193272 57808 193278 57820
rect 193858 57808 193864 57820
rect 193916 57808 193922 57860
rect 195054 57808 195060 57860
rect 195112 57848 195118 57860
rect 195882 57848 195888 57860
rect 195112 57820 195888 57848
rect 195112 57808 195118 57820
rect 195882 57808 195888 57820
rect 195940 57808 195946 57860
rect 196250 57808 196256 57860
rect 196308 57848 196314 57860
rect 196986 57848 196992 57860
rect 196308 57820 196992 57848
rect 196308 57808 196314 57820
rect 196986 57808 196992 57820
rect 197044 57808 197050 57860
rect 197354 57808 197360 57860
rect 197412 57848 197418 57860
rect 198274 57848 198280 57860
rect 197412 57820 198280 57848
rect 197412 57808 197418 57820
rect 198274 57808 198280 57820
rect 198332 57808 198338 57860
rect 198826 57808 198832 57860
rect 198884 57848 198890 57860
rect 199838 57848 199844 57860
rect 198884 57820 199844 57848
rect 198884 57808 198890 57820
rect 199838 57808 199844 57820
rect 199896 57808 199902 57860
rect 201770 57808 201776 57860
rect 201828 57848 201834 57860
rect 202506 57848 202512 57860
rect 201828 57820 202512 57848
rect 201828 57808 201834 57820
rect 202506 57808 202512 57820
rect 202564 57808 202570 57860
rect 202966 57808 202972 57860
rect 203024 57848 203030 57860
rect 204162 57848 204168 57860
rect 203024 57820 204168 57848
rect 203024 57808 203030 57820
rect 204162 57808 204168 57820
rect 204220 57808 204226 57860
rect 208486 57808 208492 57860
rect 208544 57848 208550 57860
rect 218054 57848 218060 57860
rect 208544 57820 218060 57848
rect 208544 57808 208550 57820
rect 218054 57808 218060 57820
rect 218112 57808 218118 57860
rect 95878 57740 95884 57792
rect 95936 57780 95942 57792
rect 95936 57752 96568 57780
rect 95936 57740 95942 57752
rect 93826 57616 95556 57644
rect 92842 57536 92848 57588
rect 92900 57576 92906 57588
rect 94498 57576 94504 57588
rect 92900 57548 94504 57576
rect 92900 57536 92906 57548
rect 94498 57536 94504 57548
rect 94556 57536 94562 57588
rect 95528 57576 95556 57616
rect 95602 57604 95608 57656
rect 95660 57644 95666 57656
rect 96338 57644 96344 57656
rect 95660 57616 96344 57644
rect 95660 57604 95666 57616
rect 96338 57604 96344 57616
rect 96396 57604 96402 57656
rect 96540 57644 96568 57752
rect 97000 57752 101444 57780
rect 97000 57644 97028 57752
rect 101416 57712 101444 57752
rect 101490 57740 101496 57792
rect 101548 57780 101554 57792
rect 162026 57780 162032 57792
rect 101548 57752 162032 57780
rect 101548 57740 101554 57752
rect 162026 57740 162032 57752
rect 162084 57740 162090 57792
rect 162210 57740 162216 57792
rect 162268 57780 162274 57792
rect 164510 57780 164516 57792
rect 162268 57752 164516 57780
rect 162268 57740 162274 57752
rect 164510 57740 164516 57752
rect 164568 57740 164574 57792
rect 165890 57740 165896 57792
rect 165948 57780 165954 57792
rect 166902 57780 166908 57792
rect 165948 57752 166908 57780
rect 165948 57740 165954 57752
rect 166902 57740 166908 57752
rect 166960 57740 166966 57792
rect 167086 57740 167092 57792
rect 167144 57780 167150 57792
rect 168098 57780 168104 57792
rect 167144 57752 168104 57780
rect 167144 57740 167150 57752
rect 168098 57740 168104 57752
rect 168156 57740 168162 57792
rect 169386 57740 169392 57792
rect 169444 57780 169450 57792
rect 169662 57780 169668 57792
rect 169444 57752 169668 57780
rect 169444 57740 169450 57752
rect 169662 57740 169668 57752
rect 169720 57740 169726 57792
rect 169846 57740 169852 57792
rect 169904 57780 169910 57792
rect 170858 57780 170864 57792
rect 169904 57752 170864 57780
rect 169904 57740 169910 57752
rect 170858 57740 170864 57752
rect 170916 57740 170922 57792
rect 174170 57740 174176 57792
rect 174228 57780 174234 57792
rect 174228 57752 179184 57780
rect 174228 57740 174234 57752
rect 101582 57712 101588 57724
rect 101416 57684 101588 57712
rect 101582 57672 101588 57684
rect 101640 57672 101646 57724
rect 101766 57672 101772 57724
rect 101824 57712 101830 57724
rect 102042 57712 102048 57724
rect 101824 57684 102048 57712
rect 101824 57672 101830 57684
rect 102042 57672 102048 57684
rect 102100 57672 102106 57724
rect 102318 57672 102324 57724
rect 102376 57712 102382 57724
rect 171042 57712 171048 57724
rect 102376 57684 171048 57712
rect 102376 57672 102382 57684
rect 171042 57672 171048 57684
rect 171100 57672 171106 57724
rect 171134 57672 171140 57724
rect 171192 57712 171198 57724
rect 172146 57712 172152 57724
rect 171192 57684 172152 57712
rect 171192 57672 171198 57684
rect 172146 57672 172152 57684
rect 172204 57672 172210 57724
rect 172882 57672 172888 57724
rect 172940 57712 172946 57724
rect 173618 57712 173624 57724
rect 172940 57684 173624 57712
rect 172940 57672 172946 57684
rect 173618 57672 173624 57684
rect 173676 57672 173682 57724
rect 174078 57672 174084 57724
rect 174136 57712 174142 57724
rect 174998 57712 175004 57724
rect 174136 57684 175004 57712
rect 174136 57672 174142 57684
rect 174998 57672 175004 57684
rect 175056 57672 175062 57724
rect 176654 57672 176660 57724
rect 176712 57712 176718 57724
rect 177482 57712 177488 57724
rect 176712 57684 177488 57712
rect 176712 57672 176718 57684
rect 177482 57672 177488 57684
rect 177540 57672 177546 57724
rect 178126 57672 178132 57724
rect 178184 57712 178190 57724
rect 179046 57712 179052 57724
rect 178184 57684 179052 57712
rect 178184 57672 178190 57684
rect 179046 57672 179052 57684
rect 179104 57672 179110 57724
rect 179156 57712 179184 57752
rect 179230 57740 179236 57792
rect 179288 57780 179294 57792
rect 200482 57780 200488 57792
rect 179288 57752 200488 57780
rect 179288 57740 179294 57752
rect 200482 57740 200488 57752
rect 200540 57740 200546 57792
rect 200574 57740 200580 57792
rect 200632 57780 200638 57792
rect 201218 57780 201224 57792
rect 200632 57752 201224 57780
rect 200632 57740 200638 57752
rect 201218 57740 201224 57752
rect 201276 57740 201282 57792
rect 201678 57740 201684 57792
rect 201736 57780 201742 57792
rect 202322 57780 202328 57792
rect 201736 57752 202328 57780
rect 201736 57740 201742 57752
rect 202322 57740 202328 57752
rect 202380 57740 202386 57792
rect 203242 57740 203248 57792
rect 203300 57780 203306 57792
rect 204070 57780 204076 57792
rect 203300 57752 204076 57780
rect 203300 57740 203306 57752
rect 204070 57740 204076 57752
rect 204128 57740 204134 57792
rect 210878 57740 210884 57792
rect 210936 57780 210942 57792
rect 220170 57780 220176 57792
rect 210936 57752 220176 57780
rect 210936 57740 210942 57752
rect 220170 57740 220176 57752
rect 220228 57740 220234 57792
rect 221200 57780 221228 57888
rect 221274 57876 221280 57928
rect 221332 57916 221338 57928
rect 225782 57916 225788 57928
rect 221332 57888 225788 57916
rect 221332 57876 221338 57888
rect 225782 57876 225788 57888
rect 225840 57876 225846 57928
rect 221826 57808 221832 57860
rect 221884 57848 221890 57860
rect 222930 57848 222936 57860
rect 221884 57820 222936 57848
rect 221884 57808 221890 57820
rect 222930 57808 222936 57820
rect 222988 57808 222994 57860
rect 223022 57808 223028 57860
rect 223080 57848 223086 57860
rect 228358 57848 228364 57860
rect 223080 57820 228364 57848
rect 223080 57808 223086 57820
rect 228358 57808 228364 57820
rect 228416 57808 228422 57860
rect 224310 57780 224316 57792
rect 221200 57752 224316 57780
rect 224310 57740 224316 57752
rect 224368 57740 224374 57792
rect 213270 57712 213276 57724
rect 179156 57684 213276 57712
rect 213270 57672 213276 57684
rect 213328 57672 213334 57724
rect 213362 57672 213368 57724
rect 213420 57712 213426 57724
rect 215110 57712 215116 57724
rect 213420 57684 215116 57712
rect 213420 57672 213426 57684
rect 215110 57672 215116 57684
rect 215168 57672 215174 57724
rect 215202 57672 215208 57724
rect 215260 57712 215266 57724
rect 223390 57712 223396 57724
rect 215260 57684 223396 57712
rect 215260 57672 215266 57684
rect 223390 57672 223396 57684
rect 223448 57672 223454 57724
rect 96540 57616 97028 57644
rect 97074 57604 97080 57656
rect 97132 57644 97138 57656
rect 97132 57616 98500 57644
rect 97132 57604 97138 57616
rect 97258 57576 97264 57588
rect 95528 57548 97264 57576
rect 97258 57536 97264 57548
rect 97316 57536 97322 57588
rect 98472 57576 98500 57616
rect 98546 57604 98552 57656
rect 98604 57644 98610 57656
rect 99282 57644 99288 57656
rect 98604 57616 99288 57644
rect 98604 57604 98610 57616
rect 99282 57604 99288 57616
rect 99340 57604 99346 57656
rect 100018 57604 100024 57656
rect 100076 57644 100082 57656
rect 100570 57644 100576 57656
rect 100076 57616 100576 57644
rect 100076 57604 100082 57616
rect 100570 57604 100576 57616
rect 100628 57604 100634 57656
rect 101122 57604 101128 57656
rect 101180 57644 101186 57656
rect 101858 57644 101864 57656
rect 101180 57616 101864 57644
rect 101180 57604 101186 57616
rect 101858 57604 101864 57616
rect 101916 57604 101922 57656
rect 103238 57604 103244 57656
rect 103296 57644 103302 57656
rect 172698 57644 172704 57656
rect 103296 57616 172704 57644
rect 103296 57604 103302 57616
rect 172698 57604 172704 57616
rect 172756 57604 172762 57656
rect 172790 57604 172796 57656
rect 172848 57644 172854 57656
rect 173526 57644 173532 57656
rect 172848 57616 173532 57644
rect 172848 57604 172854 57616
rect 173526 57604 173532 57616
rect 173584 57604 173590 57656
rect 174630 57604 174636 57656
rect 174688 57644 174694 57656
rect 175182 57644 175188 57656
rect 174688 57616 175188 57644
rect 174688 57604 174694 57616
rect 175182 57604 175188 57616
rect 175240 57604 175246 57656
rect 177022 57604 177028 57656
rect 177080 57644 177086 57656
rect 177574 57644 177580 57656
rect 177080 57616 177580 57644
rect 177080 57604 177086 57616
rect 177574 57604 177580 57616
rect 177632 57604 177638 57656
rect 177666 57604 177672 57656
rect 177724 57644 177730 57656
rect 177942 57644 177948 57656
rect 177724 57616 177948 57644
rect 177724 57604 177730 57616
rect 177942 57604 177948 57616
rect 178000 57604 178006 57656
rect 178770 57604 178776 57656
rect 178828 57644 178834 57656
rect 179230 57644 179236 57656
rect 178828 57616 179236 57644
rect 178828 57604 178834 57616
rect 179230 57604 179236 57616
rect 179288 57604 179294 57656
rect 179598 57604 179604 57656
rect 179656 57644 179662 57656
rect 180426 57644 180432 57656
rect 179656 57616 180432 57644
rect 179656 57604 179662 57616
rect 180426 57604 180432 57616
rect 180484 57604 180490 57656
rect 182266 57604 182272 57656
rect 182324 57644 182330 57656
rect 183094 57644 183100 57656
rect 182324 57616 183100 57644
rect 182324 57604 182330 57616
rect 183094 57604 183100 57616
rect 183152 57604 183158 57656
rect 183922 57604 183928 57656
rect 183980 57644 183986 57656
rect 184842 57644 184848 57656
rect 183980 57616 184848 57644
rect 183980 57604 183986 57616
rect 184842 57604 184848 57616
rect 184900 57604 184906 57656
rect 185026 57604 185032 57656
rect 185084 57644 185090 57656
rect 185762 57644 185768 57656
rect 185084 57616 185768 57644
rect 185084 57604 185090 57616
rect 185762 57604 185768 57616
rect 185820 57604 185826 57656
rect 188614 57604 188620 57656
rect 188672 57644 188678 57656
rect 188982 57644 188988 57656
rect 188672 57616 188988 57644
rect 188672 57604 188678 57616
rect 188982 57604 188988 57616
rect 189040 57604 189046 57656
rect 189350 57604 189356 57656
rect 189408 57644 189414 57656
rect 190086 57644 190092 57656
rect 189408 57616 190092 57644
rect 189408 57604 189414 57616
rect 190086 57604 190092 57616
rect 190144 57604 190150 57656
rect 190362 57604 190368 57656
rect 190420 57644 190426 57656
rect 216030 57644 216036 57656
rect 190420 57616 216036 57644
rect 190420 57604 190426 57616
rect 216030 57604 216036 57616
rect 216088 57604 216094 57656
rect 217226 57604 217232 57656
rect 217284 57644 217290 57656
rect 223942 57644 223948 57656
rect 217284 57616 223948 57644
rect 217284 57604 217290 57616
rect 223942 57604 223948 57616
rect 224000 57604 224006 57656
rect 103054 57576 103060 57588
rect 98472 57548 103060 57576
rect 103054 57536 103060 57548
rect 103112 57536 103118 57588
rect 104342 57536 104348 57588
rect 104400 57576 104406 57588
rect 104710 57576 104716 57588
rect 104400 57548 104716 57576
rect 104400 57536 104406 57548
rect 104710 57536 104716 57548
rect 104768 57536 104774 57588
rect 106734 57536 106740 57588
rect 106792 57576 106798 57588
rect 107470 57576 107476 57588
rect 106792 57548 107476 57576
rect 106792 57536 106798 57548
rect 107470 57536 107476 57548
rect 107528 57536 107534 57588
rect 108206 57536 108212 57588
rect 108264 57576 108270 57588
rect 113726 57576 113732 57588
rect 108264 57548 113732 57576
rect 108264 57536 108270 57548
rect 113726 57536 113732 57548
rect 113784 57536 113790 57588
rect 113818 57536 113824 57588
rect 113876 57576 113882 57588
rect 142522 57576 142528 57588
rect 113876 57548 142528 57576
rect 113876 57536 113882 57548
rect 142522 57536 142528 57548
rect 142580 57536 142586 57588
rect 142614 57536 142620 57588
rect 142672 57576 142678 57588
rect 143442 57576 143448 57588
rect 142672 57548 143448 57576
rect 142672 57536 142678 57548
rect 143442 57536 143448 57548
rect 143500 57536 143506 57588
rect 143534 57536 143540 57588
rect 143592 57576 143598 57588
rect 143592 57548 146616 57576
rect 143592 57536 143598 57548
rect 92676 57480 93256 57508
rect 70268 57412 76236 57440
rect 70268 57400 70274 57412
rect 77202 57400 77208 57452
rect 77260 57440 77266 57452
rect 78674 57440 78680 57452
rect 77260 57412 78680 57440
rect 77260 57400 77266 57412
rect 78674 57400 78680 57412
rect 78732 57400 78738 57452
rect 81618 57400 81624 57452
rect 81676 57440 81682 57452
rect 82722 57440 82728 57452
rect 81676 57412 82728 57440
rect 81676 57400 81682 57412
rect 82722 57400 82728 57412
rect 82780 57400 82786 57452
rect 83090 57400 83096 57452
rect 83148 57440 83154 57452
rect 93118 57440 93124 57452
rect 83148 57412 93124 57440
rect 83148 57400 83154 57412
rect 93118 57400 93124 57412
rect 93176 57400 93182 57452
rect 93228 57440 93256 57480
rect 93854 57468 93860 57520
rect 93912 57508 93918 57520
rect 95050 57508 95056 57520
rect 93912 57480 95056 57508
rect 93912 57468 93918 57480
rect 95050 57468 95056 57480
rect 95108 57468 95114 57520
rect 95326 57468 95332 57520
rect 95384 57508 95390 57520
rect 96430 57508 96436 57520
rect 95384 57480 96436 57508
rect 95384 57468 95390 57480
rect 96430 57468 96436 57480
rect 96488 57468 96494 57520
rect 96706 57468 96712 57520
rect 96764 57508 96770 57520
rect 100754 57508 100760 57520
rect 96764 57480 100760 57508
rect 96764 57468 96770 57480
rect 100754 57468 100760 57480
rect 100812 57468 100818 57520
rect 100846 57468 100852 57520
rect 100904 57508 100910 57520
rect 101950 57508 101956 57520
rect 100904 57480 101956 57508
rect 100904 57468 100910 57480
rect 101950 57468 101956 57480
rect 102008 57468 102014 57520
rect 102134 57468 102140 57520
rect 102192 57508 102198 57520
rect 133046 57508 133052 57520
rect 102192 57480 133052 57508
rect 102192 57468 102198 57480
rect 133046 57468 133052 57480
rect 133104 57468 133110 57520
rect 133230 57468 133236 57520
rect 133288 57508 133294 57520
rect 133690 57508 133696 57520
rect 133288 57480 133696 57508
rect 133288 57468 133294 57480
rect 133690 57468 133696 57480
rect 133748 57468 133754 57520
rect 134150 57468 134156 57520
rect 134208 57508 134214 57520
rect 134886 57508 134892 57520
rect 134208 57480 134892 57508
rect 134208 57468 134214 57480
rect 134886 57468 134892 57480
rect 134944 57468 134950 57520
rect 135898 57468 135904 57520
rect 135956 57508 135962 57520
rect 136358 57508 136364 57520
rect 135956 57480 136364 57508
rect 135956 57468 135962 57480
rect 136358 57468 136364 57480
rect 136416 57468 136422 57520
rect 136450 57468 136456 57520
rect 136508 57508 136514 57520
rect 137186 57508 137192 57520
rect 136508 57480 137192 57508
rect 136508 57468 136514 57480
rect 137186 57468 137192 57480
rect 137244 57468 137250 57520
rect 138106 57468 138112 57520
rect 138164 57508 138170 57520
rect 139118 57508 139124 57520
rect 138164 57480 139124 57508
rect 138164 57468 138170 57480
rect 139118 57468 139124 57480
rect 139176 57468 139182 57520
rect 139946 57468 139952 57520
rect 140004 57508 140010 57520
rect 140774 57508 140780 57520
rect 140004 57480 140780 57508
rect 140004 57468 140010 57480
rect 140774 57468 140780 57480
rect 140832 57468 140838 57520
rect 141142 57468 141148 57520
rect 141200 57508 141206 57520
rect 141970 57508 141976 57520
rect 141200 57480 141976 57508
rect 141200 57468 141206 57480
rect 141970 57468 141976 57480
rect 142028 57468 142034 57520
rect 142246 57468 142252 57520
rect 142304 57508 142310 57520
rect 144178 57508 144184 57520
rect 142304 57480 144184 57508
rect 142304 57468 142310 57480
rect 144178 57468 144184 57480
rect 144236 57468 144242 57520
rect 144270 57468 144276 57520
rect 144328 57508 144334 57520
rect 144822 57508 144828 57520
rect 144328 57480 144828 57508
rect 144328 57468 144334 57480
rect 144822 57468 144828 57480
rect 144880 57468 144886 57520
rect 145190 57468 145196 57520
rect 145248 57508 145254 57520
rect 146110 57508 146116 57520
rect 145248 57480 146116 57508
rect 145248 57468 145254 57480
rect 146110 57468 146116 57480
rect 146168 57468 146174 57520
rect 146588 57508 146616 57548
rect 146662 57536 146668 57588
rect 146720 57576 146726 57588
rect 147490 57576 147496 57588
rect 146720 57548 147496 57576
rect 146720 57536 146726 57548
rect 147490 57536 147496 57548
rect 147548 57536 147554 57588
rect 147674 57536 147680 57588
rect 147732 57576 147738 57588
rect 152182 57576 152188 57588
rect 147732 57548 152188 57576
rect 147732 57536 147738 57548
rect 152182 57536 152188 57548
rect 152240 57536 152246 57588
rect 152458 57536 152464 57588
rect 152516 57576 152522 57588
rect 222930 57576 222936 57588
rect 152516 57548 222936 57576
rect 152516 57536 152522 57548
rect 222930 57536 222936 57548
rect 222988 57536 222994 57588
rect 223022 57536 223028 57588
rect 223080 57576 223086 57588
rect 225874 57576 225880 57588
rect 223080 57548 225880 57576
rect 223080 57536 223086 57548
rect 225874 57536 225880 57548
rect 225932 57536 225938 57588
rect 147306 57508 147312 57520
rect 146588 57480 147312 57508
rect 147306 57468 147312 57480
rect 147364 57468 147370 57520
rect 148042 57468 148048 57520
rect 148100 57508 148106 57520
rect 148962 57508 148968 57520
rect 148100 57480 148968 57508
rect 148100 57468 148106 57480
rect 148962 57468 148968 57480
rect 149020 57468 149026 57520
rect 150250 57468 150256 57520
rect 150308 57508 150314 57520
rect 214558 57508 214564 57520
rect 150308 57480 214564 57508
rect 150308 57468 150314 57480
rect 214558 57468 214564 57480
rect 214616 57468 214622 57520
rect 215110 57468 215116 57520
rect 215168 57508 215174 57520
rect 216766 57508 216772 57520
rect 215168 57480 216772 57508
rect 215168 57468 215174 57480
rect 216766 57468 216772 57480
rect 216824 57468 216830 57520
rect 219434 57468 219440 57520
rect 219492 57508 219498 57520
rect 226150 57508 226156 57520
rect 219492 57480 226156 57508
rect 219492 57468 219498 57480
rect 226150 57468 226156 57480
rect 226208 57468 226214 57520
rect 101398 57440 101404 57452
rect 93228 57412 101404 57440
rect 101398 57400 101404 57412
rect 101456 57400 101462 57452
rect 101582 57400 101588 57452
rect 101640 57440 101646 57452
rect 113818 57440 113824 57452
rect 101640 57412 113824 57440
rect 101640 57400 101646 57412
rect 113818 57400 113824 57412
rect 113876 57400 113882 57452
rect 113910 57400 113916 57452
rect 113968 57440 113974 57452
rect 118602 57440 118608 57452
rect 113968 57412 118608 57440
rect 113968 57400 113974 57412
rect 118602 57400 118608 57412
rect 118660 57400 118666 57452
rect 118786 57400 118792 57452
rect 118844 57440 118850 57452
rect 128262 57440 128268 57452
rect 118844 57412 128268 57440
rect 118844 57400 118850 57412
rect 128262 57400 128268 57412
rect 128320 57400 128326 57452
rect 128538 57400 128544 57452
rect 128596 57440 128602 57452
rect 129642 57440 129648 57452
rect 128596 57412 129648 57440
rect 128596 57400 128602 57412
rect 129642 57400 129648 57412
rect 129700 57400 129706 57452
rect 130746 57400 130752 57452
rect 130804 57440 130810 57452
rect 130930 57440 130936 57452
rect 130804 57412 130936 57440
rect 130804 57400 130810 57412
rect 130930 57400 130936 57412
rect 130988 57400 130994 57452
rect 131114 57400 131120 57452
rect 131172 57440 131178 57452
rect 132034 57440 132040 57452
rect 131172 57412 132040 57440
rect 131172 57400 131178 57412
rect 132034 57400 132040 57412
rect 132092 57400 132098 57452
rect 132770 57400 132776 57452
rect 132828 57440 132834 57452
rect 133782 57440 133788 57452
rect 132828 57412 133788 57440
rect 132828 57400 132834 57412
rect 133782 57400 133788 57412
rect 133840 57400 133846 57452
rect 134426 57400 134432 57452
rect 134484 57440 134490 57452
rect 134978 57440 134984 57452
rect 134484 57412 134984 57440
rect 134484 57400 134490 57412
rect 134978 57400 134984 57412
rect 135036 57400 135042 57452
rect 135622 57400 135628 57452
rect 135680 57440 135686 57452
rect 136542 57440 136548 57452
rect 135680 57412 136548 57440
rect 135680 57400 135686 57412
rect 136542 57400 136548 57412
rect 136600 57400 136606 57452
rect 136726 57400 136732 57452
rect 136784 57440 136790 57452
rect 137830 57440 137836 57452
rect 136784 57412 137836 57440
rect 136784 57400 136790 57412
rect 137830 57400 137836 57412
rect 137888 57400 137894 57452
rect 139394 57400 139400 57452
rect 139452 57440 139458 57452
rect 140590 57440 140596 57452
rect 139452 57412 140596 57440
rect 139452 57400 139458 57412
rect 140590 57400 140596 57412
rect 140648 57400 140654 57452
rect 140958 57400 140964 57452
rect 141016 57440 141022 57452
rect 222378 57440 222384 57452
rect 141016 57412 222384 57440
rect 141016 57400 141022 57412
rect 222378 57400 222384 57412
rect 222436 57400 222442 57452
rect 27522 57332 27528 57384
rect 27580 57372 27586 57384
rect 66438 57372 66444 57384
rect 27580 57344 66444 57372
rect 27580 57332 27586 57344
rect 66438 57332 66444 57344
rect 66496 57332 66502 57384
rect 67542 57332 67548 57384
rect 67600 57372 67606 57384
rect 76374 57372 76380 57384
rect 67600 57344 76380 57372
rect 67600 57332 67606 57344
rect 76374 57332 76380 57344
rect 76432 57332 76438 57384
rect 87138 57332 87144 57384
rect 87196 57372 87202 57384
rect 93946 57372 93952 57384
rect 87196 57344 93952 57372
rect 87196 57332 87202 57344
rect 93946 57332 93952 57344
rect 94004 57332 94010 57384
rect 94590 57332 94596 57384
rect 94648 57372 94654 57384
rect 103606 57372 103612 57384
rect 94648 57344 103612 57372
rect 94648 57332 94654 57344
rect 103606 57332 103612 57344
rect 103664 57332 103670 57384
rect 103790 57332 103796 57384
rect 103848 57372 103854 57384
rect 104526 57372 104532 57384
rect 103848 57344 104532 57372
rect 103848 57332 103854 57344
rect 104526 57332 104532 57344
rect 104584 57332 104590 57384
rect 105814 57332 105820 57384
rect 105872 57372 105878 57384
rect 117314 57372 117320 57384
rect 105872 57344 117320 57372
rect 105872 57332 105878 57344
rect 117314 57332 117320 57344
rect 117372 57332 117378 57384
rect 118970 57332 118976 57384
rect 119028 57372 119034 57384
rect 201770 57372 201776 57384
rect 119028 57344 201776 57372
rect 119028 57332 119034 57344
rect 201770 57332 201776 57344
rect 201828 57332 201834 57384
rect 202046 57332 202052 57384
rect 202104 57372 202110 57384
rect 202782 57372 202788 57384
rect 202104 57344 202788 57372
rect 202104 57332 202110 57344
rect 202782 57332 202788 57344
rect 202840 57332 202846 57384
rect 203978 57332 203984 57384
rect 204036 57372 204042 57384
rect 208486 57372 208492 57384
rect 204036 57344 208492 57372
rect 204036 57332 204042 57344
rect 208486 57332 208492 57344
rect 208544 57332 208550 57384
rect 210234 57332 210240 57384
rect 210292 57372 210298 57384
rect 214374 57372 214380 57384
rect 210292 57344 214380 57372
rect 210292 57332 210298 57344
rect 214374 57332 214380 57344
rect 214432 57332 214438 57384
rect 214466 57332 214472 57384
rect 214524 57372 214530 57384
rect 225322 57372 225328 57384
rect 214524 57344 225328 57372
rect 214524 57332 214530 57344
rect 225322 57332 225328 57344
rect 225380 57332 225386 57384
rect 6822 57264 6828 57316
rect 6880 57304 6886 57316
rect 59262 57304 59268 57316
rect 6880 57276 59268 57304
rect 6880 57264 6886 57276
rect 59262 57264 59268 57276
rect 59320 57264 59326 57316
rect 59446 57264 59452 57316
rect 59504 57304 59510 57316
rect 60458 57304 60464 57316
rect 59504 57276 60464 57304
rect 59504 57264 59510 57276
rect 60458 57264 60464 57276
rect 60516 57264 60522 57316
rect 62022 57264 62028 57316
rect 62080 57304 62086 57316
rect 75178 57304 75184 57316
rect 62080 57276 75184 57304
rect 62080 57264 62086 57276
rect 75178 57264 75184 57276
rect 75236 57264 75242 57316
rect 82170 57264 82176 57316
rect 82228 57304 82234 57316
rect 90174 57304 90180 57316
rect 82228 57276 90180 57304
rect 82228 57264 82234 57276
rect 90174 57264 90180 57276
rect 90232 57264 90238 57316
rect 91830 57264 91836 57316
rect 91888 57304 91894 57316
rect 118510 57304 118516 57316
rect 91888 57276 118516 57304
rect 91888 57264 91894 57276
rect 118510 57264 118516 57276
rect 118568 57264 118574 57316
rect 120442 57264 120448 57316
rect 120500 57304 120506 57316
rect 121178 57304 121184 57316
rect 120500 57276 121184 57304
rect 120500 57264 120506 57276
rect 121178 57264 121184 57276
rect 121236 57264 121242 57316
rect 122834 57264 122840 57316
rect 122892 57304 122898 57316
rect 123294 57304 123300 57316
rect 122892 57276 123300 57304
rect 122892 57264 122898 57276
rect 123294 57264 123300 57276
rect 123352 57264 123358 57316
rect 124398 57264 124404 57316
rect 124456 57304 124462 57316
rect 125042 57304 125048 57316
rect 124456 57276 125048 57304
rect 124456 57264 124462 57276
rect 125042 57264 125048 57276
rect 125100 57264 125106 57316
rect 125686 57264 125692 57316
rect 125744 57304 125750 57316
rect 126606 57304 126612 57316
rect 125744 57276 126612 57304
rect 125744 57264 125750 57276
rect 126606 57264 126612 57276
rect 126664 57264 126670 57316
rect 127066 57264 127072 57316
rect 127124 57304 127130 57316
rect 127986 57304 127992 57316
rect 127124 57276 127992 57304
rect 127124 57264 127130 57276
rect 127986 57264 127992 57276
rect 128044 57264 128050 57316
rect 128170 57264 128176 57316
rect 128228 57304 128234 57316
rect 129826 57304 129832 57316
rect 128228 57276 129832 57304
rect 128228 57264 128234 57276
rect 129826 57264 129832 57276
rect 129884 57264 129890 57316
rect 130010 57264 130016 57316
rect 130068 57304 130074 57316
rect 131022 57304 131028 57316
rect 130068 57276 131028 57304
rect 130068 57264 130074 57276
rect 131022 57264 131028 57276
rect 131080 57264 131086 57316
rect 131482 57264 131488 57316
rect 131540 57304 131546 57316
rect 132126 57304 132132 57316
rect 131540 57276 132132 57304
rect 131540 57264 131546 57276
rect 132126 57264 132132 57276
rect 132184 57264 132190 57316
rect 132494 57264 132500 57316
rect 132552 57304 132558 57316
rect 223022 57304 223028 57316
rect 132552 57276 223028 57304
rect 132552 57264 132558 57276
rect 223022 57264 223028 57276
rect 223080 57264 223086 57316
rect 24762 57196 24768 57248
rect 24820 57236 24826 57248
rect 65886 57236 65892 57248
rect 24820 57208 65892 57236
rect 24820 57196 24826 57208
rect 65886 57196 65892 57208
rect 65944 57196 65950 57248
rect 68922 57196 68928 57248
rect 68980 57236 68986 57248
rect 76466 57236 76472 57248
rect 68980 57208 76472 57236
rect 68980 57196 68986 57208
rect 76466 57196 76472 57208
rect 76524 57196 76530 57248
rect 83734 57196 83740 57248
rect 83792 57236 83798 57248
rect 96706 57236 96712 57248
rect 83792 57208 96712 57236
rect 83792 57196 83798 57208
rect 96706 57196 96712 57208
rect 96764 57196 96770 57248
rect 104158 57236 104164 57248
rect 98656 57208 104164 57236
rect 43438 57128 43444 57180
rect 43496 57168 43502 57180
rect 61838 57168 61844 57180
rect 43496 57140 61844 57168
rect 43496 57128 43502 57140
rect 61838 57128 61844 57140
rect 61896 57128 61902 57180
rect 61930 57128 61936 57180
rect 61988 57168 61994 57180
rect 64874 57168 64880 57180
rect 61988 57140 64880 57168
rect 61988 57128 61994 57140
rect 64874 57128 64880 57140
rect 64932 57128 64938 57180
rect 65242 57128 65248 57180
rect 65300 57168 65306 57180
rect 65300 57140 65840 57168
rect 65300 57128 65306 57140
rect 46842 57060 46848 57112
rect 46900 57100 46906 57112
rect 65812 57100 65840 57140
rect 68646 57128 68652 57180
rect 68704 57168 68710 57180
rect 74074 57168 74080 57180
rect 68704 57140 74080 57168
rect 68704 57128 68710 57140
rect 74074 57128 74080 57140
rect 74132 57128 74138 57180
rect 89806 57128 89812 57180
rect 89864 57168 89870 57180
rect 98656 57168 98684 57208
rect 104158 57196 104164 57208
rect 104216 57196 104222 57248
rect 104986 57196 104992 57248
rect 105044 57236 105050 57248
rect 108206 57236 108212 57248
rect 105044 57208 108212 57236
rect 105044 57196 105050 57208
rect 108206 57196 108212 57208
rect 108264 57196 108270 57248
rect 108298 57196 108304 57248
rect 108356 57236 108362 57248
rect 147674 57236 147680 57248
rect 108356 57208 147680 57236
rect 108356 57196 108362 57208
rect 147674 57196 147680 57208
rect 147732 57196 147738 57248
rect 147950 57196 147956 57248
rect 148008 57236 148014 57248
rect 151814 57236 151820 57248
rect 148008 57208 151820 57236
rect 148008 57196 148014 57208
rect 151814 57196 151820 57208
rect 151872 57196 151878 57248
rect 155402 57196 155408 57248
rect 155460 57236 155466 57248
rect 166442 57236 166448 57248
rect 155460 57208 166448 57236
rect 155460 57196 155466 57208
rect 166442 57196 166448 57208
rect 166500 57196 166506 57248
rect 166810 57196 166816 57248
rect 166868 57236 166874 57248
rect 401594 57236 401600 57248
rect 166868 57208 401600 57236
rect 166868 57196 166874 57208
rect 401594 57196 401600 57208
rect 401652 57196 401658 57248
rect 89864 57140 98684 57168
rect 89864 57128 89870 57140
rect 103514 57128 103520 57180
rect 103572 57168 103578 57180
rect 143258 57168 143264 57180
rect 103572 57140 143264 57168
rect 103572 57128 103578 57140
rect 143258 57128 143264 57140
rect 143316 57128 143322 57180
rect 143534 57128 143540 57180
rect 143592 57168 143598 57180
rect 144638 57168 144644 57180
rect 143592 57140 144644 57168
rect 143592 57128 143598 57140
rect 144638 57128 144644 57140
rect 144696 57128 144702 57180
rect 144822 57128 144828 57180
rect 144880 57168 144886 57180
rect 146294 57168 146300 57180
rect 144880 57140 146300 57168
rect 144880 57128 144886 57140
rect 146294 57128 146300 57140
rect 146352 57128 146358 57180
rect 146386 57128 146392 57180
rect 146444 57168 146450 57180
rect 152458 57168 152464 57180
rect 146444 57140 152464 57168
rect 146444 57128 146450 57140
rect 152458 57128 152464 57140
rect 152516 57128 152522 57180
rect 156138 57168 156144 57180
rect 152568 57140 156144 57168
rect 74350 57100 74356 57112
rect 46900 57072 65656 57100
rect 65812 57072 74356 57100
rect 46900 57060 46906 57072
rect 49602 56992 49608 57044
rect 49660 57032 49666 57044
rect 63770 57032 63776 57044
rect 49660 57004 63776 57032
rect 49660 56992 49666 57004
rect 63770 56992 63776 57004
rect 63828 56992 63834 57044
rect 65628 57032 65656 57072
rect 74350 57060 74356 57072
rect 74408 57060 74414 57112
rect 96154 57060 96160 57112
rect 96212 57100 96218 57112
rect 96522 57100 96528 57112
rect 96212 57072 96528 57100
rect 96212 57060 96218 57072
rect 96522 57060 96528 57072
rect 96580 57060 96586 57112
rect 98270 57060 98276 57112
rect 98328 57100 98334 57112
rect 99006 57100 99012 57112
rect 98328 57072 99012 57100
rect 98328 57060 98334 57072
rect 99006 57060 99012 57072
rect 99064 57060 99070 57112
rect 99098 57060 99104 57112
rect 99156 57100 99162 57112
rect 99156 57072 103008 57100
rect 99156 57060 99162 57072
rect 71406 57032 71412 57044
rect 65260 57004 65564 57032
rect 65628 57004 71412 57032
rect 48222 56924 48228 56976
rect 48280 56964 48286 56976
rect 65260 56964 65288 57004
rect 48280 56936 65288 56964
rect 65536 56964 65564 57004
rect 71406 56992 71412 57004
rect 71464 56992 71470 57044
rect 79870 56992 79876 57044
rect 79928 57032 79934 57044
rect 80422 57032 80428 57044
rect 79928 57004 80428 57032
rect 79928 56992 79934 57004
rect 80422 56992 80428 57004
rect 80480 56992 80486 57044
rect 88886 56992 88892 57044
rect 88944 57032 88950 57044
rect 102870 57032 102876 57044
rect 88944 57004 102876 57032
rect 88944 56992 88950 57004
rect 102870 56992 102876 57004
rect 102928 56992 102934 57044
rect 71498 56964 71504 56976
rect 65536 56936 71504 56964
rect 48280 56924 48286 56936
rect 71498 56924 71504 56936
rect 71556 56924 71562 56976
rect 74810 56924 74816 56976
rect 74868 56964 74874 56976
rect 74994 56964 75000 56976
rect 74868 56936 75000 56964
rect 74868 56924 74874 56936
rect 74994 56924 75000 56936
rect 75052 56924 75058 56976
rect 93946 56924 93952 56976
rect 94004 56964 94010 56976
rect 102778 56964 102784 56976
rect 94004 56936 102784 56964
rect 94004 56924 94010 56936
rect 102778 56924 102784 56936
rect 102836 56924 102842 56976
rect 102980 56964 103008 57072
rect 103698 57060 103704 57112
rect 103756 57100 103762 57112
rect 104802 57100 104808 57112
rect 103756 57072 104808 57100
rect 103756 57060 103762 57072
rect 104802 57060 104808 57072
rect 104860 57060 104866 57112
rect 105170 57060 105176 57112
rect 105228 57100 105234 57112
rect 152568 57100 152596 57140
rect 156138 57128 156144 57140
rect 156196 57128 156202 57180
rect 210878 57168 210884 57180
rect 157306 57140 210884 57168
rect 105228 57072 152596 57100
rect 105228 57060 105234 57072
rect 153654 57060 153660 57112
rect 153712 57100 153718 57112
rect 154482 57100 154488 57112
rect 153712 57072 154488 57100
rect 153712 57060 153718 57072
rect 154482 57060 154488 57072
rect 154540 57060 154546 57112
rect 156322 57060 156328 57112
rect 156380 57100 156386 57112
rect 157306 57100 157334 57140
rect 210878 57128 210884 57140
rect 210936 57128 210942 57180
rect 212258 57128 212264 57180
rect 212316 57168 212322 57180
rect 212316 57140 213684 57168
rect 212316 57128 212322 57140
rect 156380 57072 157334 57100
rect 156380 57060 156386 57072
rect 162026 57060 162032 57112
rect 162084 57100 162090 57112
rect 168558 57100 168564 57112
rect 162084 57072 168564 57100
rect 162084 57060 162090 57072
rect 168558 57060 168564 57072
rect 168616 57060 168622 57112
rect 168650 57060 168656 57112
rect 168708 57100 168714 57112
rect 213362 57100 213368 57112
rect 168708 57072 213368 57100
rect 168708 57060 168714 57072
rect 213362 57060 213368 57072
rect 213420 57060 213426 57112
rect 213656 57100 213684 57140
rect 213730 57128 213736 57180
rect 213788 57168 213794 57180
rect 213788 57140 216720 57168
rect 213788 57128 213794 57140
rect 215386 57100 215392 57112
rect 213656 57072 215392 57100
rect 215386 57060 215392 57072
rect 215444 57060 215450 57112
rect 215478 57060 215484 57112
rect 215536 57100 215542 57112
rect 216582 57100 216588 57112
rect 215536 57072 216588 57100
rect 215536 57060 215542 57072
rect 216582 57060 216588 57072
rect 216640 57060 216646 57112
rect 216692 57100 216720 57140
rect 216766 57128 216772 57180
rect 216824 57168 216830 57180
rect 216824 57140 222148 57168
rect 216824 57128 216830 57140
rect 222010 57100 222016 57112
rect 216692 57072 222016 57100
rect 222010 57060 222016 57072
rect 222068 57060 222074 57112
rect 222120 57100 222148 57140
rect 222194 57128 222200 57180
rect 222252 57168 222258 57180
rect 300118 57168 300124 57180
rect 222252 57140 300124 57168
rect 222252 57128 222258 57140
rect 300118 57128 300124 57140
rect 300176 57128 300182 57180
rect 224126 57100 224132 57112
rect 222120 57072 224132 57100
rect 224126 57060 224132 57072
rect 224184 57060 224190 57112
rect 103054 56992 103060 57044
rect 103112 57032 103118 57044
rect 132678 57032 132684 57044
rect 103112 57004 132684 57032
rect 103112 56992 103118 57004
rect 132678 56992 132684 57004
rect 132736 56992 132742 57044
rect 132862 56992 132868 57044
rect 132920 57032 132926 57044
rect 142154 57032 142160 57044
rect 132920 57004 142160 57032
rect 132920 56992 132926 57004
rect 142154 56992 142160 57004
rect 142212 56992 142218 57044
rect 142246 56992 142252 57044
rect 142304 57032 142310 57044
rect 142304 57004 161152 57032
rect 142304 56992 142310 57004
rect 133782 56964 133788 56976
rect 102980 56936 133788 56964
rect 133782 56924 133788 56936
rect 133840 56924 133846 56976
rect 135438 56964 135444 56976
rect 133892 56936 135444 56964
rect 53742 56856 53748 56908
rect 53800 56896 53806 56908
rect 65150 56896 65156 56908
rect 53800 56868 65156 56896
rect 53800 56856 53806 56868
rect 65150 56856 65156 56868
rect 65208 56856 65214 56908
rect 65518 56856 65524 56908
rect 65576 56896 65582 56908
rect 71774 56896 71780 56908
rect 65576 56868 71780 56896
rect 65576 56856 65582 56868
rect 71774 56856 71780 56868
rect 71832 56856 71838 56908
rect 76558 56856 76564 56908
rect 76616 56896 76622 56908
rect 78122 56896 78128 56908
rect 76616 56868 78128 56896
rect 76616 56856 76622 56868
rect 78122 56856 78128 56868
rect 78180 56856 78186 56908
rect 93302 56856 93308 56908
rect 93360 56896 93366 56908
rect 133892 56896 133920 56936
rect 135438 56924 135444 56936
rect 135496 56924 135502 56976
rect 137002 56924 137008 56976
rect 137060 56964 137066 56976
rect 141326 56964 141332 56976
rect 137060 56936 141332 56964
rect 137060 56924 137066 56936
rect 141326 56924 141332 56936
rect 141384 56924 141390 56976
rect 141418 56924 141424 56976
rect 141476 56964 141482 56976
rect 146938 56964 146944 56976
rect 141476 56936 146944 56964
rect 141476 56924 141482 56936
rect 146938 56924 146944 56936
rect 146996 56924 147002 56976
rect 147306 56924 147312 56976
rect 147364 56964 147370 56976
rect 150250 56964 150256 56976
rect 147364 56936 150256 56964
rect 147364 56924 147370 56936
rect 150250 56924 150256 56936
rect 150308 56924 150314 56976
rect 150434 56924 150440 56976
rect 150492 56964 150498 56976
rect 151538 56964 151544 56976
rect 150492 56936 151544 56964
rect 150492 56924 150498 56936
rect 151538 56924 151544 56936
rect 151596 56924 151602 56976
rect 151906 56924 151912 56976
rect 151964 56964 151970 56976
rect 153102 56964 153108 56976
rect 151964 56936 153108 56964
rect 151964 56924 151970 56936
rect 153102 56924 153108 56936
rect 153160 56924 153166 56976
rect 153378 56924 153384 56976
rect 153436 56964 153442 56976
rect 154206 56964 154212 56976
rect 153436 56936 154212 56964
rect 153436 56924 153442 56936
rect 154206 56924 154212 56936
rect 154264 56924 154270 56976
rect 154574 56924 154580 56976
rect 154632 56964 154638 56976
rect 155862 56964 155868 56976
rect 154632 56936 155868 56964
rect 154632 56924 154638 56936
rect 155862 56924 155868 56936
rect 155920 56924 155926 56976
rect 155954 56924 155960 56976
rect 156012 56964 156018 56976
rect 157058 56964 157064 56976
rect 156012 56936 157064 56964
rect 156012 56924 156018 56936
rect 157058 56924 157064 56936
rect 157116 56924 157122 56976
rect 161124 56964 161152 57004
rect 161566 56992 161572 57044
rect 161624 57032 161630 57044
rect 166350 57032 166356 57044
rect 161624 57004 166356 57032
rect 161624 56992 161630 57004
rect 166350 56992 166356 57004
rect 166408 56992 166414 57044
rect 166902 56992 166908 57044
rect 166960 57032 166966 57044
rect 166960 57004 213684 57032
rect 166960 56992 166966 57004
rect 162762 56964 162768 56976
rect 161124 56936 162768 56964
rect 162762 56924 162768 56936
rect 162820 56924 162826 56976
rect 163314 56924 163320 56976
rect 163372 56964 163378 56976
rect 166810 56964 166816 56976
rect 163372 56936 166816 56964
rect 163372 56924 163378 56936
rect 166810 56924 166816 56936
rect 166868 56924 166874 56976
rect 167178 56924 167184 56976
rect 167236 56964 167242 56976
rect 213546 56964 213552 56976
rect 167236 56936 213552 56964
rect 167236 56924 167242 56936
rect 213546 56924 213552 56936
rect 213604 56924 213610 56976
rect 213656 56964 213684 57004
rect 214558 56992 214564 57044
rect 214616 57032 214622 57044
rect 220262 57032 220268 57044
rect 214616 57004 220268 57032
rect 214616 56992 214622 57004
rect 220262 56992 220268 57004
rect 220320 56992 220326 57044
rect 220722 56992 220728 57044
rect 220780 57032 220786 57044
rect 302234 57032 302240 57044
rect 220780 57004 302240 57032
rect 220780 56992 220786 57004
rect 302234 56992 302240 57004
rect 302292 56992 302298 57044
rect 215938 56964 215944 56976
rect 213656 56936 215944 56964
rect 215938 56924 215944 56936
rect 215996 56924 216002 56976
rect 216582 56924 216588 56976
rect 216640 56964 216646 56976
rect 277486 56964 277492 56976
rect 216640 56936 277492 56964
rect 216640 56924 216646 56936
rect 277486 56924 277492 56936
rect 277544 56924 277550 56976
rect 93360 56868 133920 56896
rect 93360 56856 93366 56868
rect 133966 56856 133972 56908
rect 134024 56896 134030 56908
rect 134702 56896 134708 56908
rect 134024 56868 134708 56896
rect 134024 56856 134030 56868
rect 134702 56856 134708 56868
rect 134760 56856 134766 56908
rect 134794 56856 134800 56908
rect 134852 56896 134858 56908
rect 138658 56896 138664 56908
rect 134852 56868 138664 56896
rect 134852 56856 134858 56868
rect 138658 56856 138664 56868
rect 138716 56856 138722 56908
rect 138750 56856 138756 56908
rect 138808 56896 138814 56908
rect 142062 56896 142068 56908
rect 138808 56868 142068 56896
rect 138808 56856 138814 56868
rect 142062 56856 142068 56868
rect 142120 56856 142126 56908
rect 142172 56868 142384 56896
rect 53650 56788 53656 56840
rect 53708 56828 53714 56840
rect 63402 56828 63408 56840
rect 53708 56800 63408 56828
rect 53708 56788 53714 56800
rect 63402 56788 63408 56800
rect 63460 56788 63466 56840
rect 65610 56788 65616 56840
rect 65668 56828 65674 56840
rect 72878 56828 72884 56840
rect 65668 56800 72884 56828
rect 65668 56788 65674 56800
rect 72878 56788 72884 56800
rect 72936 56788 72942 56840
rect 89162 56788 89168 56840
rect 89220 56828 89226 56840
rect 89530 56828 89536 56840
rect 89220 56800 89536 56828
rect 89220 56788 89226 56800
rect 89530 56788 89536 56800
rect 89588 56788 89594 56840
rect 90726 56788 90732 56840
rect 90784 56828 90790 56840
rect 91002 56828 91008 56840
rect 90784 56800 91008 56828
rect 90784 56788 90790 56800
rect 91002 56788 91008 56800
rect 91060 56788 91066 56840
rect 91554 56788 91560 56840
rect 91612 56828 91618 56840
rect 94590 56828 94596 56840
rect 91612 56800 94596 56828
rect 91612 56788 91618 56800
rect 94590 56788 94596 56800
rect 94648 56788 94654 56840
rect 94682 56788 94688 56840
rect 94740 56828 94746 56840
rect 99098 56828 99104 56840
rect 94740 56800 99104 56828
rect 94740 56788 94746 56800
rect 99098 56788 99104 56800
rect 99156 56788 99162 56840
rect 99742 56788 99748 56840
rect 99800 56828 99806 56840
rect 105170 56828 105176 56840
rect 99800 56800 105176 56828
rect 99800 56788 99806 56800
rect 105170 56788 105176 56800
rect 105228 56788 105234 56840
rect 105262 56788 105268 56840
rect 105320 56828 105326 56840
rect 106182 56828 106188 56840
rect 105320 56800 106188 56828
rect 105320 56788 105326 56800
rect 106182 56788 106188 56800
rect 106240 56788 106246 56840
rect 107838 56788 107844 56840
rect 107896 56828 107902 56840
rect 108758 56828 108764 56840
rect 107896 56800 108764 56828
rect 107896 56788 107902 56800
rect 108758 56788 108764 56800
rect 108816 56788 108822 56840
rect 110230 56788 110236 56840
rect 110288 56828 110294 56840
rect 113634 56828 113640 56840
rect 110288 56800 113640 56828
rect 110288 56788 110294 56800
rect 113634 56788 113640 56800
rect 113692 56788 113698 56840
rect 113726 56788 113732 56840
rect 113784 56828 113790 56840
rect 132494 56828 132500 56840
rect 113784 56800 132500 56828
rect 113784 56788 113790 56800
rect 132494 56788 132500 56800
rect 132552 56788 132558 56840
rect 132678 56788 132684 56840
rect 132736 56828 132742 56840
rect 142172 56828 142200 56868
rect 132736 56800 142200 56828
rect 142356 56828 142384 56868
rect 142522 56856 142528 56908
rect 142580 56896 142586 56908
rect 144914 56896 144920 56908
rect 142580 56868 144920 56896
rect 142580 56856 142586 56868
rect 144914 56856 144920 56868
rect 144972 56856 144978 56908
rect 145098 56856 145104 56908
rect 145156 56896 145162 56908
rect 180886 56896 180892 56908
rect 145156 56868 157104 56896
rect 145156 56856 145162 56868
rect 146570 56828 146576 56840
rect 142356 56800 146576 56828
rect 132736 56788 132742 56800
rect 146570 56788 146576 56800
rect 146628 56788 146634 56840
rect 146662 56788 146668 56840
rect 146720 56828 146726 56840
rect 156046 56828 156052 56840
rect 146720 56800 156052 56828
rect 146720 56788 146726 56800
rect 156046 56788 156052 56800
rect 156104 56788 156110 56840
rect 157076 56828 157104 56868
rect 157260 56868 180892 56896
rect 157260 56828 157288 56868
rect 180886 56856 180892 56868
rect 180944 56856 180950 56908
rect 180978 56856 180984 56908
rect 181036 56896 181042 56908
rect 181898 56896 181904 56908
rect 181036 56868 181904 56896
rect 181036 56856 181042 56868
rect 181898 56856 181904 56868
rect 181956 56856 181962 56908
rect 182542 56856 182548 56908
rect 182600 56896 182606 56908
rect 183278 56896 183284 56908
rect 182600 56868 183284 56896
rect 182600 56856 182606 56868
rect 183278 56856 183284 56868
rect 183336 56856 183342 56908
rect 186314 56856 186320 56908
rect 186372 56896 186378 56908
rect 187234 56896 187240 56908
rect 186372 56868 187240 56896
rect 186372 56856 186378 56868
rect 187234 56856 187240 56868
rect 187292 56856 187298 56908
rect 190730 56856 190736 56908
rect 190788 56896 190794 56908
rect 191650 56896 191656 56908
rect 190788 56868 191656 56896
rect 190788 56856 190794 56868
rect 191650 56856 191656 56868
rect 191708 56856 191714 56908
rect 191834 56856 191840 56908
rect 191892 56896 191898 56908
rect 193030 56896 193036 56908
rect 191892 56868 193036 56896
rect 191892 56856 191898 56868
rect 193030 56856 193036 56868
rect 193088 56856 193094 56908
rect 193582 56856 193588 56908
rect 193640 56896 193646 56908
rect 194226 56896 194232 56908
rect 193640 56868 194232 56896
rect 193640 56856 193646 56868
rect 194226 56856 194232 56868
rect 194284 56856 194290 56908
rect 194594 56856 194600 56908
rect 194652 56896 194658 56908
rect 195698 56896 195704 56908
rect 194652 56868 195704 56896
rect 194652 56856 194658 56868
rect 195698 56856 195704 56868
rect 195756 56856 195762 56908
rect 198274 56856 198280 56908
rect 198332 56896 198338 56908
rect 198550 56896 198556 56908
rect 198332 56868 198556 56896
rect 198332 56856 198338 56868
rect 198550 56856 198556 56868
rect 198608 56856 198614 56908
rect 198734 56856 198740 56908
rect 198792 56896 198798 56908
rect 200022 56896 200028 56908
rect 198792 56868 200028 56896
rect 198792 56856 198798 56868
rect 200022 56856 200028 56868
rect 200080 56856 200086 56908
rect 201770 56856 201776 56908
rect 201828 56896 201834 56908
rect 203518 56896 203524 56908
rect 201828 56868 203524 56896
rect 201828 56856 201834 56868
rect 203518 56856 203524 56868
rect 203576 56856 203582 56908
rect 204714 56856 204720 56908
rect 204772 56896 204778 56908
rect 204772 56868 204944 56896
rect 204772 56856 204778 56868
rect 157076 56800 157288 56828
rect 157444 56800 172468 56828
rect 55122 56720 55128 56772
rect 55180 56760 55186 56772
rect 64782 56760 64788 56772
rect 55180 56732 64788 56760
rect 55180 56720 55186 56732
rect 64782 56720 64788 56732
rect 64840 56720 64846 56772
rect 65334 56720 65340 56772
rect 65392 56760 65398 56772
rect 73154 56760 73160 56772
rect 65392 56732 73160 56760
rect 65392 56720 65398 56732
rect 73154 56720 73160 56732
rect 73212 56720 73218 56772
rect 84838 56720 84844 56772
rect 84896 56760 84902 56772
rect 86218 56760 86224 56772
rect 84896 56732 86224 56760
rect 84896 56720 84902 56732
rect 86218 56720 86224 56732
rect 86276 56720 86282 56772
rect 98822 56720 98828 56772
rect 98880 56760 98886 56772
rect 99190 56760 99196 56772
rect 98880 56732 99196 56760
rect 98880 56720 98886 56732
rect 99190 56720 99196 56732
rect 99248 56720 99254 56772
rect 99374 56720 99380 56772
rect 99432 56760 99438 56772
rect 100662 56760 100668 56772
rect 99432 56732 100668 56760
rect 99432 56720 99438 56732
rect 100662 56720 100668 56732
rect 100720 56720 100726 56772
rect 100754 56720 100760 56772
rect 100812 56760 100818 56772
rect 103054 56760 103060 56772
rect 100812 56732 103060 56760
rect 100812 56720 100818 56732
rect 103054 56720 103060 56732
rect 103112 56720 103118 56772
rect 103606 56720 103612 56772
rect 103664 56760 103670 56772
rect 105538 56760 105544 56772
rect 103664 56732 105544 56760
rect 103664 56720 103670 56732
rect 105538 56720 105544 56732
rect 105596 56720 105602 56772
rect 106366 56720 106372 56772
rect 106424 56760 106430 56772
rect 107562 56760 107568 56772
rect 106424 56732 107568 56760
rect 106424 56720 106430 56732
rect 107562 56720 107568 56732
rect 107620 56720 107626 56772
rect 107654 56720 107660 56772
rect 107712 56760 107718 56772
rect 108482 56760 108488 56772
rect 107712 56732 108488 56760
rect 107712 56720 107718 56732
rect 108482 56720 108488 56732
rect 108540 56720 108546 56772
rect 113910 56760 113916 56772
rect 108776 56732 108988 56760
rect 59262 56652 59268 56704
rect 59320 56692 59326 56704
rect 69658 56692 69664 56704
rect 59320 56664 65196 56692
rect 59320 56652 59326 56664
rect 57238 56584 57244 56636
rect 57296 56624 57302 56636
rect 64690 56624 64696 56636
rect 57296 56596 64696 56624
rect 57296 56584 57302 56596
rect 64690 56584 64696 56596
rect 64748 56584 64754 56636
rect 65168 56624 65196 56664
rect 65720 56664 69664 56692
rect 65242 56624 65248 56636
rect 65168 56596 65248 56624
rect 65242 56584 65248 56596
rect 65300 56584 65306 56636
rect 64874 56516 64880 56568
rect 64932 56556 64938 56568
rect 65720 56556 65748 56664
rect 69658 56652 69664 56664
rect 69716 56652 69722 56704
rect 70302 56652 70308 56704
rect 70360 56692 70366 56704
rect 76926 56692 76932 56704
rect 70360 56664 76932 56692
rect 70360 56652 70366 56664
rect 76926 56652 76932 56664
rect 76984 56652 76990 56704
rect 90082 56652 90088 56704
rect 90140 56692 90146 56704
rect 91002 56692 91008 56704
rect 90140 56664 91008 56692
rect 90140 56652 90146 56664
rect 91002 56652 91008 56664
rect 91060 56652 91066 56704
rect 97994 56652 98000 56704
rect 98052 56692 98058 56704
rect 99098 56692 99104 56704
rect 98052 56664 99104 56692
rect 98052 56652 98058 56664
rect 99098 56652 99104 56664
rect 99156 56652 99162 56704
rect 102594 56652 102600 56704
rect 102652 56692 102658 56704
rect 103330 56692 103336 56704
rect 102652 56664 103336 56692
rect 102652 56652 102658 56664
rect 103330 56652 103336 56664
rect 103388 56652 103394 56704
rect 104066 56652 104072 56704
rect 104124 56692 104130 56704
rect 108776 56692 108804 56732
rect 104124 56664 108804 56692
rect 104124 56652 104130 56664
rect 73430 56624 73436 56636
rect 64932 56528 65748 56556
rect 65812 56596 73436 56624
rect 64932 56516 64938 56528
rect 64782 56448 64788 56500
rect 64840 56488 64846 56500
rect 65812 56488 65840 56596
rect 73430 56584 73436 56596
rect 73488 56584 73494 56636
rect 97626 56584 97632 56636
rect 97684 56624 97690 56636
rect 108298 56624 108304 56636
rect 97684 56596 108304 56624
rect 97684 56584 97690 56596
rect 108298 56584 108304 56596
rect 108356 56584 108362 56636
rect 108960 56624 108988 56732
rect 109236 56732 113916 56760
rect 109236 56624 109264 56732
rect 113910 56720 113916 56732
rect 113968 56720 113974 56772
rect 114094 56720 114100 56772
rect 114152 56760 114158 56772
rect 118602 56760 118608 56772
rect 114152 56732 118608 56760
rect 114152 56720 114158 56732
rect 118602 56720 118608 56732
rect 118660 56720 118666 56772
rect 118694 56720 118700 56772
rect 118752 56760 118758 56772
rect 119798 56760 119804 56772
rect 118752 56732 119804 56760
rect 118752 56720 118758 56732
rect 119798 56720 119804 56732
rect 119856 56720 119862 56772
rect 120074 56720 120080 56772
rect 120132 56760 120138 56772
rect 120718 56760 120724 56772
rect 120132 56732 120724 56760
rect 120132 56720 120138 56732
rect 120718 56720 120724 56732
rect 120776 56720 120782 56772
rect 123294 56720 123300 56772
rect 123352 56760 123358 56772
rect 123938 56760 123944 56772
rect 123352 56732 123944 56760
rect 123352 56720 123358 56732
rect 123938 56720 123944 56732
rect 123996 56720 124002 56772
rect 124582 56720 124588 56772
rect 124640 56760 124646 56772
rect 125410 56760 125416 56772
rect 124640 56732 125416 56760
rect 124640 56720 124646 56732
rect 125410 56720 125416 56732
rect 125468 56720 125474 56772
rect 125594 56720 125600 56772
rect 125652 56760 125658 56772
rect 126238 56760 126244 56772
rect 125652 56732 126244 56760
rect 125652 56720 125658 56732
rect 126238 56720 126244 56732
rect 126296 56720 126302 56772
rect 126330 56720 126336 56772
rect 126388 56760 126394 56772
rect 129734 56760 129740 56772
rect 126388 56732 129740 56760
rect 126388 56720 126394 56732
rect 129734 56720 129740 56732
rect 129792 56720 129798 56772
rect 129826 56720 129832 56772
rect 129884 56760 129890 56772
rect 130378 56760 130384 56772
rect 129884 56732 130384 56760
rect 129884 56720 129890 56732
rect 130378 56720 130384 56732
rect 130436 56720 130442 56772
rect 131206 56720 131212 56772
rect 131264 56760 131270 56772
rect 132402 56760 132408 56772
rect 131264 56732 132408 56760
rect 131264 56720 131270 56732
rect 132402 56720 132408 56732
rect 132460 56720 132466 56772
rect 133782 56720 133788 56772
rect 133840 56760 133846 56772
rect 136726 56760 136732 56772
rect 133840 56732 136732 56760
rect 133840 56720 133846 56732
rect 136726 56720 136732 56732
rect 136784 56720 136790 56772
rect 136818 56720 136824 56772
rect 136876 56760 136882 56772
rect 138014 56760 138020 56772
rect 136876 56732 138020 56760
rect 136876 56720 136882 56732
rect 138014 56720 138020 56732
rect 138072 56720 138078 56772
rect 138474 56720 138480 56772
rect 138532 56760 138538 56772
rect 139118 56760 139124 56772
rect 138532 56732 139124 56760
rect 138532 56720 138538 56732
rect 139118 56720 139124 56732
rect 139176 56720 139182 56772
rect 139210 56720 139216 56772
rect 139268 56760 139274 56772
rect 142062 56760 142068 56772
rect 139268 56732 142068 56760
rect 139268 56720 139274 56732
rect 142062 56720 142068 56732
rect 142120 56720 142126 56772
rect 146846 56760 146852 56772
rect 142172 56732 146852 56760
rect 110782 56652 110788 56704
rect 110840 56692 110846 56704
rect 110840 56664 113404 56692
rect 110840 56652 110846 56664
rect 108960 56596 109264 56624
rect 109310 56584 109316 56636
rect 109368 56624 109374 56636
rect 110322 56624 110328 56636
rect 109368 56596 110328 56624
rect 109368 56584 109374 56596
rect 110322 56584 110328 56596
rect 110380 56584 110386 56636
rect 110506 56584 110512 56636
rect 110564 56624 110570 56636
rect 111610 56624 111616 56636
rect 110564 56596 111616 56624
rect 110564 56584 110570 56596
rect 111610 56584 111616 56596
rect 111668 56584 111674 56636
rect 112254 56584 112260 56636
rect 112312 56624 112318 56636
rect 112990 56624 112996 56636
rect 112312 56596 112996 56624
rect 112312 56584 112318 56596
rect 112990 56584 112996 56596
rect 113048 56584 113054 56636
rect 113376 56624 113404 56664
rect 113450 56652 113456 56704
rect 113508 56692 113514 56704
rect 114370 56692 114376 56704
rect 113508 56664 114376 56692
rect 113508 56652 113514 56664
rect 114370 56652 114376 56664
rect 114428 56652 114434 56704
rect 115198 56652 115204 56704
rect 115256 56692 115262 56704
rect 115750 56692 115756 56704
rect 115256 56664 115756 56692
rect 115256 56652 115262 56664
rect 115750 56652 115756 56664
rect 115808 56652 115814 56704
rect 116026 56652 116032 56704
rect 116084 56692 116090 56704
rect 117130 56692 117136 56704
rect 116084 56664 117136 56692
rect 116084 56652 116090 56664
rect 117130 56652 117136 56664
rect 117188 56652 117194 56704
rect 142172 56692 142200 56732
rect 146846 56720 146852 56732
rect 146904 56720 146910 56772
rect 146938 56720 146944 56772
rect 146996 56760 147002 56772
rect 157444 56760 157472 56800
rect 146996 56732 157472 56760
rect 146996 56720 147002 56732
rect 162946 56720 162952 56772
rect 163004 56760 163010 56772
rect 164050 56760 164056 56772
rect 163004 56732 164056 56760
rect 163004 56720 163010 56732
rect 164050 56720 164056 56732
rect 164108 56720 164114 56772
rect 165614 56720 165620 56772
rect 165672 56760 165678 56772
rect 166718 56760 166724 56772
rect 165672 56732 166724 56760
rect 165672 56720 165678 56732
rect 166718 56720 166724 56732
rect 166776 56720 166782 56772
rect 166810 56720 166816 56772
rect 166868 56760 166874 56772
rect 167178 56760 167184 56772
rect 166868 56732 167184 56760
rect 166868 56720 166874 56732
rect 167178 56720 167184 56732
rect 167236 56720 167242 56772
rect 168374 56720 168380 56772
rect 168432 56760 168438 56772
rect 169110 56760 169116 56772
rect 168432 56732 169116 56760
rect 168432 56720 168438 56732
rect 169110 56720 169116 56732
rect 169168 56720 169174 56772
rect 170306 56720 170312 56772
rect 170364 56760 170370 56772
rect 171042 56760 171048 56772
rect 170364 56732 171048 56760
rect 170364 56720 170370 56732
rect 171042 56720 171048 56732
rect 171100 56720 171106 56772
rect 171410 56720 171416 56772
rect 171468 56760 171474 56772
rect 172330 56760 172336 56772
rect 171468 56732 172336 56760
rect 171468 56720 171474 56732
rect 172330 56720 172336 56732
rect 172388 56720 172394 56772
rect 172440 56760 172468 56800
rect 172698 56788 172704 56840
rect 172756 56828 172762 56840
rect 174906 56828 174912 56840
rect 172756 56800 174912 56828
rect 172756 56788 172762 56800
rect 174906 56788 174912 56800
rect 174964 56788 174970 56840
rect 175274 56788 175280 56840
rect 175332 56828 175338 56840
rect 176378 56828 176384 56840
rect 175332 56800 176384 56828
rect 175332 56788 175338 56800
rect 176378 56788 176384 56800
rect 176436 56788 176442 56840
rect 204806 56828 204812 56840
rect 176672 56800 204812 56828
rect 175734 56760 175740 56772
rect 172440 56732 175740 56760
rect 175734 56720 175740 56732
rect 175792 56720 175798 56772
rect 175826 56720 175832 56772
rect 175884 56760 175890 56772
rect 176562 56760 176568 56772
rect 175884 56732 176568 56760
rect 175884 56720 175890 56732
rect 176562 56720 176568 56732
rect 176620 56720 176626 56772
rect 117516 56664 142200 56692
rect 113376 56596 113956 56624
rect 113928 56556 113956 56596
rect 114186 56584 114192 56636
rect 114244 56624 114250 56636
rect 114462 56624 114468 56636
rect 114244 56596 114468 56624
rect 114244 56584 114250 56596
rect 114462 56584 114468 56596
rect 114520 56584 114526 56636
rect 114830 56584 114836 56636
rect 114888 56624 114894 56636
rect 115566 56624 115572 56636
rect 114888 56596 115572 56624
rect 114888 56584 114894 56596
rect 115566 56584 115572 56596
rect 115624 56584 115630 56636
rect 116854 56624 116860 56636
rect 115676 56596 116860 56624
rect 115676 56556 115704 56596
rect 116854 56584 116860 56596
rect 116912 56584 116918 56636
rect 116946 56584 116952 56636
rect 117004 56624 117010 56636
rect 117222 56624 117228 56636
rect 117004 56596 117228 56624
rect 117004 56584 117010 56596
rect 117222 56584 117228 56596
rect 117280 56584 117286 56636
rect 113928 56528 115704 56556
rect 64840 56460 65840 56488
rect 64840 56448 64846 56460
rect 113634 56448 113640 56500
rect 113692 56488 113698 56500
rect 117516 56488 117544 56664
rect 142246 56652 142252 56704
rect 142304 56692 142310 56704
rect 147766 56692 147772 56704
rect 142304 56664 147772 56692
rect 142304 56652 142310 56664
rect 147766 56652 147772 56664
rect 147824 56652 147830 56704
rect 147858 56652 147864 56704
rect 147916 56692 147922 56704
rect 148778 56692 148784 56704
rect 147916 56664 148784 56692
rect 147916 56652 147922 56664
rect 148778 56652 148784 56664
rect 148836 56652 148842 56704
rect 149606 56652 149612 56704
rect 149664 56692 149670 56704
rect 150250 56692 150256 56704
rect 149664 56664 150256 56692
rect 149664 56652 149670 56664
rect 150250 56652 150256 56664
rect 150308 56652 150314 56704
rect 151078 56652 151084 56704
rect 151136 56692 151142 56704
rect 151630 56692 151636 56704
rect 151136 56664 151636 56692
rect 151136 56652 151142 56664
rect 151630 56652 151636 56664
rect 151688 56652 151694 56704
rect 152826 56652 152832 56704
rect 152884 56692 152890 56704
rect 153010 56692 153016 56704
rect 152884 56664 153016 56692
rect 152884 56652 152890 56664
rect 153010 56652 153016 56664
rect 153068 56652 153074 56704
rect 153930 56652 153936 56704
rect 153988 56692 153994 56704
rect 154390 56692 154396 56704
rect 153988 56664 154396 56692
rect 153988 56652 153994 56664
rect 154390 56652 154396 56664
rect 154448 56652 154454 56704
rect 154850 56652 154856 56704
rect 154908 56692 154914 56704
rect 155770 56692 155776 56704
rect 154908 56664 155776 56692
rect 154908 56652 154914 56664
rect 155770 56652 155776 56664
rect 155828 56652 155834 56704
rect 156782 56652 156788 56704
rect 156840 56692 156846 56704
rect 170398 56692 170404 56704
rect 156840 56664 170404 56692
rect 156840 56652 156846 56664
rect 170398 56652 170404 56664
rect 170456 56652 170462 56704
rect 173710 56652 173716 56704
rect 173768 56692 173774 56704
rect 176672 56692 176700 56800
rect 204806 56788 204812 56800
rect 204864 56788 204870 56840
rect 204916 56828 204944 56868
rect 205266 56856 205272 56908
rect 205324 56896 205330 56908
rect 213822 56896 213828 56908
rect 205324 56868 213828 56896
rect 205324 56856 205330 56868
rect 213822 56856 213828 56868
rect 213880 56856 213886 56908
rect 214742 56856 214748 56908
rect 214800 56896 214806 56908
rect 229462 56896 229468 56908
rect 214800 56868 229468 56896
rect 214800 56856 214806 56868
rect 229462 56856 229468 56868
rect 229520 56856 229526 56908
rect 209866 56828 209872 56840
rect 204916 56800 209872 56828
rect 209866 56788 209872 56800
rect 209924 56788 209930 56840
rect 213454 56788 213460 56840
rect 213512 56828 213518 56840
rect 213512 56800 216444 56828
rect 213512 56788 213518 56800
rect 176746 56720 176752 56772
rect 176804 56760 176810 56772
rect 180702 56760 180708 56772
rect 176804 56732 180708 56760
rect 176804 56720 176810 56732
rect 180702 56720 180708 56732
rect 180760 56720 180766 56772
rect 180886 56720 180892 56772
rect 180944 56760 180950 56772
rect 182910 56760 182916 56772
rect 180944 56732 182916 56760
rect 180944 56720 180950 56732
rect 182910 56720 182916 56732
rect 182968 56720 182974 56772
rect 183002 56720 183008 56772
rect 183060 56760 183066 56772
rect 190362 56760 190368 56772
rect 183060 56732 190368 56760
rect 183060 56720 183066 56732
rect 190362 56720 190368 56732
rect 190420 56720 190426 56772
rect 193306 56720 193312 56772
rect 193364 56760 193370 56772
rect 194410 56760 194416 56772
rect 193364 56732 194416 56760
rect 193364 56720 193370 56732
rect 194410 56720 194416 56732
rect 194468 56720 194474 56772
rect 197722 56720 197728 56772
rect 197780 56760 197786 56772
rect 198550 56760 198556 56772
rect 197780 56732 198556 56760
rect 197780 56720 197786 56732
rect 198550 56720 198556 56732
rect 198608 56720 198614 56772
rect 200482 56720 200488 56772
rect 200540 56760 200546 56772
rect 200540 56732 205036 56760
rect 200540 56720 200546 56732
rect 173768 56664 176700 56692
rect 173768 56652 173774 56664
rect 179874 56652 179880 56704
rect 179932 56692 179938 56704
rect 180518 56692 180524 56704
rect 179932 56664 180524 56692
rect 179932 56652 179938 56664
rect 180518 56652 180524 56664
rect 180576 56652 180582 56704
rect 180794 56652 180800 56704
rect 180852 56692 180858 56704
rect 204714 56692 204720 56704
rect 180852 56664 204720 56692
rect 180852 56652 180858 56664
rect 204714 56652 204720 56664
rect 204772 56652 204778 56704
rect 205008 56692 205036 56732
rect 206462 56720 206468 56772
rect 206520 56760 206526 56772
rect 214466 56760 214472 56772
rect 206520 56732 214472 56760
rect 206520 56720 206526 56732
rect 214466 56720 214472 56732
rect 214524 56720 214530 56772
rect 214650 56720 214656 56772
rect 214708 56760 214714 56772
rect 216306 56760 216312 56772
rect 214708 56732 216312 56760
rect 214708 56720 214714 56732
rect 216306 56720 216312 56732
rect 216364 56720 216370 56772
rect 216416 56760 216444 56800
rect 216490 56788 216496 56840
rect 216548 56828 216554 56840
rect 221918 56828 221924 56840
rect 216548 56800 221924 56828
rect 216548 56788 216554 56800
rect 221918 56788 221924 56800
rect 221976 56788 221982 56840
rect 222010 56788 222016 56840
rect 222068 56828 222074 56840
rect 226242 56828 226248 56840
rect 222068 56800 226248 56828
rect 222068 56788 222074 56800
rect 226242 56788 226248 56800
rect 226300 56788 226306 56840
rect 225690 56760 225696 56772
rect 216416 56732 225696 56760
rect 225690 56720 225696 56732
rect 225748 56720 225754 56772
rect 208394 56692 208400 56704
rect 205008 56664 208400 56692
rect 208394 56652 208400 56664
rect 208452 56652 208458 56704
rect 208486 56652 208492 56704
rect 208544 56692 208550 56704
rect 214742 56692 214748 56704
rect 208544 56664 214748 56692
rect 208544 56652 208550 56664
rect 214742 56652 214748 56664
rect 214800 56652 214806 56704
rect 215386 56652 215392 56704
rect 215444 56692 215450 56704
rect 221826 56692 221832 56704
rect 215444 56664 221832 56692
rect 215444 56652 215450 56664
rect 221826 56652 221832 56664
rect 221884 56652 221890 56704
rect 221918 56652 221924 56704
rect 221976 56692 221982 56704
rect 225966 56692 225972 56704
rect 221976 56664 225972 56692
rect 221976 56652 221982 56664
rect 225966 56652 225972 56664
rect 226024 56652 226030 56704
rect 142154 56624 142160 56636
rect 113692 56460 117544 56488
rect 117608 56596 142160 56624
rect 113692 56448 113698 56460
rect 117314 56380 117320 56432
rect 117372 56420 117378 56432
rect 117608 56420 117636 56596
rect 142154 56584 142160 56596
rect 142212 56584 142218 56636
rect 156690 56624 156696 56636
rect 142264 56596 156696 56624
rect 118510 56516 118516 56568
rect 118568 56556 118574 56568
rect 120718 56556 120724 56568
rect 118568 56528 120724 56556
rect 118568 56516 118574 56528
rect 120718 56516 120724 56528
rect 120776 56516 120782 56568
rect 128262 56516 128268 56568
rect 128320 56556 128326 56568
rect 129826 56556 129832 56568
rect 128320 56528 129832 56556
rect 128320 56516 128326 56528
rect 129826 56516 129832 56528
rect 129884 56516 129890 56568
rect 139854 56448 139860 56500
rect 139912 56488 139918 56500
rect 142264 56488 142292 56596
rect 156690 56584 156696 56596
rect 156748 56584 156754 56636
rect 158070 56584 158076 56636
rect 158128 56624 158134 56636
rect 158622 56624 158628 56636
rect 158128 56596 158628 56624
rect 158128 56584 158134 56596
rect 158622 56584 158628 56596
rect 158680 56584 158686 56636
rect 158898 56584 158904 56636
rect 158956 56624 158962 56636
rect 160002 56624 160008 56636
rect 158956 56596 160008 56624
rect 158956 56584 158962 56596
rect 160002 56584 160008 56596
rect 160060 56584 160066 56636
rect 160922 56584 160928 56636
rect 160980 56624 160986 56636
rect 161382 56624 161388 56636
rect 160980 56596 161388 56624
rect 160980 56584 160986 56596
rect 161382 56584 161388 56596
rect 161440 56584 161446 56636
rect 162118 56584 162124 56636
rect 162176 56624 162182 56636
rect 162670 56624 162676 56636
rect 162176 56596 162676 56624
rect 162176 56584 162182 56596
rect 162670 56584 162676 56596
rect 162728 56584 162734 56636
rect 162762 56584 162768 56636
rect 162820 56624 162826 56636
rect 162820 56596 163820 56624
rect 162820 56584 162826 56596
rect 163792 56556 163820 56596
rect 163866 56584 163872 56636
rect 163924 56624 163930 56636
rect 164142 56624 164148 56636
rect 163924 56596 164148 56624
rect 163924 56584 163930 56596
rect 164142 56584 164148 56596
rect 164200 56584 164206 56636
rect 164602 56624 164608 56636
rect 164252 56596 164608 56624
rect 164252 56556 164280 56596
rect 164602 56584 164608 56596
rect 164660 56584 164666 56636
rect 164694 56584 164700 56636
rect 164752 56624 164758 56636
rect 165430 56624 165436 56636
rect 164752 56596 165436 56624
rect 164752 56584 164758 56596
rect 165430 56584 165436 56596
rect 165488 56584 165494 56636
rect 166534 56584 166540 56636
rect 166592 56624 166598 56636
rect 166810 56624 166816 56636
rect 166592 56596 166816 56624
rect 166592 56584 166598 56596
rect 166810 56584 166816 56596
rect 166868 56584 166874 56636
rect 219618 56624 219624 56636
rect 166920 56596 219624 56624
rect 163792 56528 164280 56556
rect 166442 56516 166448 56568
rect 166500 56556 166506 56568
rect 166920 56556 166948 56596
rect 219618 56584 219624 56596
rect 219676 56584 219682 56636
rect 219894 56584 219900 56636
rect 219952 56624 219958 56636
rect 276658 56624 276664 56636
rect 219952 56596 276664 56624
rect 219952 56584 219958 56596
rect 276658 56584 276664 56596
rect 276716 56584 276722 56636
rect 166500 56528 166948 56556
rect 166500 56516 166506 56528
rect 174906 56516 174912 56568
rect 174964 56556 174970 56568
rect 175274 56556 175280 56568
rect 174964 56528 175280 56556
rect 174964 56516 174970 56528
rect 175274 56516 175280 56528
rect 175332 56516 175338 56568
rect 182910 56516 182916 56568
rect 182968 56556 182974 56568
rect 184198 56556 184204 56568
rect 182968 56528 184204 56556
rect 182968 56516 182974 56528
rect 184198 56516 184204 56528
rect 184256 56516 184262 56568
rect 184382 56516 184388 56568
rect 184440 56556 184446 56568
rect 450538 56556 450544 56568
rect 184440 56528 450544 56556
rect 184440 56516 184446 56528
rect 450538 56516 450544 56528
rect 450596 56516 450602 56568
rect 139912 56460 142292 56488
rect 139912 56448 139918 56460
rect 180242 56448 180248 56500
rect 180300 56488 180306 56500
rect 447778 56488 447784 56500
rect 180300 56460 447784 56488
rect 180300 56448 180306 56460
rect 447778 56448 447784 56460
rect 447836 56448 447842 56500
rect 117372 56392 117636 56420
rect 117372 56380 117378 56392
rect 142062 56380 142068 56432
rect 142120 56420 142126 56432
rect 142614 56420 142620 56432
rect 142120 56392 142620 56420
rect 142120 56380 142126 56392
rect 142614 56380 142620 56392
rect 142672 56380 142678 56432
rect 175734 56380 175740 56432
rect 175792 56420 175798 56432
rect 178126 56420 178132 56432
rect 175792 56392 178132 56420
rect 175792 56380 175798 56392
rect 178126 56380 178132 56392
rect 178184 56380 178190 56432
rect 182082 56380 182088 56432
rect 182140 56420 182146 56432
rect 454678 56420 454684 56432
rect 182140 56392 454684 56420
rect 182140 56380 182146 56392
rect 454678 56380 454684 56392
rect 454736 56380 454742 56432
rect 182818 56312 182824 56364
rect 182876 56352 182882 56364
rect 461578 56352 461584 56364
rect 182876 56324 461584 56352
rect 182876 56312 182882 56324
rect 461578 56312 461584 56324
rect 461636 56312 461642 56364
rect 178402 56244 178408 56296
rect 178460 56284 178466 56296
rect 479518 56284 479524 56296
rect 178460 56256 479524 56284
rect 178460 56244 178466 56256
rect 479518 56244 479524 56256
rect 479576 56244 479582 56296
rect 74810 56176 74816 56228
rect 74868 56216 74874 56228
rect 75638 56216 75644 56228
rect 74868 56188 75644 56216
rect 74868 56176 74874 56188
rect 75638 56176 75644 56188
rect 75696 56176 75702 56228
rect 181070 56176 181076 56228
rect 181128 56216 181134 56228
rect 184382 56216 184388 56228
rect 181128 56188 184388 56216
rect 181128 56176 181134 56188
rect 184382 56176 184388 56188
rect 184440 56176 184446 56228
rect 184566 56176 184572 56228
rect 184624 56216 184630 56228
rect 468478 56216 468484 56228
rect 184624 56188 468484 56216
rect 184624 56176 184630 56188
rect 468478 56176 468484 56188
rect 468536 56176 468542 56228
rect 179322 56108 179328 56160
rect 179380 56148 179386 56160
rect 483014 56148 483020 56160
rect 179380 56120 483020 56148
rect 179380 56108 179386 56120
rect 483014 56108 483020 56120
rect 483072 56108 483078 56160
rect 183738 56040 183744 56092
rect 183796 56080 183802 56092
rect 500954 56080 500960 56092
rect 183796 56052 500960 56080
rect 183796 56040 183802 56052
rect 500954 56040 500960 56052
rect 501012 56040 501018 56092
rect 185486 55972 185492 56024
rect 185544 56012 185550 56024
rect 507854 56012 507860 56024
rect 185544 55984 507860 56012
rect 185544 55972 185550 55984
rect 507854 55972 507860 55984
rect 507912 55972 507918 56024
rect 129734 55904 129740 55956
rect 129792 55944 129798 55956
rect 178034 55944 178040 55956
rect 129792 55916 178040 55944
rect 129792 55904 129798 55916
rect 178034 55904 178040 55916
rect 178092 55904 178098 55956
rect 189258 55904 189264 55956
rect 189316 55944 189322 55956
rect 519538 55944 519544 55956
rect 189316 55916 519544 55944
rect 189316 55904 189322 55916
rect 519538 55904 519544 55916
rect 519596 55904 519602 55956
rect 55766 55836 55772 55888
rect 55824 55876 55830 55888
rect 580350 55876 580356 55888
rect 55824 55848 580356 55876
rect 55824 55836 55830 55848
rect 580350 55836 580356 55848
rect 580408 55836 580414 55888
rect 112806 55768 112812 55820
rect 112864 55768 112870 55820
rect 167362 55768 167368 55820
rect 167420 55808 167426 55820
rect 434714 55808 434720 55820
rect 167420 55780 434720 55808
rect 167420 55768 167426 55780
rect 434714 55768 434720 55780
rect 434772 55768 434778 55820
rect 63494 55564 63500 55616
rect 63552 55604 63558 55616
rect 64230 55604 64236 55616
rect 63552 55576 64236 55604
rect 63552 55564 63558 55576
rect 64230 55564 64236 55576
rect 64288 55564 64294 55616
rect 63678 55496 63684 55548
rect 63736 55536 63742 55548
rect 64506 55536 64512 55548
rect 63736 55508 64512 55536
rect 63736 55496 63742 55508
rect 64506 55496 64512 55508
rect 64564 55496 64570 55548
rect 112824 55536 112852 55768
rect 127894 55700 127900 55752
rect 127952 55740 127958 55752
rect 128170 55740 128176 55752
rect 127952 55712 128176 55740
rect 127952 55700 127958 55712
rect 128170 55700 128176 55712
rect 128228 55700 128234 55752
rect 152366 55700 152372 55752
rect 152424 55740 152430 55752
rect 152826 55740 152832 55752
rect 152424 55712 152832 55740
rect 152424 55700 152430 55712
rect 152826 55700 152832 55712
rect 152884 55700 152890 55752
rect 163590 55700 163596 55752
rect 163648 55740 163654 55752
rect 417418 55740 417424 55752
rect 163648 55712 417424 55740
rect 163648 55700 163654 55712
rect 417418 55700 417424 55712
rect 417476 55700 417482 55752
rect 116302 55632 116308 55684
rect 116360 55672 116366 55684
rect 227714 55672 227720 55684
rect 116360 55644 227720 55672
rect 116360 55632 116366 55644
rect 227714 55632 227720 55644
rect 227772 55632 227778 55684
rect 114554 55564 114560 55616
rect 114612 55604 114618 55616
rect 220814 55604 220820 55616
rect 114612 55576 220820 55604
rect 114612 55564 114618 55576
rect 220814 55564 220820 55576
rect 220872 55564 220878 55616
rect 213914 55536 213920 55548
rect 112824 55508 213920 55536
rect 213914 55496 213920 55508
rect 213972 55496 213978 55548
rect 111058 55428 111064 55480
rect 111116 55468 111122 55480
rect 207014 55468 207020 55480
rect 111116 55440 207020 55468
rect 111116 55428 111122 55440
rect 207014 55428 207020 55440
rect 207072 55428 207078 55480
rect 111978 55360 111984 55412
rect 112036 55400 112042 55412
rect 209774 55400 209780 55412
rect 112036 55372 209780 55400
rect 112036 55360 112042 55372
rect 209774 55360 209780 55372
rect 209832 55360 209838 55412
rect 112714 55292 112720 55344
rect 112772 55332 112778 55344
rect 112898 55332 112904 55344
rect 112772 55304 112904 55332
rect 112772 55292 112778 55304
rect 112898 55292 112904 55304
rect 112956 55292 112962 55344
rect 158254 55292 158260 55344
rect 158312 55332 158318 55344
rect 158530 55332 158536 55344
rect 158312 55304 158536 55332
rect 158312 55292 158318 55304
rect 158530 55292 158536 55304
rect 158588 55292 158594 55344
rect 137094 55156 137100 55208
rect 137152 55196 137158 55208
rect 313274 55196 313280 55208
rect 137152 55168 313280 55196
rect 137152 55156 137158 55168
rect 313274 55156 313280 55168
rect 313332 55156 313338 55208
rect 138290 55088 138296 55140
rect 138348 55128 138354 55140
rect 316034 55128 316040 55140
rect 138348 55100 316040 55128
rect 138348 55088 138354 55100
rect 316034 55088 316040 55100
rect 316092 55088 316098 55140
rect 138106 55020 138112 55072
rect 138164 55060 138170 55072
rect 320174 55060 320180 55072
rect 138164 55032 320180 55060
rect 138164 55020 138170 55032
rect 320174 55020 320180 55032
rect 320232 55020 320238 55072
rect 140774 54952 140780 55004
rect 140832 54992 140838 55004
rect 324314 54992 324320 55004
rect 140832 54964 324320 54992
rect 140832 54952 140838 54964
rect 324314 54952 324320 54964
rect 324372 54952 324378 55004
rect 140866 54884 140872 54936
rect 140924 54924 140930 54936
rect 327074 54924 327080 54936
rect 140924 54896 327080 54924
rect 140924 54884 140930 54896
rect 327074 54884 327080 54896
rect 327132 54884 327138 54936
rect 157610 54816 157616 54868
rect 157668 54856 157674 54868
rect 158530 54856 158536 54868
rect 157668 54828 158536 54856
rect 157668 54816 157674 54828
rect 158530 54816 158536 54828
rect 158588 54816 158594 54868
rect 160094 54816 160100 54868
rect 160152 54856 160158 54868
rect 405734 54856 405740 54868
rect 160152 54828 405740 54856
rect 160152 54816 160158 54828
rect 405734 54816 405740 54828
rect 405792 54816 405798 54868
rect 161842 54748 161848 54800
rect 161900 54788 161906 54800
rect 412634 54788 412640 54800
rect 161900 54760 412640 54788
rect 161900 54748 161906 54760
rect 412634 54748 412640 54760
rect 412692 54748 412698 54800
rect 166166 54680 166172 54732
rect 166224 54720 166230 54732
rect 430574 54720 430580 54732
rect 166224 54692 430580 54720
rect 166224 54680 166230 54692
rect 430574 54680 430580 54692
rect 430632 54680 430638 54732
rect 60642 54612 60648 54664
rect 60700 54652 60706 54664
rect 74994 54652 75000 54664
rect 60700 54624 75000 54652
rect 60700 54612 60706 54624
rect 74994 54612 75000 54624
rect 75052 54612 75058 54664
rect 166994 54612 167000 54664
rect 167052 54652 167058 54664
rect 438854 54652 438860 54664
rect 167052 54624 438860 54652
rect 167052 54612 167058 54624
rect 438854 54612 438860 54624
rect 438912 54612 438918 54664
rect 50982 54544 50988 54596
rect 51040 54584 51046 54596
rect 71866 54584 71872 54596
rect 51040 54556 71872 54584
rect 51040 54544 51046 54556
rect 71866 54544 71872 54556
rect 71924 54544 71930 54596
rect 185026 54544 185032 54596
rect 185084 54584 185090 54596
rect 475378 54584 475384 54596
rect 185084 54556 475384 54584
rect 185084 54544 185090 54556
rect 475378 54544 475384 54556
rect 475436 54544 475442 54596
rect 38562 54476 38568 54528
rect 38620 54516 38626 54528
rect 69382 54516 69388 54528
rect 38620 54488 69388 54516
rect 38620 54476 38626 54488
rect 69382 54476 69388 54488
rect 69440 54476 69446 54528
rect 189350 54476 189356 54528
rect 189408 54516 189414 54528
rect 526438 54516 526444 54528
rect 189408 54488 526444 54516
rect 189408 54476 189414 54488
rect 526438 54476 526444 54488
rect 526496 54476 526502 54528
rect 137186 54408 137192 54460
rect 137244 54448 137250 54460
rect 309134 54448 309140 54460
rect 137244 54420 309140 54448
rect 137244 54408 137250 54420
rect 309134 54408 309140 54420
rect 309192 54408 309198 54460
rect 133966 54340 133972 54392
rect 134024 54380 134030 54392
rect 302234 54380 302240 54392
rect 134024 54352 302240 54380
rect 134024 54340 134030 54352
rect 302234 54340 302240 54352
rect 302292 54340 302298 54392
rect 131114 54272 131120 54324
rect 131172 54312 131178 54324
rect 132310 54312 132316 54324
rect 131172 54284 132316 54312
rect 131172 54272 131178 54284
rect 132310 54272 132316 54284
rect 132368 54272 132374 54324
rect 132770 54272 132776 54324
rect 132828 54312 132834 54324
rect 299474 54312 299480 54324
rect 132828 54284 299480 54312
rect 132828 54272 132834 54284
rect 299474 54272 299480 54284
rect 299532 54272 299538 54324
rect 129734 54204 129740 54256
rect 129792 54244 129798 54256
rect 218054 54244 218060 54256
rect 129792 54216 218060 54244
rect 129792 54204 129798 54216
rect 218054 54204 218060 54216
rect 218112 54204 218118 54256
rect 161382 53728 161388 53780
rect 161440 53768 161446 53780
rect 407758 53768 407764 53780
rect 161440 53740 407764 53768
rect 161440 53728 161446 53740
rect 407758 53728 407764 53740
rect 407816 53728 407822 53780
rect 162578 53660 162584 53712
rect 162636 53700 162642 53712
rect 414658 53700 414664 53712
rect 162636 53672 414664 53700
rect 162636 53660 162642 53672
rect 414658 53660 414664 53672
rect 414716 53660 414722 53712
rect 164418 53592 164424 53644
rect 164476 53632 164482 53644
rect 421558 53632 421564 53644
rect 164476 53604 421564 53632
rect 164476 53592 164482 53604
rect 421558 53592 421564 53604
rect 421616 53592 421622 53644
rect 186774 53524 186780 53576
rect 186832 53564 186838 53576
rect 443638 53564 443644 53576
rect 186832 53536 443644 53564
rect 186832 53524 186838 53536
rect 443638 53524 443644 53536
rect 443696 53524 443702 53576
rect 165338 53456 165344 53508
rect 165396 53496 165402 53508
rect 425698 53496 425704 53508
rect 165396 53468 425704 53496
rect 165396 53456 165402 53468
rect 425698 53456 425704 53468
rect 425756 53456 425762 53508
rect 171502 53388 171508 53440
rect 171560 53428 171566 53440
rect 452654 53428 452660 53440
rect 171560 53400 452660 53428
rect 171560 53388 171566 53400
rect 452654 53388 452660 53400
rect 452712 53388 452718 53440
rect 183922 53320 183928 53372
rect 183980 53360 183986 53372
rect 472618 53360 472624 53372
rect 183980 53332 472624 53360
rect 183980 53320 183986 53332
rect 472618 53320 472624 53332
rect 472676 53320 472682 53372
rect 183830 53252 183836 53304
rect 183888 53292 183894 53304
rect 502334 53292 502340 53304
rect 183888 53264 502340 53292
rect 183888 53252 183894 53264
rect 502334 53252 502340 53264
rect 502392 53252 502398 53304
rect 186590 53184 186596 53236
rect 186648 53224 186654 53236
rect 512638 53224 512644 53236
rect 186648 53196 512644 53224
rect 186648 53184 186654 53196
rect 512638 53184 512644 53196
rect 512696 53184 512702 53236
rect 188154 53116 188160 53168
rect 188212 53156 188218 53168
rect 520274 53156 520280 53168
rect 188212 53128 520280 53156
rect 188212 53116 188218 53128
rect 520274 53116 520280 53128
rect 520332 53116 520338 53168
rect 190822 53048 190828 53100
rect 190880 53088 190886 53100
rect 530578 53088 530584 53100
rect 190880 53060 530584 53088
rect 190880 53048 190886 53060
rect 530578 53048 530584 53060
rect 530636 53048 530642 53100
rect 119246 52980 119252 53032
rect 119304 53020 119310 53032
rect 240134 53020 240140 53032
rect 119304 52992 240140 53020
rect 119304 52980 119310 52992
rect 240134 52980 240140 52992
rect 240192 52980 240198 53032
rect 116578 52912 116584 52964
rect 116636 52952 116642 52964
rect 229094 52952 229100 52964
rect 116636 52924 229100 52952
rect 116636 52912 116642 52924
rect 229094 52912 229100 52924
rect 229152 52912 229158 52964
rect 115842 52844 115848 52896
rect 115900 52884 115906 52896
rect 226334 52884 226340 52896
rect 115900 52856 226340 52884
rect 115900 52844 115906 52856
rect 226334 52844 226340 52856
rect 226392 52844 226398 52896
rect 123478 52776 123484 52828
rect 123536 52816 123542 52828
rect 233234 52816 233240 52828
rect 123536 52788 233240 52816
rect 123536 52776 123542 52788
rect 233234 52776 233240 52788
rect 233292 52776 233298 52828
rect 142890 52708 142896 52760
rect 142948 52748 142954 52760
rect 235994 52748 236000 52760
rect 142948 52720 236000 52748
rect 142948 52708 142954 52720
rect 235994 52708 236000 52720
rect 236052 52708 236058 52760
rect 156138 52640 156144 52692
rect 156196 52680 156202 52692
rect 160186 52680 160192 52692
rect 156196 52652 160192 52680
rect 156196 52640 156202 52652
rect 160186 52640 160192 52652
rect 160244 52640 160250 52692
rect 121914 52368 121920 52420
rect 121972 52408 121978 52420
rect 251174 52408 251180 52420
rect 121972 52380 251180 52408
rect 121972 52368 121978 52380
rect 251174 52368 251180 52380
rect 251232 52368 251238 52420
rect 122742 52300 122748 52352
rect 122800 52340 122806 52352
rect 253934 52340 253940 52352
rect 122800 52312 253940 52340
rect 122800 52300 122806 52312
rect 253934 52300 253940 52312
rect 253992 52300 253998 52352
rect 142798 52232 142804 52284
rect 142856 52272 142862 52284
rect 335354 52272 335360 52284
rect 142856 52244 335360 52272
rect 142856 52232 142862 52244
rect 335354 52232 335360 52244
rect 335412 52232 335418 52284
rect 143718 52164 143724 52216
rect 143776 52204 143782 52216
rect 339494 52204 339500 52216
rect 143776 52176 339500 52204
rect 143776 52164 143782 52176
rect 339494 52164 339500 52176
rect 339552 52164 339558 52216
rect 143534 52096 143540 52148
rect 143592 52136 143598 52148
rect 342254 52136 342260 52148
rect 143592 52108 342260 52136
rect 143592 52096 143598 52108
rect 342254 52096 342260 52108
rect 342312 52096 342318 52148
rect 145466 52028 145472 52080
rect 145524 52068 145530 52080
rect 346394 52068 346400 52080
rect 145524 52040 346400 52068
rect 145524 52028 145530 52040
rect 346394 52028 346400 52040
rect 346452 52028 346458 52080
rect 148134 51960 148140 52012
rect 148192 52000 148198 52012
rect 357526 52000 357532 52012
rect 148192 51972 357532 52000
rect 148192 51960 148198 51972
rect 357526 51960 357532 51972
rect 357584 51960 357590 52012
rect 149882 51892 149888 51944
rect 149940 51932 149946 51944
rect 364334 51932 364340 51944
rect 149940 51904 364340 51932
rect 149940 51892 149946 51904
rect 364334 51892 364340 51904
rect 364392 51892 364398 51944
rect 168374 51824 168380 51876
rect 168432 51864 168438 51876
rect 436738 51864 436744 51876
rect 168432 51836 436744 51864
rect 168432 51824 168438 51836
rect 436738 51824 436744 51836
rect 436796 51824 436802 51876
rect 192110 51756 192116 51808
rect 192168 51796 192174 51808
rect 535454 51796 535460 51808
rect 192168 51768 535460 51796
rect 192168 51756 192174 51768
rect 535454 51756 535460 51768
rect 535512 51756 535518 51808
rect 193214 51688 193220 51740
rect 193272 51728 193278 51740
rect 542354 51728 542360 51740
rect 193272 51700 542360 51728
rect 193272 51688 193278 51700
rect 542354 51688 542360 51700
rect 542412 51688 542418 51740
rect 143902 51620 143908 51672
rect 143960 51660 143966 51672
rect 247034 51660 247040 51672
rect 143960 51632 247040 51660
rect 143960 51620 143966 51632
rect 247034 51620 247040 51632
rect 247092 51620 247098 51672
rect 177114 51348 177120 51400
rect 177172 51388 177178 51400
rect 177942 51388 177948 51400
rect 177172 51360 177948 51388
rect 177172 51348 177178 51360
rect 177942 51348 177948 51360
rect 178000 51348 178006 51400
rect 172790 51008 172796 51060
rect 172848 51048 172854 51060
rect 432598 51048 432604 51060
rect 172848 51020 432604 51048
rect 172848 51008 172854 51020
rect 432598 51008 432604 51020
rect 432656 51008 432662 51060
rect 169754 50940 169760 50992
rect 169812 50980 169818 50992
rect 445754 50980 445760 50992
rect 169812 50952 445760 50980
rect 169812 50940 169818 50952
rect 445754 50940 445760 50952
rect 445812 50940 445818 50992
rect 169846 50872 169852 50924
rect 169904 50912 169910 50924
rect 448514 50912 448520 50924
rect 169904 50884 448520 50912
rect 169904 50872 169910 50884
rect 448514 50872 448520 50884
rect 448572 50872 448578 50924
rect 172606 50804 172612 50856
rect 172664 50844 172670 50856
rect 456794 50844 456800 50856
rect 172664 50816 456800 50844
rect 172664 50804 172670 50816
rect 456794 50804 456800 50816
rect 456852 50804 456858 50856
rect 174262 50736 174268 50788
rect 174320 50776 174326 50788
rect 463694 50776 463700 50788
rect 174320 50748 463700 50776
rect 174320 50736 174326 50748
rect 463694 50736 463700 50748
rect 463752 50736 463758 50788
rect 196434 50668 196440 50720
rect 196492 50708 196498 50720
rect 533338 50708 533344 50720
rect 196492 50680 533344 50708
rect 196492 50668 196498 50680
rect 533338 50668 533344 50680
rect 533396 50668 533402 50720
rect 194594 50600 194600 50652
rect 194652 50640 194658 50652
rect 537478 50640 537484 50652
rect 194652 50612 537484 50640
rect 194652 50600 194658 50612
rect 537478 50600 537484 50612
rect 537536 50600 537542 50652
rect 197538 50532 197544 50584
rect 197596 50572 197602 50584
rect 544378 50572 544384 50584
rect 197596 50544 544384 50572
rect 197596 50532 197602 50544
rect 544378 50532 544384 50544
rect 544436 50532 544442 50584
rect 194686 50464 194692 50516
rect 194744 50504 194750 50516
rect 194744 50476 199976 50504
rect 194744 50464 194750 50476
rect 199194 50396 199200 50448
rect 199252 50436 199258 50448
rect 199948 50436 199976 50476
rect 200022 50464 200028 50516
rect 200080 50504 200086 50516
rect 539594 50504 539600 50516
rect 200080 50476 539600 50504
rect 200080 50464 200086 50476
rect 539594 50464 539600 50476
rect 539652 50464 539658 50516
rect 546494 50436 546500 50448
rect 199252 50408 199884 50436
rect 199948 50408 546500 50436
rect 199252 50396 199258 50408
rect 106366 50328 106372 50380
rect 106424 50368 106430 50380
rect 107562 50368 107568 50380
rect 106424 50340 107568 50368
rect 106424 50328 106430 50340
rect 107562 50328 107568 50340
rect 107620 50328 107626 50380
rect 107654 50328 107660 50380
rect 107712 50368 107718 50380
rect 108942 50368 108948 50380
rect 107712 50340 108948 50368
rect 107712 50328 107718 50340
rect 108942 50328 108948 50340
rect 109000 50328 109006 50380
rect 109034 50328 109040 50380
rect 109092 50368 109098 50380
rect 110138 50368 110144 50380
rect 109092 50340 110144 50368
rect 109092 50328 109098 50340
rect 110138 50328 110144 50340
rect 110196 50328 110202 50380
rect 130102 50328 130108 50380
rect 130160 50368 130166 50380
rect 130930 50368 130936 50380
rect 130160 50340 130936 50368
rect 130160 50328 130166 50340
rect 130930 50328 130936 50340
rect 130988 50328 130994 50380
rect 135254 50328 135260 50380
rect 135312 50368 135318 50380
rect 136450 50368 136456 50380
rect 135312 50340 136456 50368
rect 135312 50328 135318 50340
rect 136450 50328 136456 50340
rect 136508 50328 136514 50380
rect 187694 50328 187700 50380
rect 187752 50368 187758 50380
rect 188798 50368 188804 50380
rect 187752 50340 188804 50368
rect 187752 50328 187758 50340
rect 188798 50328 188804 50340
rect 188856 50328 188862 50380
rect 196066 50328 196072 50380
rect 196124 50368 196130 50380
rect 197170 50368 197176 50380
rect 196124 50340 197176 50368
rect 196124 50328 196130 50340
rect 197170 50328 197176 50340
rect 197228 50328 197234 50380
rect 198734 50328 198740 50380
rect 198792 50368 198798 50380
rect 199746 50368 199752 50380
rect 198792 50340 199752 50368
rect 198792 50328 198798 50340
rect 199746 50328 199752 50340
rect 199804 50328 199810 50380
rect 199856 50368 199884 50408
rect 546494 50396 546500 50408
rect 546552 50396 546558 50448
rect 564434 50368 564440 50380
rect 199856 50340 564440 50368
rect 564434 50328 564440 50340
rect 564492 50328 564498 50380
rect 147674 50260 147680 50312
rect 147732 50300 147738 50312
rect 360194 50300 360200 50312
rect 147732 50272 360200 50300
rect 147732 50260 147738 50272
rect 360194 50260 360200 50272
rect 360252 50260 360258 50312
rect 137922 50192 137928 50244
rect 137980 50232 137986 50244
rect 280154 50232 280160 50244
rect 137980 50204 280160 50232
rect 137980 50192 137986 50204
rect 280154 50192 280160 50204
rect 280212 50192 280218 50244
rect 192202 50124 192208 50176
rect 192260 50164 192266 50176
rect 200022 50164 200028 50176
rect 192260 50136 200028 50164
rect 192260 50124 192266 50136
rect 200022 50124 200028 50136
rect 200080 50124 200086 50176
rect 200114 50124 200120 50176
rect 200172 50164 200178 50176
rect 201310 50164 201316 50176
rect 200172 50136 201316 50164
rect 200172 50124 200178 50136
rect 201310 50124 201316 50136
rect 201368 50124 201374 50176
rect 201678 50124 201684 50176
rect 201736 50164 201742 50176
rect 202598 50164 202604 50176
rect 201736 50136 202604 50164
rect 201736 50124 201742 50136
rect 202598 50124 202604 50136
rect 202656 50124 202662 50176
rect 201586 50056 201592 50108
rect 201644 50096 201650 50108
rect 202690 50096 202696 50108
rect 201644 50068 202696 50096
rect 201644 50056 201650 50068
rect 202690 50056 202696 50068
rect 202748 50056 202754 50108
rect 151814 49308 151820 49360
rect 151872 49348 151878 49360
rect 291194 49348 291200 49360
rect 151872 49320 291200 49348
rect 151872 49308 151878 49320
rect 291194 49308 291200 49320
rect 291252 49308 291258 49360
rect 178126 49240 178132 49292
rect 178184 49280 178190 49292
rect 329834 49280 329840 49292
rect 178184 49252 329840 49280
rect 178184 49240 178190 49252
rect 329834 49240 329840 49252
rect 329892 49240 329898 49292
rect 156690 49172 156696 49224
rect 156748 49212 156754 49224
rect 322934 49212 322940 49224
rect 156748 49184 322940 49212
rect 156748 49172 156754 49184
rect 322934 49172 322940 49184
rect 322992 49172 322998 49224
rect 141326 49104 141332 49156
rect 141384 49144 141390 49156
rect 311894 49144 311900 49156
rect 141384 49116 311900 49144
rect 141384 49104 141390 49116
rect 311894 49104 311900 49116
rect 311952 49104 311958 49156
rect 156046 49036 156052 49088
rect 156104 49076 156110 49088
rect 340874 49076 340880 49088
rect 156104 49048 340880 49076
rect 156104 49036 156110 49048
rect 340874 49036 340880 49048
rect 340932 49036 340938 49088
rect 197354 48968 197360 49020
rect 197412 49008 197418 49020
rect 560294 49008 560300 49020
rect 197412 48980 560300 49008
rect 197412 48968 197418 48980
rect 560294 48968 560300 48980
rect 560352 48968 560358 49020
rect 242342 46860 242348 46912
rect 242400 46900 242406 46912
rect 579982 46900 579988 46912
rect 242400 46872 579988 46900
rect 242400 46860 242406 46872
rect 579982 46860 579988 46872
rect 580040 46860 580046 46912
rect 124398 46316 124404 46368
rect 124456 46356 124462 46368
rect 125502 46356 125508 46368
rect 124456 46328 125508 46356
rect 124456 46316 124462 46328
rect 125502 46316 125508 46328
rect 125560 46316 125566 46368
rect 124582 46248 124588 46300
rect 124640 46288 124646 46300
rect 125318 46288 125324 46300
rect 124640 46260 125324 46288
rect 124640 46248 124646 46260
rect 125318 46248 125324 46260
rect 125376 46248 125382 46300
rect 125778 46248 125784 46300
rect 125836 46288 125842 46300
rect 126882 46288 126888 46300
rect 125836 46260 126888 46288
rect 125836 46248 125842 46260
rect 126882 46248 126888 46260
rect 126940 46248 126946 46300
rect 126974 46248 126980 46300
rect 127032 46288 127038 46300
rect 128262 46288 128268 46300
rect 127032 46260 128268 46288
rect 127032 46248 127038 46260
rect 128262 46248 128268 46260
rect 128320 46248 128326 46300
rect 118878 46180 118884 46232
rect 118936 46220 118942 46232
rect 119890 46220 119896 46232
rect 118936 46192 119896 46220
rect 118936 46180 118942 46192
rect 119890 46180 119896 46192
rect 119948 46180 119954 46232
rect 120074 46180 120080 46232
rect 120132 46220 120138 46232
rect 121362 46220 121368 46232
rect 120132 46192 121368 46220
rect 120132 46180 120138 46192
rect 121362 46180 121368 46192
rect 121420 46180 121426 46232
rect 122834 46180 122840 46232
rect 122892 46220 122898 46232
rect 124122 46220 124128 46232
rect 122892 46192 124128 46220
rect 122892 46180 122898 46192
rect 124122 46180 124128 46192
rect 124180 46180 124186 46232
rect 124490 46180 124496 46232
rect 124548 46220 124554 46232
rect 125226 46220 125232 46232
rect 124548 46192 125232 46220
rect 124548 46180 124554 46192
rect 125226 46180 125232 46192
rect 125284 46180 125290 46232
rect 125594 46180 125600 46232
rect 125652 46220 125658 46232
rect 126698 46220 126704 46232
rect 125652 46192 126704 46220
rect 125652 46180 125658 46192
rect 126698 46180 126704 46192
rect 126756 46180 126762 46232
rect 127066 46180 127072 46232
rect 127124 46220 127130 46232
rect 128078 46220 128084 46232
rect 127124 46192 128084 46220
rect 127124 46180 127130 46192
rect 128078 46180 128084 46192
rect 128136 46180 128142 46232
rect 124306 46112 124312 46164
rect 124364 46152 124370 46164
rect 125410 46152 125416 46164
rect 124364 46124 125416 46152
rect 124364 46112 124370 46124
rect 125410 46112 125416 46124
rect 125468 46112 125474 46164
rect 119338 45364 119344 45416
rect 119396 45404 119402 45416
rect 119706 45404 119712 45416
rect 119396 45376 119712 45404
rect 119396 45364 119402 45376
rect 119706 45364 119712 45376
rect 119764 45364 119770 45416
rect 2866 33056 2872 33108
rect 2924 33096 2930 33108
rect 15838 33096 15844 33108
rect 2924 33068 15844 33096
rect 2924 33056 2930 33068
rect 15838 33056 15844 33068
rect 15896 33056 15902 33108
rect 130378 24080 130384 24132
rect 130436 24120 130442 24132
rect 242894 24120 242900 24132
rect 130436 24092 242900 24120
rect 130436 24080 130442 24092
rect 242894 24080 242900 24092
rect 242952 24080 242958 24132
rect 3418 20612 3424 20664
rect 3476 20652 3482 20664
rect 29638 20652 29644 20664
rect 3476 20624 29644 20652
rect 3476 20612 3482 20624
rect 29638 20612 29644 20624
rect 29696 20612 29702 20664
rect 55674 20612 55680 20664
rect 55732 20652 55738 20664
rect 580074 20652 580080 20664
rect 55732 20624 580080 20652
rect 55732 20612 55738 20624
rect 580074 20612 580080 20624
rect 580132 20612 580138 20664
rect 204898 20068 204904 20120
rect 204956 20108 204962 20120
rect 440234 20108 440240 20120
rect 204956 20080 440240 20108
rect 204956 20068 204962 20080
rect 440234 20068 440240 20080
rect 440292 20068 440298 20120
rect 209038 20000 209044 20052
rect 209096 20040 209102 20052
rect 454034 20040 454040 20052
rect 209096 20012 454040 20040
rect 209096 20000 209102 20012
rect 454034 20000 454040 20012
rect 454092 20000 454098 20052
rect 216030 19932 216036 19984
rect 216088 19972 216094 19984
rect 467834 19972 467840 19984
rect 216088 19944 467840 19972
rect 216088 19932 216094 19944
rect 467834 19932 467840 19944
rect 467892 19932 467898 19984
rect 115658 18844 115664 18896
rect 115716 18884 115722 18896
rect 224954 18884 224960 18896
rect 115716 18856 224960 18884
rect 115716 18844 115722 18856
rect 224954 18844 224960 18856
rect 225012 18844 225018 18896
rect 164878 18776 164884 18828
rect 164936 18816 164942 18828
rect 318794 18816 318800 18828
rect 164936 18788 318800 18816
rect 164936 18776 164942 18788
rect 318794 18776 318800 18788
rect 318852 18776 318858 18828
rect 160738 18708 160744 18760
rect 160796 18748 160802 18760
rect 325694 18748 325700 18760
rect 160796 18720 325700 18748
rect 160796 18708 160802 18720
rect 325694 18708 325700 18720
rect 325752 18708 325758 18760
rect 170398 18640 170404 18692
rect 170456 18680 170462 18692
rect 361574 18680 361580 18692
rect 170456 18652 361580 18680
rect 170456 18640 170462 18652
rect 361574 18640 361580 18652
rect 361632 18640 361638 18692
rect 213270 18572 213276 18624
rect 213328 18612 213334 18624
rect 460934 18612 460940 18624
rect 213328 18584 460940 18612
rect 213328 18572 213334 18584
rect 460934 18572 460940 18584
rect 460992 18572 460998 18624
rect 126514 17892 126520 17944
rect 126572 17932 126578 17944
rect 269114 17932 269120 17944
rect 126572 17904 269120 17932
rect 126572 17892 126578 17904
rect 269114 17892 269120 17904
rect 269172 17892 269178 17944
rect 127894 17824 127900 17876
rect 127952 17864 127958 17876
rect 273254 17864 273260 17876
rect 127952 17836 273260 17864
rect 127952 17824 127958 17836
rect 273254 17824 273260 17836
rect 273312 17824 273318 17876
rect 127986 17756 127992 17808
rect 128044 17796 128050 17808
rect 276014 17796 276020 17808
rect 128044 17768 276020 17796
rect 128044 17756 128050 17768
rect 276014 17756 276020 17768
rect 276072 17756 276078 17808
rect 130746 17688 130752 17740
rect 130804 17728 130810 17740
rect 287054 17728 287060 17740
rect 130804 17700 287060 17728
rect 130804 17688 130810 17700
rect 287054 17688 287060 17700
rect 287112 17688 287118 17740
rect 184198 17620 184204 17672
rect 184256 17660 184262 17672
rect 343634 17660 343640 17672
rect 184256 17632 343640 17660
rect 184256 17620 184262 17632
rect 343634 17620 343640 17632
rect 343692 17620 343698 17672
rect 133598 17552 133604 17604
rect 133656 17592 133662 17604
rect 298094 17592 298100 17604
rect 133656 17564 298100 17592
rect 133656 17552 133662 17564
rect 298094 17552 298100 17564
rect 298152 17552 298158 17604
rect 134978 17484 134984 17536
rect 135036 17524 135042 17536
rect 300854 17524 300860 17536
rect 135036 17496 300860 17524
rect 135036 17484 135042 17496
rect 300854 17484 300860 17496
rect 300912 17484 300918 17536
rect 136266 17416 136272 17468
rect 136324 17456 136330 17468
rect 307754 17456 307760 17468
rect 136324 17428 307760 17456
rect 136324 17416 136330 17428
rect 307754 17416 307760 17428
rect 307812 17416 307818 17468
rect 137738 17348 137744 17400
rect 137796 17388 137802 17400
rect 316126 17388 316132 17400
rect 137796 17360 316132 17388
rect 137796 17348 137802 17360
rect 316126 17348 316132 17360
rect 316184 17348 316190 17400
rect 144178 17280 144184 17332
rect 144236 17320 144242 17332
rect 332594 17320 332600 17332
rect 144236 17292 332600 17320
rect 144236 17280 144242 17292
rect 332594 17280 332600 17292
rect 332652 17280 332658 17332
rect 141878 17212 141884 17264
rect 141936 17252 141942 17264
rect 332686 17252 332692 17264
rect 141936 17224 332692 17252
rect 141936 17212 141942 17224
rect 332686 17212 332692 17224
rect 332744 17212 332750 17264
rect 126606 17144 126612 17196
rect 126664 17184 126670 17196
rect 266354 17184 266360 17196
rect 126664 17156 266360 17184
rect 126664 17144 126670 17156
rect 266354 17144 266360 17156
rect 266412 17144 266418 17196
rect 125134 17076 125140 17128
rect 125192 17116 125198 17128
rect 262214 17116 262220 17128
rect 125192 17088 262220 17116
rect 125192 17076 125198 17088
rect 262214 17076 262220 17088
rect 262272 17076 262278 17128
rect 119798 16532 119804 16584
rect 119856 16572 119862 16584
rect 238110 16572 238116 16584
rect 119856 16544 238116 16572
rect 119856 16532 119862 16544
rect 238110 16532 238116 16544
rect 238168 16532 238174 16584
rect 119706 16464 119712 16516
rect 119764 16504 119770 16516
rect 241698 16504 241704 16516
rect 119764 16476 241704 16504
rect 119764 16464 119770 16476
rect 241698 16464 241704 16476
rect 241756 16464 241762 16516
rect 121178 16396 121184 16448
rect 121236 16436 121242 16448
rect 245194 16436 245200 16448
rect 121236 16408 245200 16436
rect 121236 16396 121242 16408
rect 245194 16396 245200 16408
rect 245252 16396 245258 16448
rect 121270 16328 121276 16380
rect 121328 16368 121334 16380
rect 248782 16368 248788 16380
rect 121328 16340 248788 16368
rect 121328 16328 121334 16340
rect 248782 16328 248788 16340
rect 248840 16328 248846 16380
rect 122558 16260 122564 16312
rect 122616 16300 122622 16312
rect 252370 16300 252376 16312
rect 122616 16272 252376 16300
rect 122616 16260 122622 16272
rect 252370 16260 252376 16272
rect 252428 16260 252434 16312
rect 123846 16192 123852 16244
rect 123904 16232 123910 16244
rect 255866 16232 255872 16244
rect 123904 16204 255872 16232
rect 123904 16192 123910 16204
rect 255866 16192 255872 16204
rect 255924 16192 255930 16244
rect 123938 16124 123944 16176
rect 123996 16164 124002 16176
rect 259454 16164 259460 16176
rect 123996 16136 259460 16164
rect 123996 16124 124002 16136
rect 259454 16124 259460 16136
rect 259512 16124 259518 16176
rect 199746 16056 199752 16108
rect 199804 16096 199810 16108
rect 568022 16096 568028 16108
rect 199804 16068 568028 16096
rect 199804 16056 199810 16068
rect 568022 16056 568028 16068
rect 568080 16056 568086 16108
rect 201126 15988 201132 16040
rect 201184 16028 201190 16040
rect 571518 16028 571524 16040
rect 201184 16000 571524 16028
rect 201184 15988 201190 16000
rect 571518 15988 571524 16000
rect 571576 15988 571582 16040
rect 202506 15920 202512 15972
rect 202564 15960 202570 15972
rect 575106 15960 575112 15972
rect 202564 15932 575112 15960
rect 202564 15920 202570 15932
rect 575106 15920 575112 15932
rect 575164 15920 575170 15972
rect 90726 15852 90732 15904
rect 90784 15892 90790 15904
rect 123570 15892 123576 15904
rect 90784 15864 123576 15892
rect 90784 15852 90790 15864
rect 123570 15852 123576 15864
rect 123628 15852 123634 15904
rect 202414 15852 202420 15904
rect 202472 15892 202478 15904
rect 578602 15892 578608 15904
rect 202472 15864 578608 15892
rect 202472 15852 202478 15864
rect 578602 15852 578608 15864
rect 578660 15852 578666 15904
rect 118510 15784 118516 15836
rect 118568 15824 118574 15836
rect 234614 15824 234620 15836
rect 118568 15796 234620 15824
rect 118568 15784 118574 15796
rect 234614 15784 234620 15796
rect 234672 15784 234678 15836
rect 117038 15716 117044 15768
rect 117096 15756 117102 15768
rect 231026 15756 231032 15768
rect 117096 15728 231032 15756
rect 117096 15716 117102 15728
rect 231026 15716 231032 15728
rect 231084 15716 231090 15768
rect 117130 15648 117136 15700
rect 117188 15688 117194 15700
rect 227530 15688 227536 15700
rect 117188 15660 227536 15688
rect 117188 15648 117194 15660
rect 227530 15648 227536 15660
rect 227588 15648 227594 15700
rect 115750 15580 115756 15632
rect 115808 15620 115814 15632
rect 223942 15620 223948 15632
rect 115808 15592 223948 15620
rect 115808 15580 115814 15592
rect 223942 15580 223948 15592
rect 224000 15580 224006 15632
rect 114278 15512 114284 15564
rect 114336 15552 114342 15564
rect 219986 15552 219992 15564
rect 114336 15524 219992 15552
rect 114336 15512 114342 15524
rect 219986 15512 219992 15524
rect 220044 15512 220050 15564
rect 114370 15444 114376 15496
rect 114428 15484 114434 15496
rect 216858 15484 216864 15496
rect 114428 15456 216864 15484
rect 114428 15444 114434 15456
rect 216858 15444 216864 15456
rect 216916 15444 216922 15496
rect 112898 15376 112904 15428
rect 112956 15416 112962 15428
rect 213086 15416 213092 15428
rect 112956 15388 213092 15416
rect 112956 15376 112962 15388
rect 213086 15376 213092 15388
rect 213144 15376 213150 15428
rect 111518 15308 111524 15360
rect 111576 15348 111582 15360
rect 209866 15348 209872 15360
rect 111576 15320 209872 15348
rect 111576 15308 111582 15320
rect 209866 15308 209872 15320
rect 209924 15308 209930 15360
rect 183278 15104 183284 15156
rect 183336 15144 183342 15156
rect 497090 15144 497096 15156
rect 183336 15116 497096 15144
rect 183336 15104 183342 15116
rect 497090 15104 497096 15116
rect 497148 15104 497154 15156
rect 183186 15036 183192 15088
rect 183244 15076 183250 15088
rect 500586 15076 500592 15088
rect 183244 15048 500592 15076
rect 183244 15036 183250 15048
rect 500586 15036 500592 15048
rect 500644 15036 500650 15088
rect 184566 14968 184572 15020
rect 184624 15008 184630 15020
rect 504174 15008 504180 15020
rect 184624 14980 504180 15008
rect 184624 14968 184630 14980
rect 504174 14968 504180 14980
rect 504232 14968 504238 15020
rect 186038 14900 186044 14952
rect 186096 14940 186102 14952
rect 507670 14940 507676 14952
rect 186096 14912 507676 14940
rect 186096 14900 186102 14912
rect 507670 14900 507676 14912
rect 507728 14900 507734 14952
rect 186130 14832 186136 14884
rect 186188 14872 186194 14884
rect 511258 14872 511264 14884
rect 186188 14844 511264 14872
rect 186188 14832 186194 14844
rect 511258 14832 511264 14844
rect 511316 14832 511322 14884
rect 187418 14764 187424 14816
rect 187476 14804 187482 14816
rect 514754 14804 514760 14816
rect 187476 14776 514760 14804
rect 187476 14764 187482 14776
rect 514754 14764 514760 14776
rect 514812 14764 514818 14816
rect 188798 14696 188804 14748
rect 188856 14736 188862 14748
rect 518342 14736 518348 14748
rect 188856 14708 518348 14736
rect 188856 14696 188862 14708
rect 518342 14696 518348 14708
rect 518400 14696 518406 14748
rect 188706 14628 188712 14680
rect 188764 14668 188770 14680
rect 521838 14668 521844 14680
rect 188764 14640 521844 14668
rect 188764 14628 188770 14640
rect 521838 14628 521844 14640
rect 521896 14628 521902 14680
rect 190270 14560 190276 14612
rect 190328 14600 190334 14612
rect 525426 14600 525432 14612
rect 190328 14572 525432 14600
rect 190328 14560 190334 14572
rect 525426 14560 525432 14572
rect 525484 14560 525490 14612
rect 190178 14492 190184 14544
rect 190236 14532 190242 14544
rect 529014 14532 529020 14544
rect 190236 14504 529020 14532
rect 190236 14492 190242 14504
rect 529014 14492 529020 14504
rect 529072 14492 529078 14544
rect 191558 14424 191564 14476
rect 191616 14464 191622 14476
rect 532510 14464 532516 14476
rect 191616 14436 532516 14464
rect 191616 14424 191622 14436
rect 532510 14424 532516 14436
rect 532568 14424 532574 14476
rect 181990 14356 181996 14408
rect 182048 14396 182054 14408
rect 493502 14396 493508 14408
rect 182048 14368 493508 14396
rect 182048 14356 182054 14368
rect 493502 14356 493508 14368
rect 493560 14356 493566 14408
rect 181898 14288 181904 14340
rect 181956 14328 181962 14340
rect 489914 14328 489920 14340
rect 181956 14300 489920 14328
rect 181956 14288 181962 14300
rect 489914 14288 489920 14300
rect 489972 14288 489978 14340
rect 180518 14220 180524 14272
rect 180576 14260 180582 14272
rect 486418 14260 486424 14272
rect 180576 14232 486424 14260
rect 180576 14220 180582 14232
rect 486418 14220 486424 14232
rect 486476 14220 486482 14272
rect 179138 14152 179144 14204
rect 179196 14192 179202 14204
rect 481634 14192 481640 14204
rect 179196 14164 481640 14192
rect 179196 14152 179202 14164
rect 481634 14152 481640 14164
rect 481692 14152 481698 14204
rect 177666 14084 177672 14136
rect 177724 14124 177730 14136
rect 478138 14124 478144 14136
rect 177724 14096 478144 14124
rect 177724 14084 177730 14096
rect 478138 14084 478144 14096
rect 478196 14084 478202 14136
rect 177574 14016 177580 14068
rect 177632 14056 177638 14068
rect 473354 14056 473360 14068
rect 177632 14028 473360 14056
rect 177632 14016 177638 14028
rect 473354 14016 473360 14028
rect 473412 14016 473418 14068
rect 176470 13948 176476 14000
rect 176528 13988 176534 14000
rect 471054 13988 471060 14000
rect 176528 13960 471060 13988
rect 176528 13948 176534 13960
rect 471054 13948 471060 13960
rect 471112 13948 471118 14000
rect 176378 13880 176384 13932
rect 176436 13920 176442 13932
rect 467466 13920 467472 13932
rect 176436 13892 467472 13920
rect 176436 13880 176442 13892
rect 467466 13880 467472 13892
rect 467524 13880 467530 13932
rect 158346 13744 158352 13796
rect 158404 13784 158410 13796
rect 396534 13784 396540 13796
rect 158404 13756 396540 13784
rect 158404 13744 158410 13756
rect 396534 13744 396540 13756
rect 396592 13744 396598 13796
rect 158254 13676 158260 13728
rect 158312 13716 158318 13728
rect 398834 13716 398840 13728
rect 158312 13688 398840 13716
rect 158312 13676 158318 13688
rect 398834 13676 398840 13688
rect 398892 13676 398898 13728
rect 159910 13608 159916 13660
rect 159968 13648 159974 13660
rect 403618 13648 403624 13660
rect 159968 13620 403624 13648
rect 159968 13608 159974 13620
rect 403618 13608 403624 13620
rect 403676 13608 403682 13660
rect 161014 13540 161020 13592
rect 161072 13580 161078 13592
rect 407206 13580 407212 13592
rect 161072 13552 407212 13580
rect 161072 13540 161078 13552
rect 407206 13540 407212 13552
rect 407264 13540 407270 13592
rect 161198 13472 161204 13524
rect 161256 13512 161262 13524
rect 410794 13512 410800 13524
rect 161256 13484 410800 13512
rect 161256 13472 161262 13484
rect 410794 13472 410800 13484
rect 410852 13472 410858 13524
rect 162670 13404 162676 13456
rect 162728 13444 162734 13456
rect 414290 13444 414296 13456
rect 162728 13416 414296 13444
rect 162728 13404 162734 13416
rect 414290 13404 414296 13416
rect 414348 13404 414354 13456
rect 164050 13336 164056 13388
rect 164108 13376 164114 13388
rect 417418 13376 417424 13388
rect 164108 13348 417424 13376
rect 164108 13336 164114 13348
rect 417418 13336 417424 13348
rect 417476 13336 417482 13388
rect 163958 13268 163964 13320
rect 164016 13308 164022 13320
rect 421374 13308 421380 13320
rect 164016 13280 421380 13308
rect 164016 13268 164022 13280
rect 421374 13268 421380 13280
rect 421432 13268 421438 13320
rect 165430 13200 165436 13252
rect 165488 13240 165494 13252
rect 423766 13240 423772 13252
rect 165488 13212 423772 13240
rect 165488 13200 165494 13212
rect 423766 13200 423772 13212
rect 423824 13200 423830 13252
rect 166718 13132 166724 13184
rect 166776 13172 166782 13184
rect 428458 13172 428464 13184
rect 166776 13144 428464 13172
rect 166776 13132 166782 13144
rect 428458 13132 428464 13144
rect 428516 13132 428522 13184
rect 166810 13064 166816 13116
rect 166868 13104 166874 13116
rect 432046 13104 432052 13116
rect 166868 13076 432052 13104
rect 166868 13064 166874 13076
rect 432046 13064 432052 13076
rect 432104 13064 432110 13116
rect 156966 12996 156972 13048
rect 157024 13036 157030 13048
rect 393038 13036 393044 13048
rect 157024 13008 393044 13036
rect 157024 12996 157030 13008
rect 393038 12996 393044 13008
rect 393096 12996 393102 13048
rect 157058 12928 157064 12980
rect 157116 12968 157122 12980
rect 389450 12968 389456 12980
rect 157116 12940 389456 12968
rect 157116 12928 157122 12940
rect 389450 12928 389456 12940
rect 389508 12928 389514 12980
rect 155586 12860 155592 12912
rect 155644 12900 155650 12912
rect 385954 12900 385960 12912
rect 155644 12872 385960 12900
rect 155644 12860 155650 12872
rect 385954 12860 385960 12872
rect 386012 12860 386018 12912
rect 154298 12792 154304 12844
rect 154356 12832 154362 12844
rect 382366 12832 382372 12844
rect 154356 12804 382372 12832
rect 154356 12792 154362 12804
rect 382366 12792 382372 12804
rect 382424 12792 382430 12844
rect 154206 12724 154212 12776
rect 154264 12764 154270 12776
rect 378870 12764 378876 12776
rect 154264 12736 378876 12764
rect 154264 12724 154270 12736
rect 378870 12724 378876 12736
rect 378928 12724 378934 12776
rect 152734 12656 152740 12708
rect 152792 12696 152798 12708
rect 373994 12696 374000 12708
rect 152792 12668 374000 12696
rect 152792 12656 152798 12668
rect 373994 12656 374000 12668
rect 374052 12656 374058 12708
rect 151354 12588 151360 12640
rect 151412 12628 151418 12640
rect 368198 12628 368204 12640
rect 151412 12600 368204 12628
rect 151412 12588 151418 12600
rect 368198 12588 368204 12600
rect 368256 12588 368262 12640
rect 132218 12384 132224 12436
rect 132276 12424 132282 12436
rect 293678 12424 293684 12436
rect 132276 12396 293684 12424
rect 132276 12384 132282 12396
rect 293678 12384 293684 12396
rect 293736 12384 293742 12436
rect 133690 12316 133696 12368
rect 133748 12356 133754 12368
rect 297266 12356 297272 12368
rect 133748 12328 297272 12356
rect 133748 12316 133754 12328
rect 297266 12316 297272 12328
rect 297324 12316 297330 12368
rect 134886 12248 134892 12300
rect 134944 12288 134950 12300
rect 299566 12288 299572 12300
rect 134944 12260 299572 12288
rect 134944 12248 134950 12260
rect 299566 12248 299572 12260
rect 299624 12248 299630 12300
rect 135070 12180 135076 12232
rect 135128 12220 135134 12232
rect 304350 12220 304356 12232
rect 135128 12192 304356 12220
rect 135128 12180 135134 12192
rect 304350 12180 304356 12192
rect 304408 12180 304414 12232
rect 136358 12112 136364 12164
rect 136416 12152 136422 12164
rect 307938 12152 307944 12164
rect 136416 12124 307944 12152
rect 136416 12112 136422 12124
rect 307938 12112 307944 12124
rect 307996 12112 308002 12164
rect 137830 12044 137836 12096
rect 137888 12084 137894 12096
rect 311434 12084 311440 12096
rect 137888 12056 311440 12084
rect 137888 12044 137894 12056
rect 311434 12044 311440 12056
rect 311492 12044 311498 12096
rect 137646 11976 137652 12028
rect 137704 12016 137710 12028
rect 315022 12016 315028 12028
rect 137704 11988 315028 12016
rect 137704 11976 137710 11988
rect 315022 11976 315028 11988
rect 315080 11976 315086 12028
rect 139118 11908 139124 11960
rect 139176 11948 139182 11960
rect 318518 11948 318524 11960
rect 139176 11920 318524 11948
rect 139176 11908 139182 11920
rect 318518 11908 318524 11920
rect 318576 11908 318582 11960
rect 140590 11840 140596 11892
rect 140648 11880 140654 11892
rect 322106 11880 322112 11892
rect 140648 11852 322112 11880
rect 140648 11840 140654 11852
rect 322106 11840 322112 11852
rect 322164 11840 322170 11892
rect 140682 11772 140688 11824
rect 140740 11812 140746 11824
rect 325602 11812 325608 11824
rect 140740 11784 325608 11812
rect 140740 11772 140746 11784
rect 325602 11772 325608 11784
rect 325660 11772 325666 11824
rect 141970 11704 141976 11756
rect 142028 11744 142034 11756
rect 329190 11744 329196 11756
rect 142028 11716 329196 11744
rect 142028 11704 142034 11716
rect 329190 11704 329196 11716
rect 329248 11704 329254 11756
rect 132126 11636 132132 11688
rect 132184 11676 132190 11688
rect 290182 11676 290188 11688
rect 132184 11648 290188 11676
rect 132184 11636 132190 11648
rect 290182 11636 290188 11648
rect 290240 11636 290246 11688
rect 130838 11568 130844 11620
rect 130896 11608 130902 11620
rect 286594 11608 286600 11620
rect 130896 11580 286600 11608
rect 130896 11568 130902 11580
rect 286594 11568 286600 11580
rect 286652 11568 286658 11620
rect 129458 11500 129464 11552
rect 129516 11540 129522 11552
rect 279510 11540 279516 11552
rect 129516 11512 279516 11540
rect 129516 11500 129522 11512
rect 279510 11500 279516 11512
rect 279568 11500 279574 11552
rect 128078 11432 128084 11484
rect 128136 11472 128142 11484
rect 276106 11472 276112 11484
rect 128136 11444 276112 11472
rect 128136 11432 128142 11444
rect 276106 11432 276112 11444
rect 276164 11432 276170 11484
rect 126698 11364 126704 11416
rect 126756 11404 126762 11416
rect 268838 11404 268844 11416
rect 126756 11376 268844 11404
rect 126756 11364 126762 11376
rect 268838 11364 268844 11376
rect 268896 11364 268902 11416
rect 125318 11296 125324 11348
rect 125376 11336 125382 11348
rect 265342 11336 265348 11348
rect 125376 11308 265348 11336
rect 125376 11296 125382 11308
rect 265342 11296 265348 11308
rect 265400 11296 265406 11348
rect 125226 11228 125232 11280
rect 125284 11268 125290 11280
rect 261754 11268 261760 11280
rect 125284 11240 261760 11268
rect 125284 11228 125290 11240
rect 261754 11228 261760 11240
rect 261812 11228 261818 11280
rect 124030 11160 124036 11212
rect 124088 11200 124094 11212
rect 258258 11200 258264 11212
rect 124088 11172 258264 11200
rect 124088 11160 124094 11172
rect 258258 11160 258264 11172
rect 258316 11160 258322 11212
rect 209774 11092 209780 11144
rect 209832 11132 209838 11144
rect 210970 11132 210976 11144
rect 209832 11104 210976 11132
rect 209832 11092 209838 11104
rect 210970 11092 210976 11104
rect 211028 11092 211034 11144
rect 194226 10956 194232 11008
rect 194284 10996 194290 11008
rect 541986 10996 541992 11008
rect 194284 10968 541992 10996
rect 194284 10956 194290 10968
rect 541986 10956 541992 10968
rect 542044 10956 542050 11008
rect 105998 10888 106004 10940
rect 106056 10928 106062 10940
rect 184934 10928 184940 10940
rect 106056 10900 184940 10928
rect 106056 10888 106062 10900
rect 184934 10888 184940 10900
rect 184992 10888 184998 10940
rect 194318 10888 194324 10940
rect 194376 10928 194382 10940
rect 545482 10928 545488 10940
rect 194376 10900 545488 10928
rect 194376 10888 194382 10900
rect 545482 10888 545488 10900
rect 545540 10888 545546 10940
rect 107194 10820 107200 10872
rect 107252 10860 107258 10872
rect 188522 10860 188528 10872
rect 107252 10832 188528 10860
rect 107252 10820 107258 10832
rect 188522 10820 188528 10832
rect 188580 10820 188586 10872
rect 195790 10820 195796 10872
rect 195848 10860 195854 10872
rect 547874 10860 547880 10872
rect 195848 10832 547880 10860
rect 195848 10820 195854 10832
rect 547874 10820 547880 10832
rect 547932 10820 547938 10872
rect 107286 10752 107292 10804
rect 107344 10792 107350 10804
rect 190822 10792 190828 10804
rect 107344 10764 190828 10792
rect 107344 10752 107350 10764
rect 190822 10752 190828 10764
rect 190880 10752 190886 10804
rect 196986 10752 196992 10804
rect 197044 10792 197050 10804
rect 552658 10792 552664 10804
rect 197044 10764 552664 10792
rect 197044 10752 197050 10764
rect 552658 10752 552664 10764
rect 552716 10752 552722 10804
rect 107378 10684 107384 10736
rect 107436 10724 107442 10736
rect 192018 10724 192024 10736
rect 107436 10696 192024 10724
rect 107436 10684 107442 10696
rect 192018 10684 192024 10696
rect 192076 10684 192082 10736
rect 197078 10684 197084 10736
rect 197136 10724 197142 10736
rect 556154 10724 556160 10736
rect 197136 10696 556160 10724
rect 197136 10684 197142 10696
rect 556154 10684 556160 10696
rect 556212 10684 556218 10736
rect 108758 10616 108764 10668
rect 108816 10656 108822 10668
rect 193214 10656 193220 10668
rect 108816 10628 193220 10656
rect 108816 10616 108822 10628
rect 193214 10616 193220 10628
rect 193272 10616 193278 10668
rect 198458 10616 198464 10668
rect 198516 10656 198522 10668
rect 559742 10656 559748 10668
rect 198516 10628 559748 10656
rect 198516 10616 198522 10628
rect 559742 10616 559748 10628
rect 559800 10616 559806 10668
rect 108666 10548 108672 10600
rect 108724 10588 108730 10600
rect 195606 10588 195612 10600
rect 108724 10560 195612 10588
rect 108724 10548 108730 10560
rect 195606 10548 195612 10560
rect 195664 10548 195670 10600
rect 199838 10548 199844 10600
rect 199896 10588 199902 10600
rect 563238 10588 563244 10600
rect 199896 10560 563244 10588
rect 199896 10548 199902 10560
rect 563238 10548 563244 10560
rect 563296 10548 563302 10600
rect 108850 10480 108856 10532
rect 108908 10520 108914 10532
rect 197906 10520 197912 10532
rect 108908 10492 197912 10520
rect 108908 10480 108914 10492
rect 197906 10480 197912 10492
rect 197964 10480 197970 10532
rect 199930 10480 199936 10532
rect 199988 10520 199994 10532
rect 566826 10520 566832 10532
rect 199988 10492 566832 10520
rect 199988 10480 199994 10492
rect 566826 10480 566832 10492
rect 566884 10480 566890 10532
rect 110138 10412 110144 10464
rect 110196 10452 110202 10464
rect 199102 10452 199108 10464
rect 110196 10424 199108 10452
rect 110196 10412 110202 10424
rect 199102 10412 199108 10424
rect 199160 10412 199166 10464
rect 201218 10412 201224 10464
rect 201276 10452 201282 10464
rect 570322 10452 570328 10464
rect 201276 10424 570328 10452
rect 201276 10412 201282 10424
rect 570322 10412 570328 10424
rect 570380 10412 570386 10464
rect 110230 10344 110236 10396
rect 110288 10384 110294 10396
rect 202690 10384 202696 10396
rect 110288 10356 202696 10384
rect 110288 10344 110294 10356
rect 202690 10344 202696 10356
rect 202748 10344 202754 10396
rect 202874 10344 202880 10396
rect 202932 10384 202938 10396
rect 572714 10384 572720 10396
rect 202932 10356 572720 10384
rect 202932 10344 202938 10356
rect 572714 10344 572720 10356
rect 572772 10344 572778 10396
rect 110046 10276 110052 10328
rect 110104 10316 110110 10328
rect 201586 10316 201592 10328
rect 110104 10288 201592 10316
rect 110104 10276 110110 10288
rect 201586 10276 201592 10288
rect 201644 10276 201650 10328
rect 202506 10276 202512 10328
rect 202564 10316 202570 10328
rect 577406 10316 577412 10328
rect 202564 10288 577412 10316
rect 202564 10276 202570 10288
rect 577406 10276 577412 10288
rect 577464 10276 577470 10328
rect 192938 10208 192944 10260
rect 192996 10248 193002 10260
rect 538398 10248 538404 10260
rect 192996 10220 538404 10248
rect 192996 10208 193002 10220
rect 538398 10208 538404 10220
rect 538456 10208 538462 10260
rect 193030 10140 193036 10192
rect 193088 10180 193094 10192
rect 534902 10180 534908 10192
rect 193088 10152 534908 10180
rect 193088 10140 193094 10152
rect 534902 10140 534908 10152
rect 534960 10140 534966 10192
rect 115566 10072 115572 10124
rect 115624 10112 115630 10124
rect 222746 10112 222752 10124
rect 115624 10084 222752 10112
rect 115624 10072 115630 10084
rect 222746 10072 222752 10084
rect 222804 10072 222810 10124
rect 114462 10004 114468 10056
rect 114520 10044 114526 10056
rect 219250 10044 219256 10056
rect 114520 10016 219256 10044
rect 114520 10004 114526 10016
rect 219250 10004 219256 10016
rect 219308 10004 219314 10056
rect 112806 9936 112812 9988
rect 112864 9976 112870 9988
rect 215662 9976 215668 9988
rect 112864 9948 215668 9976
rect 112864 9936 112870 9948
rect 215662 9936 215668 9948
rect 215720 9936 215726 9988
rect 112990 9868 112996 9920
rect 113048 9908 113054 9920
rect 212166 9908 212172 9920
rect 113048 9880 212172 9908
rect 113048 9868 113054 9880
rect 212166 9868 212172 9880
rect 212224 9868 212230 9920
rect 111426 9800 111432 9852
rect 111484 9840 111490 9852
rect 208578 9840 208584 9852
rect 111484 9812 208584 9840
rect 111484 9800 111490 9812
rect 208578 9800 208584 9812
rect 208636 9800 208642 9852
rect 111610 9732 111616 9784
rect 111668 9772 111674 9784
rect 205082 9772 205088 9784
rect 111668 9744 205088 9772
rect 111668 9732 111674 9744
rect 205082 9732 205088 9744
rect 205140 9732 205146 9784
rect 175090 9596 175096 9648
rect 175148 9636 175154 9648
rect 466270 9636 466276 9648
rect 175148 9608 466276 9636
rect 175148 9596 175154 9608
rect 466270 9596 466276 9608
rect 466328 9596 466334 9648
rect 176562 9528 176568 9580
rect 176620 9568 176626 9580
rect 469858 9568 469864 9580
rect 176620 9540 469864 9568
rect 176620 9528 176626 9540
rect 469858 9528 469864 9540
rect 469916 9528 469922 9580
rect 177758 9460 177764 9512
rect 177816 9500 177822 9512
rect 473446 9500 473452 9512
rect 177816 9472 473452 9500
rect 177816 9460 177822 9472
rect 473446 9460 473452 9472
rect 473504 9460 473510 9512
rect 177942 9392 177948 9444
rect 178000 9432 178006 9444
rect 475746 9432 475752 9444
rect 178000 9404 475752 9432
rect 178000 9392 178006 9404
rect 475746 9392 475752 9404
rect 475804 9392 475810 9444
rect 98914 9324 98920 9376
rect 98972 9364 98978 9376
rect 158898 9364 158904 9376
rect 98972 9336 158904 9364
rect 98972 9324 98978 9336
rect 158898 9324 158904 9336
rect 158956 9324 158962 9376
rect 177850 9324 177856 9376
rect 177908 9364 177914 9376
rect 476942 9364 476948 9376
rect 177908 9336 476948 9364
rect 177908 9324 177914 9336
rect 476942 9324 476948 9336
rect 477000 9324 477006 9376
rect 100478 9256 100484 9308
rect 100536 9296 100542 9308
rect 163682 9296 163688 9308
rect 100536 9268 163688 9296
rect 100536 9256 100542 9268
rect 163682 9256 163688 9268
rect 163740 9256 163746 9308
rect 179230 9256 179236 9308
rect 179288 9296 179294 9308
rect 481726 9296 481732 9308
rect 179288 9268 481732 9296
rect 179288 9256 179294 9268
rect 481726 9256 481732 9268
rect 481784 9256 481790 9308
rect 101858 9188 101864 9240
rect 101916 9228 101922 9240
rect 167178 9228 167184 9240
rect 101916 9200 167184 9228
rect 101916 9188 101922 9200
rect 167178 9188 167184 9200
rect 167236 9188 167242 9240
rect 180426 9188 180432 9240
rect 180484 9228 180490 9240
rect 485222 9228 485228 9240
rect 180484 9200 485228 9228
rect 180484 9188 180490 9200
rect 485222 9188 485228 9200
rect 485280 9188 485286 9240
rect 101766 9120 101772 9172
rect 101824 9160 101830 9172
rect 170766 9160 170772 9172
rect 101824 9132 170772 9160
rect 101824 9120 101830 9132
rect 170766 9120 170772 9132
rect 170824 9120 170830 9172
rect 180610 9120 180616 9172
rect 180668 9160 180674 9172
rect 488810 9160 488816 9172
rect 180668 9132 488816 9160
rect 180668 9120 180674 9132
rect 488810 9120 488816 9132
rect 488868 9120 488874 9172
rect 103330 9052 103336 9104
rect 103388 9092 103394 9104
rect 174262 9092 174268 9104
rect 103388 9064 174268 9092
rect 103388 9052 103394 9064
rect 174262 9052 174268 9064
rect 174320 9052 174326 9104
rect 181806 9052 181812 9104
rect 181864 9092 181870 9104
rect 492306 9092 492312 9104
rect 181864 9064 492312 9092
rect 181864 9052 181870 9064
rect 492306 9052 492312 9064
rect 492364 9052 492370 9104
rect 86218 8984 86224 9036
rect 86276 9024 86282 9036
rect 101030 9024 101036 9036
rect 86276 8996 101036 9024
rect 86276 8984 86282 8996
rect 101030 8984 101036 8996
rect 101088 8984 101094 9036
rect 104434 8984 104440 9036
rect 104492 9024 104498 9036
rect 177850 9024 177856 9036
rect 104492 8996 177856 9024
rect 104492 8984 104498 8996
rect 177850 8984 177856 8996
rect 177908 8984 177914 9036
rect 183094 8984 183100 9036
rect 183152 9024 183158 9036
rect 495894 9024 495900 9036
rect 183152 8996 495900 9024
rect 183152 8984 183158 8996
rect 495894 8984 495900 8996
rect 495952 8984 495958 9036
rect 86586 8916 86592 8968
rect 86644 8956 86650 8968
rect 104526 8956 104532 8968
rect 86644 8928 104532 8956
rect 86644 8916 86650 8928
rect 104526 8916 104532 8928
rect 104584 8916 104590 8968
rect 104618 8916 104624 8968
rect 104676 8956 104682 8968
rect 181438 8956 181444 8968
rect 104676 8928 181444 8956
rect 104676 8916 104682 8928
rect 181438 8916 181444 8928
rect 181496 8916 181502 8968
rect 183370 8916 183376 8968
rect 183428 8956 183434 8968
rect 499390 8956 499396 8968
rect 183428 8928 499396 8956
rect 183428 8916 183434 8928
rect 499390 8916 499396 8928
rect 499448 8916 499454 8968
rect 174998 8848 175004 8900
rect 175056 8888 175062 8900
rect 462774 8888 462780 8900
rect 175056 8860 462780 8888
rect 175056 8848 175062 8860
rect 462774 8848 462780 8860
rect 462832 8848 462838 8900
rect 173710 8780 173716 8832
rect 173768 8820 173774 8832
rect 459186 8820 459192 8832
rect 173768 8792 459192 8820
rect 173768 8780 173774 8792
rect 459186 8780 459192 8792
rect 459244 8780 459250 8832
rect 172238 8712 172244 8764
rect 172296 8752 172302 8764
rect 455690 8752 455696 8764
rect 172296 8724 455696 8752
rect 172296 8712 172302 8724
rect 455690 8712 455696 8724
rect 455748 8712 455754 8764
rect 172330 8644 172336 8696
rect 172388 8684 172394 8696
rect 452102 8684 452108 8696
rect 172388 8656 452108 8684
rect 172388 8644 172394 8656
rect 452102 8644 452108 8656
rect 452160 8644 452166 8696
rect 170950 8576 170956 8628
rect 171008 8616 171014 8628
rect 448606 8616 448612 8628
rect 171008 8588 448612 8616
rect 171008 8576 171014 8588
rect 448606 8576 448612 8588
rect 448664 8576 448670 8628
rect 169478 8508 169484 8560
rect 169536 8548 169542 8560
rect 445018 8548 445024 8560
rect 169536 8520 445024 8548
rect 169536 8508 169542 8520
rect 445018 8508 445024 8520
rect 445076 8508 445082 8560
rect 169570 8440 169576 8492
rect 169628 8480 169634 8492
rect 441522 8480 441528 8492
rect 169628 8452 441528 8480
rect 169628 8440 169634 8452
rect 441522 8440 441528 8452
rect 441580 8440 441586 8492
rect 168190 8372 168196 8424
rect 168248 8412 168254 8424
rect 437934 8412 437940 8424
rect 168248 8384 437940 8412
rect 168248 8372 168254 8384
rect 437934 8372 437940 8384
rect 437992 8372 437998 8424
rect 93118 8304 93124 8356
rect 93176 8344 93182 8356
rect 93946 8344 93952 8356
rect 93176 8316 93952 8344
rect 93176 8304 93182 8316
rect 93946 8304 93952 8316
rect 94004 8304 94010 8356
rect 168098 8304 168104 8356
rect 168156 8344 168162 8356
rect 434438 8344 434444 8356
rect 168156 8316 434444 8344
rect 168156 8304 168162 8316
rect 434438 8304 434444 8316
rect 434496 8304 434502 8356
rect 150250 8236 150256 8288
rect 150308 8276 150314 8288
rect 363506 8276 363512 8288
rect 150308 8248 363512 8276
rect 150308 8236 150314 8248
rect 363506 8236 363512 8248
rect 363564 8236 363570 8288
rect 151538 8168 151544 8220
rect 151596 8208 151602 8220
rect 367002 8208 367008 8220
rect 151596 8180 367008 8208
rect 151596 8168 151602 8180
rect 367002 8168 367008 8180
rect 367060 8168 367066 8220
rect 151446 8100 151452 8152
rect 151504 8140 151510 8152
rect 370590 8140 370596 8152
rect 151504 8112 370596 8140
rect 151504 8100 151510 8112
rect 370590 8100 370596 8112
rect 370648 8100 370654 8152
rect 152826 8032 152832 8084
rect 152884 8072 152890 8084
rect 374086 8072 374092 8084
rect 152884 8044 374092 8072
rect 152884 8032 152890 8044
rect 374086 8032 374092 8044
rect 374144 8032 374150 8084
rect 93578 7964 93584 8016
rect 93636 8004 93642 8016
rect 134150 8004 134156 8016
rect 93636 7976 134156 8004
rect 93636 7964 93642 7976
rect 134150 7964 134156 7976
rect 134208 7964 134214 8016
rect 152918 7964 152924 8016
rect 152976 8004 152982 8016
rect 377674 8004 377680 8016
rect 152976 7976 377680 8004
rect 152976 7964 152982 7976
rect 377674 7964 377680 7976
rect 377732 7964 377738 8016
rect 95050 7896 95056 7948
rect 95108 7936 95114 7948
rect 137646 7936 137652 7948
rect 95108 7908 137652 7936
rect 95108 7896 95114 7908
rect 137646 7896 137652 7908
rect 137704 7896 137710 7948
rect 154390 7896 154396 7948
rect 154448 7936 154454 7948
rect 381170 7936 381176 7948
rect 154448 7908 381176 7936
rect 154448 7896 154454 7908
rect 381170 7896 381176 7908
rect 381228 7896 381234 7948
rect 95142 7828 95148 7880
rect 95200 7868 95206 7880
rect 141234 7868 141240 7880
rect 95200 7840 141240 7868
rect 95200 7828 95206 7840
rect 141234 7828 141240 7840
rect 141292 7828 141298 7880
rect 155770 7828 155776 7880
rect 155828 7868 155834 7880
rect 384758 7868 384764 7880
rect 155828 7840 384764 7868
rect 155828 7828 155834 7840
rect 384758 7828 384764 7840
rect 384816 7828 384822 7880
rect 96338 7760 96344 7812
rect 96396 7800 96402 7812
rect 144730 7800 144736 7812
rect 96396 7772 144736 7800
rect 96396 7760 96402 7772
rect 144730 7760 144736 7772
rect 144788 7760 144794 7812
rect 155678 7760 155684 7812
rect 155736 7800 155742 7812
rect 388254 7800 388260 7812
rect 155736 7772 388260 7800
rect 155736 7760 155742 7772
rect 388254 7760 388260 7772
rect 388312 7760 388318 7812
rect 96246 7692 96252 7744
rect 96304 7732 96310 7744
rect 148226 7732 148232 7744
rect 96304 7704 148232 7732
rect 96304 7692 96310 7704
rect 148226 7692 148232 7704
rect 148284 7692 148290 7744
rect 157150 7692 157156 7744
rect 157208 7732 157214 7744
rect 391842 7732 391848 7744
rect 157208 7704 391848 7732
rect 157208 7692 157214 7704
rect 391842 7692 391848 7704
rect 391900 7692 391906 7744
rect 97902 7624 97908 7676
rect 97960 7664 97966 7676
rect 151814 7664 151820 7676
rect 97960 7636 151820 7664
rect 97960 7624 97966 7636
rect 151814 7624 151820 7636
rect 151872 7624 151878 7676
rect 158530 7624 158536 7676
rect 158588 7664 158594 7676
rect 395338 7664 395344 7676
rect 158588 7636 395344 7664
rect 158588 7624 158594 7636
rect 395338 7624 395344 7636
rect 395396 7624 395402 7676
rect 99006 7556 99012 7608
rect 99064 7596 99070 7608
rect 155402 7596 155408 7608
rect 99064 7568 155408 7596
rect 99064 7556 99070 7568
rect 155402 7556 155408 7568
rect 155460 7556 155466 7608
rect 158438 7556 158444 7608
rect 158496 7596 158502 7608
rect 398926 7596 398932 7608
rect 158496 7568 398932 7596
rect 158496 7556 158502 7568
rect 398926 7556 398932 7568
rect 398984 7556 398990 7608
rect 148870 7488 148876 7540
rect 148928 7528 148934 7540
rect 359918 7528 359924 7540
rect 148928 7500 359924 7528
rect 148928 7488 148934 7500
rect 359918 7488 359924 7500
rect 359976 7488 359982 7540
rect 148778 7420 148784 7472
rect 148836 7460 148842 7472
rect 356330 7460 356336 7472
rect 148836 7432 356336 7460
rect 148836 7420 148842 7432
rect 356330 7420 356336 7432
rect 356388 7420 356394 7472
rect 147306 7352 147312 7404
rect 147364 7392 147370 7404
rect 352834 7392 352840 7404
rect 147364 7364 352840 7392
rect 147364 7352 147370 7364
rect 352834 7352 352840 7364
rect 352892 7352 352898 7404
rect 146110 7284 146116 7336
rect 146168 7324 146174 7336
rect 345750 7324 345756 7336
rect 146168 7296 345756 7324
rect 146168 7284 146174 7296
rect 345750 7284 345756 7296
rect 345808 7284 345814 7336
rect 144822 7216 144828 7268
rect 144880 7256 144886 7268
rect 342162 7256 342168 7268
rect 144880 7228 342168 7256
rect 144880 7216 144886 7228
rect 342162 7216 342168 7228
rect 342220 7216 342226 7268
rect 143350 7148 143356 7200
rect 143408 7188 143414 7200
rect 338666 7188 338672 7200
rect 143408 7160 338672 7188
rect 143408 7148 143414 7160
rect 338666 7148 338672 7160
rect 338724 7148 338730 7200
rect 143442 7080 143448 7132
rect 143500 7120 143506 7132
rect 335078 7120 335084 7132
rect 143500 7092 335084 7120
rect 143500 7080 143506 7092
rect 335078 7080 335084 7092
rect 335136 7080 335142 7132
rect 141786 7012 141792 7064
rect 141844 7052 141850 7064
rect 331582 7052 331588 7064
rect 141844 7024 331588 7052
rect 141844 7012 141850 7024
rect 331582 7012 331588 7024
rect 331640 7012 331646 7064
rect 3418 6808 3424 6860
rect 3476 6848 3482 6860
rect 22738 6848 22744 6860
rect 3476 6820 22744 6848
rect 3476 6808 3482 6820
rect 22738 6808 22744 6820
rect 22796 6808 22802 6860
rect 125502 6808 125508 6860
rect 125560 6848 125566 6860
rect 264146 6848 264152 6860
rect 125560 6820 264152 6848
rect 125560 6808 125566 6820
rect 264146 6808 264152 6820
rect 264204 6808 264210 6860
rect 126882 6740 126888 6792
rect 126940 6780 126946 6792
rect 267734 6780 267740 6792
rect 126940 6752 267740 6780
rect 126940 6740 126946 6752
rect 267734 6740 267740 6752
rect 267792 6740 267798 6792
rect 126790 6672 126796 6724
rect 126848 6712 126854 6724
rect 271230 6712 271236 6724
rect 126848 6684 271236 6712
rect 126848 6672 126854 6684
rect 271230 6672 271236 6684
rect 271288 6672 271294 6724
rect 128170 6604 128176 6656
rect 128228 6644 128234 6656
rect 274818 6644 274824 6656
rect 128228 6616 274824 6644
rect 128228 6604 128234 6616
rect 274818 6604 274824 6616
rect 274876 6604 274882 6656
rect 129642 6536 129648 6588
rect 129700 6576 129706 6588
rect 278314 6576 278320 6588
rect 129700 6548 278320 6576
rect 129700 6536 129706 6548
rect 278314 6536 278320 6548
rect 278372 6536 278378 6588
rect 129550 6468 129556 6520
rect 129608 6508 129614 6520
rect 281902 6508 281908 6520
rect 129608 6480 281908 6508
rect 129608 6468 129614 6480
rect 281902 6468 281908 6480
rect 281960 6468 281966 6520
rect 130930 6400 130936 6452
rect 130988 6440 130994 6452
rect 285398 6440 285404 6452
rect 130988 6412 285404 6440
rect 130988 6400 130994 6412
rect 285398 6400 285404 6412
rect 285456 6400 285462 6452
rect 132402 6332 132408 6384
rect 132460 6372 132466 6384
rect 288986 6372 288992 6384
rect 132460 6344 288992 6372
rect 132460 6332 132466 6344
rect 288986 6332 288992 6344
rect 289044 6332 289050 6384
rect 132310 6264 132316 6316
rect 132368 6304 132374 6316
rect 292574 6304 292580 6316
rect 132368 6276 292580 6304
rect 132368 6264 132374 6276
rect 292574 6264 292580 6276
rect 292632 6264 292638 6316
rect 105538 6196 105544 6248
rect 105596 6236 105602 6248
rect 128170 6236 128176 6248
rect 105596 6208 128176 6236
rect 105596 6196 105602 6208
rect 128170 6196 128176 6208
rect 128228 6196 128234 6248
rect 133506 6196 133512 6248
rect 133564 6236 133570 6248
rect 296070 6236 296076 6248
rect 133564 6208 296076 6236
rect 133564 6196 133570 6208
rect 296070 6196 296076 6208
rect 296128 6196 296134 6248
rect 92198 6128 92204 6180
rect 92256 6168 92262 6180
rect 130562 6168 130568 6180
rect 92256 6140 130568 6168
rect 92256 6128 92262 6140
rect 130562 6128 130568 6140
rect 130620 6128 130626 6180
rect 151630 6128 151636 6180
rect 151688 6168 151694 6180
rect 369394 6168 369400 6180
rect 151688 6140 369400 6168
rect 151688 6128 151694 6140
rect 369394 6128 369400 6140
rect 369452 6128 369458 6180
rect 125410 6060 125416 6112
rect 125468 6100 125474 6112
rect 260650 6100 260656 6112
rect 125468 6072 260656 6100
rect 125468 6060 125474 6072
rect 260650 6060 260656 6072
rect 260708 6060 260714 6112
rect 124122 5992 124128 6044
rect 124180 6032 124186 6044
rect 257062 6032 257068 6044
rect 124180 6004 257068 6032
rect 124180 5992 124186 6004
rect 257062 5992 257068 6004
rect 257120 5992 257126 6044
rect 122650 5924 122656 5976
rect 122708 5964 122714 5976
rect 253474 5964 253480 5976
rect 122708 5936 253480 5964
rect 122708 5924 122714 5936
rect 253474 5924 253480 5936
rect 253532 5924 253538 5976
rect 122374 5856 122380 5908
rect 122432 5896 122438 5908
rect 249978 5896 249984 5908
rect 122432 5868 249984 5896
rect 122432 5856 122438 5868
rect 249978 5856 249984 5868
rect 250036 5856 250042 5908
rect 121362 5788 121368 5840
rect 121420 5828 121426 5840
rect 246390 5828 246396 5840
rect 121420 5800 246396 5828
rect 121420 5788 121426 5800
rect 246390 5788 246396 5800
rect 246448 5788 246454 5840
rect 119614 5720 119620 5772
rect 119672 5760 119678 5772
rect 242986 5760 242992 5772
rect 119672 5732 242992 5760
rect 119672 5720 119678 5732
rect 242986 5720 242992 5732
rect 243044 5720 243050 5772
rect 119890 5652 119896 5704
rect 119948 5692 119954 5704
rect 239306 5692 239312 5704
rect 119948 5664 239312 5692
rect 119948 5652 119954 5664
rect 239306 5652 239312 5664
rect 239364 5652 239370 5704
rect 118602 5584 118608 5636
rect 118660 5624 118666 5636
rect 235810 5624 235816 5636
rect 118660 5596 235816 5624
rect 118660 5584 118666 5596
rect 235810 5584 235816 5596
rect 235868 5584 235874 5636
rect 116946 5516 116952 5568
rect 117004 5556 117010 5568
rect 232222 5556 232228 5568
rect 117004 5528 232228 5556
rect 117004 5516 117010 5528
rect 232222 5516 232228 5528
rect 232280 5516 232286 5568
rect 276014 5516 276020 5568
rect 276072 5556 276078 5568
rect 277118 5556 277124 5568
rect 276072 5528 277124 5556
rect 276072 5516 276078 5528
rect 277118 5516 277124 5528
rect 277176 5516 277182 5568
rect 299566 5516 299572 5568
rect 299624 5556 299630 5568
rect 300762 5556 300768 5568
rect 299624 5528 300768 5556
rect 299624 5516 299630 5528
rect 300762 5516 300768 5528
rect 300820 5516 300826 5568
rect 101950 5448 101956 5500
rect 102008 5488 102014 5500
rect 166074 5488 166080 5500
rect 102008 5460 166080 5488
rect 102008 5448 102014 5460
rect 166074 5448 166080 5460
rect 166132 5448 166138 5500
rect 191466 5448 191472 5500
rect 191524 5488 191530 5500
rect 533706 5488 533712 5500
rect 191524 5460 533712 5488
rect 191524 5448 191530 5460
rect 533706 5448 533712 5460
rect 533764 5448 533770 5500
rect 102042 5380 102048 5432
rect 102100 5420 102106 5432
rect 169570 5420 169576 5432
rect 102100 5392 169576 5420
rect 102100 5380 102106 5392
rect 169570 5380 169576 5392
rect 169628 5380 169634 5432
rect 192754 5380 192760 5432
rect 192812 5420 192818 5432
rect 537202 5420 537208 5432
rect 192812 5392 537208 5420
rect 192812 5380 192818 5392
rect 537202 5380 537208 5392
rect 537260 5380 537266 5432
rect 103422 5312 103428 5364
rect 103480 5352 103486 5364
rect 173158 5352 173164 5364
rect 103480 5324 173164 5352
rect 103480 5312 103486 5324
rect 173158 5312 173164 5324
rect 173216 5312 173222 5364
rect 194410 5312 194416 5364
rect 194468 5352 194474 5364
rect 540790 5352 540796 5364
rect 194468 5324 540796 5352
rect 194468 5312 194474 5324
rect 540790 5312 540796 5324
rect 540848 5312 540854 5364
rect 104802 5244 104808 5296
rect 104860 5284 104866 5296
rect 176654 5284 176660 5296
rect 104860 5256 176660 5284
rect 104860 5244 104866 5256
rect 176654 5244 176660 5256
rect 176712 5244 176718 5296
rect 196894 5244 196900 5296
rect 196952 5284 196958 5296
rect 204898 5284 204904 5296
rect 196952 5256 204904 5284
rect 196952 5244 196958 5256
rect 204898 5244 204904 5256
rect 204956 5244 204962 5296
rect 204990 5244 204996 5296
rect 205048 5284 205054 5296
rect 544286 5284 544292 5296
rect 205048 5256 544292 5284
rect 205048 5244 205054 5256
rect 544286 5244 544292 5256
rect 544344 5244 544350 5296
rect 104710 5176 104716 5228
rect 104768 5216 104774 5228
rect 180242 5216 180248 5228
rect 104768 5188 180248 5216
rect 104768 5176 104774 5188
rect 180242 5176 180248 5188
rect 180300 5176 180306 5228
rect 195882 5176 195888 5228
rect 195940 5216 195946 5228
rect 547966 5216 547972 5228
rect 195940 5188 547972 5216
rect 195940 5176 195946 5188
rect 547966 5176 547972 5188
rect 548024 5176 548030 5228
rect 106182 5108 106188 5160
rect 106240 5148 106246 5160
rect 183738 5148 183744 5160
rect 106240 5120 183744 5148
rect 106240 5108 106246 5120
rect 183738 5108 183744 5120
rect 183796 5108 183802 5160
rect 187234 5108 187240 5160
rect 187292 5148 187298 5160
rect 195330 5148 195336 5160
rect 187292 5120 195336 5148
rect 187292 5108 187298 5120
rect 195330 5108 195336 5120
rect 195388 5108 195394 5160
rect 197170 5108 197176 5160
rect 197228 5148 197234 5160
rect 551462 5148 551468 5160
rect 197228 5120 551468 5148
rect 197228 5108 197234 5120
rect 551462 5108 551468 5120
rect 551520 5108 551526 5160
rect 106090 5040 106096 5092
rect 106148 5080 106154 5092
rect 187326 5080 187332 5092
rect 106148 5052 187332 5080
rect 106148 5040 106154 5052
rect 187326 5040 187332 5052
rect 187384 5040 187390 5092
rect 200298 5080 200304 5092
rect 194336 5052 200304 5080
rect 107470 4972 107476 5024
rect 107528 5012 107534 5024
rect 189718 5012 189724 5024
rect 107528 4984 189724 5012
rect 107528 4972 107534 4984
rect 189718 4972 189724 4984
rect 189776 4972 189782 5024
rect 194336 5012 194364 5052
rect 200298 5040 200304 5052
rect 200356 5040 200362 5092
rect 201310 5040 201316 5092
rect 201368 5080 201374 5092
rect 204806 5080 204812 5092
rect 201368 5052 204812 5080
rect 201368 5040 201374 5052
rect 204806 5040 204812 5052
rect 204864 5040 204870 5092
rect 204898 5040 204904 5092
rect 204956 5080 204962 5092
rect 554958 5080 554964 5092
rect 204956 5052 554964 5080
rect 204956 5040 204962 5052
rect 554958 5040 554964 5052
rect 555016 5040 555022 5092
rect 193968 4984 194364 5012
rect 107562 4904 107568 4956
rect 107620 4944 107626 4956
rect 193306 4944 193312 4956
rect 107620 4916 193312 4944
rect 107620 4904 107626 4916
rect 193306 4904 193312 4916
rect 193364 4904 193370 4956
rect 108942 4836 108948 4888
rect 109000 4876 109006 4888
rect 193858 4876 193864 4888
rect 109000 4848 193864 4876
rect 109000 4836 109006 4848
rect 193858 4836 193864 4848
rect 193916 4836 193922 4888
rect 110322 4768 110328 4820
rect 110380 4808 110386 4820
rect 193968 4808 193996 4984
rect 198550 4972 198556 5024
rect 198608 5012 198614 5024
rect 558546 5012 558552 5024
rect 198608 4984 558552 5012
rect 198608 4972 198614 4984
rect 558546 4972 558552 4984
rect 558604 4972 558610 5024
rect 194134 4904 194140 4956
rect 194192 4944 194198 4956
rect 194192 4916 197216 4944
rect 194192 4904 194198 4916
rect 194042 4836 194048 4888
rect 194100 4876 194106 4888
rect 196802 4876 196808 4888
rect 194100 4848 196808 4876
rect 194100 4836 194106 4848
rect 196802 4836 196808 4848
rect 196860 4836 196866 4888
rect 197188 4876 197216 4916
rect 198274 4904 198280 4956
rect 198332 4944 198338 4956
rect 562042 4944 562048 4956
rect 198332 4916 562048 4944
rect 198332 4904 198338 4916
rect 562042 4904 562048 4916
rect 562100 4904 562106 4956
rect 204714 4876 204720 4888
rect 197188 4848 204720 4876
rect 204714 4836 204720 4848
rect 204772 4836 204778 4888
rect 204990 4836 204996 4888
rect 205048 4876 205054 4888
rect 569126 4876 569132 4888
rect 205048 4848 569132 4876
rect 205048 4836 205054 4848
rect 569126 4836 569132 4848
rect 569184 4836 569190 4888
rect 110380 4780 193996 4808
rect 110380 4768 110386 4780
rect 195054 4768 195060 4820
rect 195112 4808 195118 4820
rect 203886 4808 203892 4820
rect 195112 4780 203892 4808
rect 195112 4768 195118 4780
rect 203886 4768 203892 4780
rect 203944 4768 203950 4820
rect 204162 4768 204168 4820
rect 204220 4808 204226 4820
rect 580994 4808 581000 4820
rect 204220 4780 581000 4808
rect 204220 4768 204226 4780
rect 580994 4768 581000 4780
rect 581052 4768 581058 4820
rect 100570 4700 100576 4752
rect 100628 4740 100634 4752
rect 162486 4740 162492 4752
rect 100628 4712 162492 4740
rect 100628 4700 100634 4712
rect 162486 4700 162492 4712
rect 162544 4700 162550 4752
rect 191650 4700 191656 4752
rect 191708 4740 191714 4752
rect 530118 4740 530124 4752
rect 191708 4712 530124 4740
rect 191708 4700 191714 4712
rect 530118 4700 530124 4712
rect 530176 4700 530182 4752
rect 99190 4632 99196 4684
rect 99248 4672 99254 4684
rect 157794 4672 157800 4684
rect 99248 4644 157800 4672
rect 99248 4632 99254 4644
rect 157794 4632 157800 4644
rect 157852 4632 157858 4684
rect 190086 4632 190092 4684
rect 190144 4672 190150 4684
rect 526622 4672 526628 4684
rect 190144 4644 526628 4672
rect 190144 4632 190150 4644
rect 526622 4632 526628 4644
rect 526680 4632 526686 4684
rect 96522 4564 96528 4616
rect 96580 4604 96586 4616
rect 147122 4604 147128 4616
rect 96580 4576 147128 4604
rect 96580 4564 96586 4576
rect 147122 4564 147128 4576
rect 147180 4564 147186 4616
rect 147214 4564 147220 4616
rect 147272 4604 147278 4616
rect 195054 4604 195060 4616
rect 147272 4576 195060 4604
rect 147272 4564 147278 4576
rect 195054 4564 195060 4576
rect 195112 4564 195118 4616
rect 195146 4564 195152 4616
rect 195204 4604 195210 4616
rect 523034 4604 523040 4616
rect 195204 4576 523040 4604
rect 195204 4564 195210 4576
rect 523034 4564 523040 4576
rect 523092 4564 523098 4616
rect 99098 4496 99104 4548
rect 99156 4536 99162 4548
rect 154206 4536 154212 4548
rect 99156 4508 154212 4536
rect 99156 4496 99162 4508
rect 154206 4496 154212 4508
rect 154264 4496 154270 4548
rect 188890 4496 188896 4548
rect 188948 4536 188954 4548
rect 519538 4536 519544 4548
rect 188948 4508 519544 4536
rect 188948 4496 188954 4508
rect 519538 4496 519544 4508
rect 519596 4496 519602 4548
rect 96430 4428 96436 4480
rect 96488 4468 96494 4480
rect 143534 4468 143540 4480
rect 96488 4440 143540 4468
rect 96488 4428 96494 4440
rect 143534 4428 143540 4440
rect 143592 4428 143598 4480
rect 146938 4428 146944 4480
rect 146996 4468 147002 4480
rect 182542 4468 182548 4480
rect 146996 4440 182548 4468
rect 146996 4428 147002 4440
rect 182542 4428 182548 4440
rect 182600 4428 182606 4480
rect 188614 4428 188620 4480
rect 188672 4468 188678 4480
rect 195146 4468 195152 4480
rect 188672 4440 195152 4468
rect 188672 4428 188678 4440
rect 195146 4428 195152 4440
rect 195204 4428 195210 4480
rect 515950 4468 515956 4480
rect 195256 4440 515956 4468
rect 93762 4360 93768 4412
rect 93820 4400 93826 4412
rect 136450 4400 136456 4412
rect 93820 4372 136456 4400
rect 93820 4360 93826 4372
rect 136450 4360 136456 4372
rect 136508 4360 136514 4412
rect 142798 4360 142804 4412
rect 142856 4400 142862 4412
rect 186130 4400 186136 4412
rect 142856 4372 186136 4400
rect 142856 4360 142862 4372
rect 186130 4360 186136 4372
rect 186188 4360 186194 4412
rect 187510 4360 187516 4412
rect 187568 4400 187574 4412
rect 195256 4400 195284 4440
rect 515950 4428 515956 4440
rect 516008 4428 516014 4480
rect 187568 4372 195284 4400
rect 187568 4360 187574 4372
rect 195330 4360 195336 4412
rect 195388 4400 195394 4412
rect 512454 4400 512460 4412
rect 195388 4372 512460 4400
rect 195388 4360 195394 4372
rect 512454 4360 512460 4372
rect 512512 4360 512518 4412
rect 93670 4292 93676 4344
rect 93728 4332 93734 4344
rect 132954 4332 132960 4344
rect 93728 4304 132960 4332
rect 93728 4292 93734 4304
rect 132954 4292 132960 4304
rect 133012 4292 133018 4344
rect 173802 4292 173808 4344
rect 173860 4332 173866 4344
rect 458082 4332 458088 4344
rect 173860 4304 458088 4332
rect 173860 4292 173866 4304
rect 458082 4292 458088 4304
rect 458140 4292 458146 4344
rect 92290 4224 92296 4276
rect 92348 4264 92354 4276
rect 126974 4264 126980 4276
rect 92348 4236 126980 4264
rect 92348 4224 92354 4236
rect 126974 4224 126980 4236
rect 127032 4224 127038 4276
rect 172146 4224 172152 4276
rect 172204 4264 172210 4276
rect 450906 4264 450912 4276
rect 172204 4236 450912 4264
rect 172204 4224 172210 4236
rect 450906 4224 450912 4236
rect 450964 4224 450970 4276
rect 99282 4156 99288 4208
rect 99340 4196 99346 4208
rect 99340 4168 103468 4196
rect 99340 4156 99346 4168
rect 21818 4088 21824 4140
rect 21876 4128 21882 4140
rect 21876 4100 22094 4128
rect 21876 4088 21882 4100
rect 22066 4060 22094 4100
rect 24210 4088 24216 4140
rect 24268 4128 24274 4140
rect 24762 4128 24768 4140
rect 24268 4100 24768 4128
rect 24268 4088 24274 4100
rect 24762 4088 24768 4100
rect 24820 4088 24826 4140
rect 27706 4088 27712 4140
rect 27764 4128 27770 4140
rect 28902 4128 28908 4140
rect 27764 4100 28908 4128
rect 27764 4088 27770 4100
rect 28902 4088 28908 4100
rect 28960 4088 28966 4140
rect 28994 4088 29000 4140
rect 29052 4128 29058 4140
rect 65150 4128 65156 4140
rect 29052 4100 65156 4128
rect 29052 4088 29058 4100
rect 65150 4088 65156 4100
rect 65208 4088 65214 4140
rect 84010 4088 84016 4140
rect 84068 4128 84074 4140
rect 96246 4128 96252 4140
rect 84068 4100 96252 4128
rect 84068 4088 84074 4100
rect 96246 4088 96252 4100
rect 96304 4088 96310 4140
rect 97258 4088 97264 4140
rect 97316 4128 97322 4140
rect 103330 4128 103336 4140
rect 97316 4100 103336 4128
rect 97316 4088 97322 4100
rect 103330 4088 103336 4100
rect 103388 4088 103394 4140
rect 103440 4128 103468 4168
rect 171042 4156 171048 4208
rect 171100 4196 171106 4208
rect 447410 4196 447416 4208
rect 171100 4168 447416 4196
rect 171100 4156 171106 4168
rect 447410 4156 447416 4168
rect 447468 4156 447474 4208
rect 156598 4128 156604 4140
rect 103440 4100 156604 4128
rect 156598 4088 156604 4100
rect 156656 4088 156662 4140
rect 220170 4088 220176 4140
rect 220228 4128 220234 4140
rect 390646 4128 390652 4140
rect 220228 4100 390652 4128
rect 220228 4088 220234 4100
rect 390646 4088 390652 4100
rect 390704 4088 390710 4140
rect 436738 4088 436744 4140
rect 436796 4128 436802 4140
rect 442626 4128 442632 4140
rect 436796 4100 442632 4128
rect 436796 4088 436802 4100
rect 442626 4088 442632 4100
rect 442684 4088 442690 4140
rect 479518 4088 479524 4140
rect 479576 4128 479582 4140
rect 480530 4128 480536 4140
rect 479576 4100 480536 4128
rect 479576 4088 479582 4100
rect 480530 4088 480536 4100
rect 480588 4088 480594 4140
rect 65058 4060 65064 4072
rect 22066 4032 65064 4060
rect 65058 4020 65064 4032
rect 65116 4020 65122 4072
rect 85390 4020 85396 4072
rect 85448 4060 85454 4072
rect 94406 4060 94412 4072
rect 85448 4032 94412 4060
rect 85448 4020 85454 4032
rect 94406 4020 94412 4032
rect 94464 4020 94470 4072
rect 94498 4020 94504 4072
rect 94556 4060 94562 4072
rect 99834 4060 99840 4072
rect 94556 4032 99840 4060
rect 94556 4020 94562 4032
rect 99834 4020 99840 4032
rect 99892 4020 99898 4072
rect 100662 4020 100668 4072
rect 100720 4060 100726 4072
rect 160094 4060 160100 4072
rect 100720 4032 160100 4060
rect 100720 4020 100726 4032
rect 160094 4020 160100 4032
rect 160152 4020 160158 4072
rect 215938 4020 215944 4072
rect 215996 4060 216002 4072
rect 404814 4060 404820 4072
rect 215996 4032 404820 4060
rect 215996 4020 216002 4032
rect 404814 4020 404820 4032
rect 404872 4020 404878 4072
rect 26878 3952 26884 4004
rect 26936 3992 26942 4004
rect 63678 3992 63684 4004
rect 26936 3964 63684 3992
rect 26936 3952 26942 3964
rect 63678 3952 63684 3964
rect 63736 3952 63742 4004
rect 88242 3952 88248 4004
rect 88300 3992 88306 4004
rect 114002 3992 114008 4004
rect 88300 3964 114008 3992
rect 88300 3952 88306 3964
rect 114002 3952 114008 3964
rect 114060 3952 114066 4004
rect 146202 3952 146208 4004
rect 146260 3992 146266 4004
rect 348050 3992 348056 4004
rect 146260 3964 348056 3992
rect 146260 3952 146266 3964
rect 348050 3952 348056 3964
rect 348108 3952 348114 4004
rect 475378 3952 475384 4004
rect 475436 3992 475442 4004
rect 510062 3992 510068 4004
rect 475436 3964 510068 3992
rect 475436 3952 475442 3964
rect 510062 3952 510068 3964
rect 510120 3952 510126 4004
rect 18230 3884 18236 3936
rect 18288 3924 18294 3936
rect 63494 3924 63500 3936
rect 18288 3896 63500 3924
rect 18288 3884 18294 3896
rect 63494 3884 63500 3896
rect 63552 3884 63558 3936
rect 89622 3884 89628 3936
rect 89680 3924 89686 3936
rect 115198 3924 115204 3936
rect 89680 3896 115204 3924
rect 89680 3884 89686 3896
rect 115198 3884 115204 3896
rect 115256 3884 115262 3936
rect 147490 3884 147496 3936
rect 147548 3924 147554 3936
rect 351638 3924 351644 3936
rect 147548 3896 351644 3924
rect 147548 3884 147554 3896
rect 351638 3884 351644 3896
rect 351696 3884 351702 3936
rect 472618 3884 472624 3936
rect 472676 3924 472682 3936
rect 506474 3924 506480 3936
rect 472676 3896 506480 3924
rect 472676 3884 472682 3896
rect 506474 3884 506480 3896
rect 506532 3884 506538 3936
rect 20622 3816 20628 3868
rect 20680 3856 20686 3868
rect 64966 3856 64972 3868
rect 20680 3828 64972 3856
rect 20680 3816 20686 3828
rect 64966 3816 64972 3828
rect 65024 3816 65030 3868
rect 89530 3816 89536 3868
rect 89588 3856 89594 3868
rect 118786 3856 118792 3868
rect 89588 3828 118792 3856
rect 89588 3816 89594 3828
rect 118786 3816 118792 3828
rect 118844 3816 118850 3868
rect 147398 3816 147404 3868
rect 147456 3856 147462 3868
rect 354030 3856 354036 3868
rect 147456 3828 354036 3856
rect 147456 3816 147462 3828
rect 354030 3816 354036 3828
rect 354088 3816 354094 3868
rect 468478 3816 468484 3868
rect 468536 3856 468542 3868
rect 505370 3856 505376 3868
rect 468536 3828 505376 3856
rect 468536 3816 468542 3828
rect 505370 3816 505376 3828
rect 505428 3816 505434 3868
rect 15930 3748 15936 3800
rect 15988 3788 15994 3800
rect 55674 3788 55680 3800
rect 15988 3760 55680 3788
rect 15988 3748 15994 3760
rect 55674 3748 55680 3760
rect 55732 3748 55738 3800
rect 55766 3748 55772 3800
rect 55824 3788 55830 3800
rect 61010 3788 61016 3800
rect 55824 3760 61016 3788
rect 55824 3748 55830 3760
rect 61010 3748 61016 3760
rect 61068 3748 61074 3800
rect 89346 3748 89352 3800
rect 89404 3788 89410 3800
rect 116394 3788 116400 3800
rect 89404 3760 116400 3788
rect 89404 3748 89410 3760
rect 116394 3748 116400 3760
rect 116452 3748 116458 3800
rect 147582 3748 147588 3800
rect 147640 3788 147646 3800
rect 355226 3788 355232 3800
rect 147640 3760 355232 3788
rect 147640 3748 147646 3760
rect 355226 3748 355232 3760
rect 355284 3748 355290 3800
rect 421558 3748 421564 3800
rect 421616 3788 421622 3800
rect 423674 3788 423680 3800
rect 421616 3760 423680 3788
rect 421616 3748 421622 3760
rect 423674 3748 423680 3760
rect 423732 3748 423738 3800
rect 432598 3748 432604 3800
rect 432656 3788 432662 3800
rect 460382 3788 460388 3800
rect 432656 3760 460388 3788
rect 432656 3748 432662 3760
rect 460382 3748 460388 3760
rect 460440 3748 460446 3800
rect 461670 3748 461676 3800
rect 461728 3788 461734 3800
rect 498194 3788 498200 3800
rect 461728 3760 498200 3788
rect 461728 3748 461734 3760
rect 498194 3748 498200 3760
rect 498252 3748 498258 3800
rect 12250 3680 12256 3732
rect 12308 3720 12314 3732
rect 59998 3720 60004 3732
rect 12308 3692 60004 3720
rect 12308 3680 12314 3692
rect 59998 3680 60004 3692
rect 60056 3680 60062 3732
rect 60826 3680 60832 3732
rect 60884 3720 60890 3732
rect 74902 3720 74908 3732
rect 60884 3692 74908 3720
rect 60884 3680 60890 3692
rect 74902 3680 74908 3692
rect 74960 3680 74966 3732
rect 81158 3680 81164 3732
rect 81216 3720 81222 3732
rect 85666 3720 85672 3732
rect 81216 3692 85672 3720
rect 81216 3680 81222 3692
rect 85666 3680 85672 3692
rect 85724 3680 85730 3732
rect 89438 3680 89444 3732
rect 89496 3720 89502 3732
rect 119890 3720 119896 3732
rect 89496 3692 119896 3720
rect 89496 3680 89502 3692
rect 119890 3680 119896 3692
rect 119948 3680 119954 3732
rect 120718 3680 120724 3732
rect 120776 3720 120782 3732
rect 129366 3720 129372 3732
rect 120776 3692 129372 3720
rect 120776 3680 120782 3692
rect 129366 3680 129372 3692
rect 129424 3680 129430 3732
rect 148594 3680 148600 3732
rect 148652 3720 148658 3732
rect 358722 3720 358728 3732
rect 148652 3692 358728 3720
rect 148652 3680 148658 3692
rect 358722 3680 358728 3692
rect 358780 3680 358786 3732
rect 447778 3680 447784 3732
rect 447836 3720 447842 3732
rect 447836 3692 450032 3720
rect 447836 3680 447842 3692
rect 7650 3612 7656 3664
rect 7708 3652 7714 3664
rect 55766 3652 55772 3664
rect 7708 3624 55772 3652
rect 7708 3612 7714 3624
rect 55766 3612 55772 3624
rect 55824 3612 55830 3664
rect 60734 3652 60740 3664
rect 55876 3624 60740 3652
rect 5258 3544 5264 3596
rect 5316 3584 5322 3596
rect 55876 3584 55904 3624
rect 60734 3612 60740 3624
rect 60792 3612 60798 3664
rect 74810 3652 74816 3664
rect 64846 3624 74816 3652
rect 59446 3584 59452 3596
rect 5316 3556 55904 3584
rect 55968 3556 59452 3584
rect 5316 3544 5322 3556
rect 2866 3476 2872 3528
rect 2924 3516 2930 3528
rect 55968 3516 55996 3556
rect 59446 3544 59452 3556
rect 59504 3544 59510 3596
rect 59722 3544 59728 3596
rect 59780 3584 59786 3596
rect 63862 3584 63868 3596
rect 59780 3556 63868 3584
rect 59780 3544 59786 3556
rect 63862 3544 63868 3556
rect 63920 3544 63926 3596
rect 64322 3544 64328 3596
rect 64380 3584 64386 3596
rect 64846 3584 64874 3624
rect 74810 3612 74816 3624
rect 74868 3612 74874 3664
rect 91002 3612 91008 3664
rect 91060 3652 91066 3664
rect 122282 3652 122288 3664
rect 91060 3624 122288 3652
rect 91060 3612 91066 3624
rect 122282 3612 122288 3624
rect 122340 3612 122346 3664
rect 150342 3612 150348 3664
rect 150400 3652 150406 3664
rect 365806 3652 365812 3664
rect 150400 3624 365812 3652
rect 150400 3612 150406 3624
rect 365806 3612 365812 3624
rect 365864 3612 365870 3664
rect 443638 3612 443644 3664
rect 443696 3652 443702 3664
rect 443696 3624 449940 3652
rect 443696 3612 443702 3624
rect 64380 3556 64874 3584
rect 64380 3544 64386 3556
rect 69106 3544 69112 3596
rect 69164 3584 69170 3596
rect 70210 3584 70216 3596
rect 69164 3556 70216 3584
rect 69164 3544 69170 3556
rect 70210 3544 70216 3556
rect 70268 3544 70274 3596
rect 73798 3544 73804 3596
rect 73856 3584 73862 3596
rect 76558 3584 76564 3596
rect 73856 3556 76564 3584
rect 73856 3544 73862 3556
rect 76558 3544 76564 3556
rect 76616 3544 76622 3596
rect 77386 3544 77392 3596
rect 77444 3584 77450 3596
rect 78766 3584 78772 3596
rect 77444 3556 78772 3584
rect 77444 3544 77450 3556
rect 78766 3544 78772 3556
rect 78824 3544 78830 3596
rect 82722 3544 82728 3596
rect 82780 3584 82786 3596
rect 87966 3584 87972 3596
rect 82780 3556 87972 3584
rect 82780 3544 82786 3556
rect 87966 3544 87972 3556
rect 88024 3544 88030 3596
rect 90818 3544 90824 3596
rect 90876 3584 90882 3596
rect 123478 3584 123484 3596
rect 90876 3556 123484 3584
rect 90876 3544 90882 3556
rect 123478 3544 123484 3556
rect 123536 3544 123542 3596
rect 153010 3544 153016 3596
rect 153068 3544 153074 3596
rect 153102 3544 153108 3596
rect 153160 3584 153166 3596
rect 372890 3584 372896 3596
rect 153160 3556 372896 3584
rect 153160 3544 153166 3556
rect 372890 3544 372896 3556
rect 372948 3544 372954 3596
rect 373994 3544 374000 3596
rect 374052 3584 374058 3596
rect 375282 3584 375288 3596
rect 374052 3556 375288 3584
rect 374052 3544 374058 3556
rect 375282 3544 375288 3556
rect 375340 3544 375346 3596
rect 2924 3488 55996 3516
rect 2924 3476 2930 3488
rect 56042 3476 56048 3528
rect 56100 3516 56106 3528
rect 57146 3516 57152 3528
rect 56100 3488 57152 3516
rect 56100 3476 56106 3488
rect 57146 3476 57152 3488
rect 57204 3476 57210 3528
rect 58434 3476 58440 3528
rect 58492 3516 58498 3528
rect 59262 3516 59268 3528
rect 58492 3488 59268 3516
rect 58492 3476 58498 3488
rect 59262 3476 59268 3488
rect 59320 3476 59326 3528
rect 59630 3476 59636 3528
rect 59688 3516 59694 3528
rect 60642 3516 60648 3528
rect 59688 3488 60648 3516
rect 59688 3476 59694 3488
rect 60642 3476 60648 3488
rect 60700 3476 60706 3528
rect 63218 3476 63224 3528
rect 63276 3516 63282 3528
rect 74718 3516 74724 3528
rect 63276 3488 74724 3516
rect 63276 3476 63282 3488
rect 74718 3476 74724 3488
rect 74776 3476 74782 3528
rect 76190 3476 76196 3528
rect 76248 3516 76254 3528
rect 77202 3516 77208 3528
rect 76248 3488 77208 3516
rect 76248 3476 76254 3488
rect 77202 3476 77208 3488
rect 77260 3476 77266 3528
rect 79134 3476 79140 3528
rect 79192 3516 79198 3528
rect 79686 3516 79692 3528
rect 79192 3488 79692 3516
rect 79192 3476 79198 3488
rect 79686 3476 79692 3488
rect 79744 3476 79750 3528
rect 81342 3476 81348 3528
rect 81400 3516 81406 3528
rect 84470 3516 84476 3528
rect 81400 3488 84476 3516
rect 81400 3476 81406 3488
rect 84470 3476 84476 3488
rect 84528 3476 84534 3528
rect 87598 3476 87604 3528
rect 87656 3516 87662 3528
rect 89162 3516 89168 3528
rect 87656 3488 89168 3516
rect 87656 3476 87662 3488
rect 89162 3476 89168 3488
rect 89220 3476 89226 3528
rect 90910 3476 90916 3528
rect 90968 3516 90974 3528
rect 124674 3516 124680 3528
rect 90968 3488 124680 3516
rect 90968 3476 90974 3488
rect 124674 3476 124680 3488
rect 124732 3476 124738 3528
rect 137278 3476 137284 3528
rect 137336 3516 137342 3528
rect 140038 3516 140044 3528
rect 137336 3488 140044 3516
rect 137336 3476 137342 3488
rect 140038 3476 140044 3488
rect 140096 3476 140102 3528
rect 153028 3516 153056 3544
rect 376478 3516 376484 3528
rect 153028 3488 376484 3516
rect 376478 3476 376484 3488
rect 376536 3476 376542 3528
rect 398834 3476 398840 3528
rect 398892 3516 398898 3528
rect 400122 3516 400128 3528
rect 398892 3488 400128 3516
rect 398892 3476 398898 3488
rect 400122 3476 400128 3488
rect 400180 3476 400186 3528
rect 414658 3476 414664 3528
rect 414716 3516 414722 3528
rect 416682 3516 416688 3528
rect 414716 3488 416688 3516
rect 414716 3476 414722 3488
rect 416682 3476 416688 3488
rect 416740 3476 416746 3528
rect 423766 3476 423772 3528
rect 423824 3516 423830 3528
rect 424962 3516 424968 3528
rect 423824 3488 424968 3516
rect 423824 3476 423830 3488
rect 424962 3476 424968 3488
rect 425020 3476 425026 3528
rect 425698 3476 425704 3528
rect 425756 3516 425762 3528
rect 427262 3516 427268 3528
rect 425756 3488 427268 3516
rect 425756 3476 425762 3488
rect 427262 3476 427268 3488
rect 427320 3476 427326 3528
rect 448514 3476 448520 3528
rect 448572 3516 448578 3528
rect 449802 3516 449808 3528
rect 448572 3488 449808 3516
rect 448572 3476 448578 3488
rect 449802 3476 449808 3488
rect 449860 3476 449866 3528
rect 449912 3516 449940 3624
rect 450004 3584 450032 3692
rect 454678 3680 454684 3732
rect 454736 3720 454742 3732
rect 494698 3720 494704 3732
rect 454736 3692 494704 3720
rect 454736 3680 454742 3692
rect 494698 3680 494704 3692
rect 494756 3680 494762 3732
rect 450538 3612 450544 3664
rect 450596 3652 450602 3664
rect 491110 3652 491116 3664
rect 450596 3624 491116 3652
rect 450596 3612 450602 3624
rect 491110 3612 491116 3624
rect 491168 3612 491174 3664
rect 537478 3612 537484 3664
rect 537536 3652 537542 3664
rect 550266 3652 550272 3664
rect 537536 3624 550272 3652
rect 537536 3612 537542 3624
rect 550266 3612 550272 3624
rect 550324 3612 550330 3664
rect 481542 3584 481548 3596
rect 450004 3556 481548 3584
rect 481542 3544 481548 3556
rect 481600 3544 481606 3596
rect 481634 3544 481640 3596
rect 481692 3584 481698 3596
rect 482830 3584 482836 3596
rect 481692 3556 482836 3584
rect 481692 3544 481698 3556
rect 482830 3544 482836 3556
rect 482888 3544 482894 3596
rect 517146 3584 517152 3596
rect 509206 3556 517152 3584
rect 509206 3516 509234 3556
rect 517146 3544 517152 3556
rect 517204 3544 517210 3596
rect 544378 3544 544384 3596
rect 544436 3584 544442 3596
rect 557350 3584 557356 3596
rect 544436 3556 557356 3584
rect 544436 3544 544442 3556
rect 557350 3544 557356 3556
rect 557408 3544 557414 3596
rect 449912 3488 509234 3516
rect 512638 3476 512644 3528
rect 512696 3516 512702 3528
rect 513558 3516 513564 3528
rect 512696 3488 513564 3516
rect 512696 3476 512702 3488
rect 513558 3476 513564 3488
rect 513616 3476 513622 3528
rect 526438 3476 526444 3528
rect 526496 3516 526502 3528
rect 527818 3516 527824 3528
rect 526496 3488 527824 3516
rect 526496 3476 526502 3488
rect 527818 3476 527824 3488
rect 527876 3476 527882 3528
rect 530578 3476 530584 3528
rect 530636 3516 530642 3528
rect 531314 3516 531320 3528
rect 530636 3488 531320 3516
rect 530636 3476 530642 3488
rect 531314 3476 531320 3488
rect 531372 3476 531378 3528
rect 533338 3476 533344 3528
rect 533396 3516 533402 3528
rect 553762 3516 553768 3528
rect 533396 3488 553768 3516
rect 533396 3476 533402 3488
rect 553762 3476 553768 3488
rect 553820 3476 553826 3528
rect 572714 3476 572720 3528
rect 572772 3516 572778 3528
rect 573910 3516 573916 3528
rect 572772 3488 573916 3516
rect 572772 3476 572778 3488
rect 573910 3476 573916 3488
rect 573968 3476 573974 3528
rect 1670 3408 1676 3460
rect 1728 3448 1734 3460
rect 59538 3448 59544 3460
rect 1728 3420 59544 3448
rect 1728 3408 1734 3420
rect 59538 3408 59544 3420
rect 59596 3408 59602 3460
rect 65518 3408 65524 3460
rect 65576 3448 65582 3460
rect 66162 3448 66168 3460
rect 65576 3420 66168 3448
rect 65576 3408 65582 3420
rect 66162 3408 66168 3420
rect 66220 3408 66226 3460
rect 66714 3408 66720 3460
rect 66772 3448 66778 3460
rect 67542 3448 67548 3460
rect 66772 3420 67548 3448
rect 66772 3408 66778 3420
rect 67542 3408 67548 3420
rect 67600 3408 67606 3460
rect 67910 3408 67916 3460
rect 67968 3448 67974 3460
rect 68922 3448 68928 3460
rect 67968 3420 68928 3448
rect 67968 3408 67974 3420
rect 68922 3408 68928 3420
rect 68980 3408 68986 3460
rect 72602 3408 72608 3460
rect 72660 3448 72666 3460
rect 73062 3448 73068 3460
rect 72660 3420 73068 3448
rect 72660 3408 72666 3420
rect 73062 3408 73068 3420
rect 73120 3408 73126 3460
rect 82630 3408 82636 3460
rect 82688 3448 82694 3460
rect 91554 3448 91560 3460
rect 82688 3420 91560 3448
rect 82688 3408 82694 3420
rect 91554 3408 91560 3420
rect 91612 3408 91618 3460
rect 92382 3408 92388 3460
rect 92440 3448 92446 3460
rect 131758 3448 131764 3460
rect 92440 3420 131764 3448
rect 92440 3408 92446 3420
rect 131758 3408 131764 3420
rect 131816 3408 131822 3460
rect 148318 3408 148324 3460
rect 148376 3448 148382 3460
rect 150618 3448 150624 3460
rect 148376 3420 150624 3448
rect 148376 3408 148382 3420
rect 150618 3408 150624 3420
rect 150676 3408 150682 3460
rect 154482 3408 154488 3460
rect 154540 3448 154546 3460
rect 379974 3448 379980 3460
rect 154540 3420 379980 3448
rect 154540 3408 154546 3420
rect 379974 3408 379980 3420
rect 380032 3408 380038 3460
rect 429838 3408 429844 3460
rect 429896 3448 429902 3460
rect 583386 3448 583392 3460
rect 429896 3420 583392 3448
rect 429896 3408 429902 3420
rect 583386 3408 583392 3420
rect 583444 3408 583450 3460
rect 8754 3340 8760 3392
rect 8812 3380 8818 3392
rect 9582 3380 9588 3392
rect 8812 3352 9588 3380
rect 8812 3340 8818 3352
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 9950 3340 9956 3392
rect 10008 3380 10014 3392
rect 10962 3380 10968 3392
rect 10008 3352 10968 3380
rect 10008 3340 10014 3352
rect 10962 3340 10968 3352
rect 11020 3340 11026 3392
rect 11146 3340 11152 3392
rect 11204 3380 11210 3392
rect 12342 3380 12348 3392
rect 11204 3352 12348 3380
rect 11204 3340 11210 3352
rect 12342 3340 12348 3352
rect 12400 3340 12406 3392
rect 17034 3340 17040 3392
rect 17092 3380 17098 3392
rect 17862 3380 17868 3392
rect 17092 3352 17868 3380
rect 17092 3340 17098 3352
rect 17862 3340 17868 3352
rect 17920 3340 17926 3392
rect 23014 3340 23020 3392
rect 23072 3380 23078 3392
rect 28994 3380 29000 3392
rect 23072 3352 29000 3380
rect 23072 3340 23078 3352
rect 28994 3340 29000 3352
rect 29052 3340 29058 3392
rect 32398 3340 32404 3392
rect 32456 3380 32462 3392
rect 33042 3380 33048 3392
rect 32456 3352 33048 3380
rect 32456 3340 32462 3352
rect 33042 3340 33048 3352
rect 33100 3340 33106 3392
rect 33594 3340 33600 3392
rect 33652 3380 33658 3392
rect 34422 3380 34428 3392
rect 33652 3352 34428 3380
rect 33652 3340 33658 3352
rect 34422 3340 34428 3352
rect 34480 3340 34486 3392
rect 66346 3380 66352 3392
rect 34532 3352 66352 3380
rect 19426 3272 19432 3324
rect 19484 3312 19490 3324
rect 26878 3312 26884 3324
rect 19484 3284 26884 3312
rect 19484 3272 19490 3284
rect 26878 3272 26884 3284
rect 26936 3272 26942 3324
rect 28902 3272 28908 3324
rect 28960 3312 28966 3324
rect 34532 3312 34560 3352
rect 66346 3340 66352 3352
rect 66404 3340 66410 3392
rect 88058 3340 88064 3392
rect 88116 3380 88122 3392
rect 112806 3380 112812 3392
rect 88116 3352 112812 3380
rect 88116 3340 88122 3352
rect 112806 3340 112812 3352
rect 112864 3340 112870 3392
rect 136542 3340 136548 3392
rect 136600 3380 136606 3392
rect 306742 3380 306748 3392
rect 136600 3352 306748 3380
rect 136600 3340 136606 3352
rect 306742 3340 306748 3352
rect 306800 3340 306806 3392
rect 307754 3340 307760 3392
rect 307812 3380 307818 3392
rect 309042 3380 309048 3392
rect 307812 3352 309048 3380
rect 307812 3340 307818 3352
rect 309042 3340 309048 3352
rect 309100 3340 309106 3392
rect 316034 3340 316040 3392
rect 316092 3380 316098 3392
rect 317322 3380 317328 3392
rect 316092 3352 317328 3380
rect 316092 3340 316098 3352
rect 317322 3340 317328 3352
rect 317380 3340 317386 3392
rect 332594 3340 332600 3392
rect 332652 3380 332658 3392
rect 333882 3380 333888 3392
rect 332652 3352 333888 3380
rect 332652 3340 332658 3352
rect 333882 3340 333888 3352
rect 333940 3340 333946 3392
rect 347038 3340 347044 3392
rect 347096 3380 347102 3392
rect 349246 3380 349252 3392
rect 347096 3352 349252 3380
rect 347096 3340 347102 3352
rect 349246 3340 349252 3352
rect 349304 3340 349310 3392
rect 473354 3340 473360 3392
rect 473412 3380 473418 3392
rect 474550 3380 474556 3392
rect 473412 3352 474556 3380
rect 473412 3340 473418 3352
rect 474550 3340 474556 3352
rect 474608 3340 474614 3392
rect 481542 3340 481548 3392
rect 481600 3380 481606 3392
rect 487614 3380 487620 3392
rect 481600 3352 487620 3380
rect 481600 3340 481606 3352
rect 487614 3340 487620 3352
rect 487672 3340 487678 3392
rect 547874 3340 547880 3392
rect 547932 3380 547938 3392
rect 549070 3380 549076 3392
rect 547932 3352 549076 3380
rect 547932 3340 547938 3352
rect 549070 3340 549076 3352
rect 549128 3340 549134 3392
rect 28960 3284 34560 3312
rect 28960 3272 28966 3284
rect 34790 3272 34796 3324
rect 34848 3312 34854 3324
rect 35802 3312 35808 3324
rect 34848 3284 35808 3312
rect 34848 3272 34854 3284
rect 35802 3272 35808 3284
rect 35860 3272 35866 3324
rect 40678 3272 40684 3324
rect 40736 3312 40742 3324
rect 41322 3312 41328 3324
rect 40736 3284 41328 3312
rect 40736 3272 40742 3284
rect 41322 3272 41328 3284
rect 41380 3272 41386 3324
rect 41874 3272 41880 3324
rect 41932 3312 41938 3324
rect 43438 3312 43444 3324
rect 41932 3284 43444 3312
rect 41932 3272 41938 3284
rect 43438 3272 43444 3284
rect 43496 3272 43502 3324
rect 44266 3272 44272 3324
rect 44324 3312 44330 3324
rect 45370 3312 45376 3324
rect 44324 3284 45376 3312
rect 44324 3272 44330 3284
rect 45370 3272 45376 3284
rect 45428 3272 45434 3324
rect 45462 3272 45468 3324
rect 45520 3312 45526 3324
rect 66530 3312 66536 3324
rect 45520 3284 66536 3312
rect 45520 3272 45526 3284
rect 66530 3272 66536 3284
rect 66588 3272 66594 3324
rect 88150 3272 88156 3324
rect 88208 3312 88214 3324
rect 111610 3312 111616 3324
rect 88208 3284 111616 3312
rect 88208 3272 88214 3284
rect 111610 3272 111616 3284
rect 111668 3272 111674 3324
rect 136358 3272 136364 3324
rect 136416 3312 136422 3324
rect 305546 3312 305552 3324
rect 136416 3284 305552 3312
rect 136416 3272 136422 3284
rect 305546 3272 305552 3284
rect 305604 3272 305610 3324
rect 31294 3204 31300 3256
rect 31352 3244 31358 3256
rect 67818 3244 67824 3256
rect 31352 3216 67824 3244
rect 31352 3204 31358 3216
rect 67818 3204 67824 3216
rect 67876 3204 67882 3256
rect 86770 3204 86776 3256
rect 86828 3244 86834 3256
rect 109310 3244 109316 3256
rect 86828 3216 109316 3244
rect 86828 3204 86834 3216
rect 109310 3204 109316 3216
rect 109368 3204 109374 3256
rect 193214 3204 193220 3256
rect 193272 3244 193278 3256
rect 194410 3244 194416 3256
rect 193272 3216 194416 3244
rect 193272 3204 193278 3216
rect 194410 3204 194416 3216
rect 194468 3204 194474 3256
rect 203518 3204 203524 3256
rect 203576 3244 203582 3256
rect 206186 3244 206192 3256
rect 203576 3216 206192 3244
rect 203576 3204 203582 3216
rect 206186 3204 206192 3216
rect 206244 3204 206250 3256
rect 220078 3204 220084 3256
rect 220136 3244 220142 3256
rect 387150 3244 387156 3256
rect 220136 3216 387156 3244
rect 220136 3204 220142 3216
rect 387150 3204 387156 3216
rect 387208 3204 387214 3256
rect 30098 3136 30104 3188
rect 30156 3176 30162 3188
rect 45370 3176 45376 3188
rect 30156 3148 45376 3176
rect 30156 3136 30162 3148
rect 45370 3136 45376 3148
rect 45428 3136 45434 3188
rect 69198 3176 69204 3188
rect 45480 3148 69204 3176
rect 26510 3068 26516 3120
rect 26568 3108 26574 3120
rect 27522 3108 27528 3120
rect 26568 3080 27528 3108
rect 26568 3068 26574 3080
rect 27522 3068 27528 3080
rect 27580 3068 27586 3120
rect 37182 3068 37188 3120
rect 37240 3108 37246 3120
rect 45480 3108 45508 3148
rect 69198 3136 69204 3148
rect 69256 3136 69262 3188
rect 86862 3136 86868 3188
rect 86920 3176 86926 3188
rect 108114 3176 108120 3188
rect 86920 3148 108120 3176
rect 86920 3136 86926 3148
rect 108114 3136 108120 3148
rect 108172 3136 108178 3188
rect 123570 3136 123576 3188
rect 123628 3176 123634 3188
rect 125870 3176 125876 3188
rect 123628 3148 125876 3176
rect 123628 3136 123634 3148
rect 125870 3136 125876 3148
rect 125928 3136 125934 3188
rect 131022 3136 131028 3188
rect 131080 3176 131086 3188
rect 284294 3176 284300 3188
rect 131080 3148 284300 3176
rect 131080 3136 131086 3148
rect 284294 3136 284300 3148
rect 284352 3136 284358 3188
rect 37240 3080 45508 3108
rect 37240 3068 37246 3080
rect 48958 3068 48964 3120
rect 49016 3108 49022 3120
rect 49602 3108 49608 3120
rect 49016 3080 49608 3108
rect 49016 3068 49022 3080
rect 49602 3068 49608 3080
rect 49660 3068 49666 3120
rect 50154 3068 50160 3120
rect 50212 3108 50218 3120
rect 50982 3108 50988 3120
rect 50212 3080 50988 3108
rect 50212 3068 50218 3080
rect 50982 3068 50988 3080
rect 51040 3068 51046 3120
rect 52546 3068 52552 3120
rect 52604 3108 52610 3120
rect 53650 3108 53656 3120
rect 52604 3080 53656 3108
rect 52604 3068 52610 3080
rect 53650 3068 53656 3080
rect 53708 3068 53714 3120
rect 68002 3108 68008 3120
rect 53760 3080 68008 3108
rect 25314 3000 25320 3052
rect 25372 3040 25378 3052
rect 26142 3040 26148 3052
rect 25372 3012 26148 3040
rect 25372 3000 25378 3012
rect 26142 3000 26148 3012
rect 26200 3000 26206 3052
rect 35986 3000 35992 3052
rect 36044 3040 36050 3052
rect 53760 3040 53788 3080
rect 68002 3068 68008 3080
rect 68060 3068 68066 3120
rect 86678 3068 86684 3120
rect 86736 3108 86742 3120
rect 105722 3108 105728 3120
rect 86736 3080 105728 3108
rect 86736 3068 86742 3080
rect 105722 3068 105728 3080
rect 105780 3068 105786 3120
rect 128262 3068 128268 3120
rect 128320 3108 128326 3120
rect 272426 3108 272432 3120
rect 128320 3080 272432 3108
rect 128320 3068 128326 3080
rect 272426 3068 272432 3080
rect 272484 3068 272490 3120
rect 417510 3068 417516 3120
rect 417568 3108 417574 3120
rect 420178 3108 420184 3120
rect 417568 3080 420184 3108
rect 417568 3068 417574 3080
rect 420178 3068 420184 3080
rect 420236 3068 420242 3120
rect 36044 3012 53788 3040
rect 36044 3000 36050 3012
rect 53834 3000 53840 3052
rect 53892 3040 53898 3052
rect 70578 3040 70584 3052
rect 53892 3012 70584 3040
rect 53892 3000 53898 3012
rect 70578 3000 70584 3012
rect 70636 3000 70642 3052
rect 74994 3000 75000 3052
rect 75052 3040 75058 3052
rect 76650 3040 76656 3052
rect 75052 3012 76656 3040
rect 75052 3000 75058 3012
rect 76650 3000 76656 3012
rect 76708 3000 76714 3052
rect 85482 3000 85488 3052
rect 85540 3040 85546 3052
rect 102226 3040 102232 3052
rect 85540 3012 102232 3040
rect 85540 3000 85546 3012
rect 102226 3000 102232 3012
rect 102284 3000 102290 3052
rect 104158 3000 104164 3052
rect 104216 3040 104222 3052
rect 121086 3040 121092 3052
rect 104216 3012 121092 3040
rect 104216 3000 104222 3012
rect 121086 3000 121092 3012
rect 121144 3000 121150 3052
rect 222930 3000 222936 3052
rect 222988 3040 222994 3052
rect 350442 3040 350448 3052
rect 222988 3012 350448 3040
rect 222988 3000 222994 3012
rect 350442 3000 350448 3012
rect 350500 3000 350506 3052
rect 407758 3000 407764 3052
rect 407816 3040 407822 3052
rect 409598 3040 409604 3052
rect 407816 3012 409604 3040
rect 407816 3000 407822 3012
rect 409598 3000 409604 3012
rect 409656 3000 409662 3052
rect 45462 2932 45468 2984
rect 45520 2972 45526 2984
rect 70670 2972 70676 2984
rect 45520 2944 70676 2972
rect 45520 2932 45526 2944
rect 70670 2932 70676 2944
rect 70728 2932 70734 2984
rect 84102 2932 84108 2984
rect 84160 2972 84166 2984
rect 95142 2972 95148 2984
rect 84160 2944 95148 2972
rect 84160 2932 84166 2944
rect 95142 2932 95148 2944
rect 95200 2932 95206 2984
rect 102870 2932 102876 2984
rect 102928 2972 102934 2984
rect 117590 2972 117596 2984
rect 102928 2944 117596 2972
rect 102928 2932 102934 2944
rect 117590 2932 117596 2944
rect 117648 2932 117654 2984
rect 220262 2932 220268 2984
rect 220320 2972 220326 2984
rect 337470 2972 337476 2984
rect 220320 2944 337476 2972
rect 220320 2932 220326 2944
rect 337470 2932 337476 2944
rect 337528 2932 337534 2984
rect 368474 2932 368480 2984
rect 368532 2972 368538 2984
rect 371694 2972 371700 2984
rect 368532 2944 371700 2972
rect 368532 2932 368538 2944
rect 371694 2932 371700 2944
rect 371752 2932 371758 2984
rect 51350 2864 51356 2916
rect 51408 2904 51414 2916
rect 72050 2904 72056 2916
rect 51408 2876 72056 2904
rect 51408 2864 51414 2876
rect 72050 2864 72056 2876
rect 72108 2864 72114 2916
rect 81250 2864 81256 2916
rect 81308 2904 81314 2916
rect 82078 2904 82084 2916
rect 81308 2876 82084 2904
rect 81308 2864 81314 2876
rect 82078 2864 82084 2876
rect 82136 2864 82142 2916
rect 83918 2864 83924 2916
rect 83976 2904 83982 2916
rect 92750 2904 92756 2916
rect 83976 2876 92756 2904
rect 83976 2864 83982 2876
rect 92750 2864 92756 2876
rect 92808 2864 92814 2916
rect 94406 2864 94412 2916
rect 94464 2904 94470 2916
rect 98638 2904 98644 2916
rect 94464 2876 98644 2904
rect 94464 2864 94470 2876
rect 98638 2864 98644 2876
rect 98696 2864 98702 2916
rect 102778 2864 102784 2916
rect 102836 2904 102842 2916
rect 110506 2904 110512 2916
rect 102836 2876 110512 2904
rect 102836 2864 102842 2876
rect 110506 2864 110512 2876
rect 110564 2864 110570 2916
rect 222838 2864 222844 2916
rect 222896 2904 222902 2916
rect 294874 2904 294880 2916
rect 222896 2876 294880 2904
rect 222896 2864 222902 2876
rect 294874 2864 294880 2876
rect 294932 2864 294938 2916
rect 519630 2864 519636 2916
rect 519688 2904 519694 2916
rect 524230 2904 524236 2916
rect 519688 2876 524236 2904
rect 519688 2864 519694 2876
rect 524230 2864 524236 2876
rect 524288 2864 524294 2916
rect 43070 2796 43076 2848
rect 43128 2836 43134 2848
rect 53834 2836 53840 2848
rect 43128 2808 53840 2836
rect 43128 2796 43134 2808
rect 53834 2796 53840 2808
rect 53892 2796 53898 2848
rect 57238 2796 57244 2848
rect 57296 2836 57302 2848
rect 68278 2836 68284 2848
rect 57296 2808 68284 2836
rect 57296 2796 57302 2808
rect 68278 2796 68284 2808
rect 68336 2796 68342 2848
rect 81066 2796 81072 2848
rect 81124 2836 81130 2848
rect 86862 2836 86868 2848
rect 81124 2808 86868 2836
rect 81124 2796 81130 2808
rect 86862 2796 86868 2808
rect 86920 2796 86926 2848
rect 101398 2796 101404 2848
rect 101456 2836 101462 2848
rect 106918 2836 106924 2848
rect 101456 2808 106924 2836
rect 101456 2796 101462 2808
rect 106918 2796 106924 2808
rect 106976 2796 106982 2848
rect 223022 2796 223028 2848
rect 223080 2836 223086 2848
rect 283098 2836 283104 2848
rect 223080 2808 283104 2836
rect 223080 2796 223086 2808
rect 283098 2796 283104 2808
rect 283156 2796 283162 2848
rect 242894 2728 242900 2780
rect 242952 2768 242958 2780
rect 244090 2768 244096 2780
rect 242952 2740 244096 2768
rect 242952 2728 242958 2740
rect 244090 2728 244096 2740
rect 244148 2728 244154 2780
rect 160002 2116 160008 2168
rect 160060 2156 160066 2168
rect 401318 2156 401324 2168
rect 160060 2128 401324 2156
rect 160060 2116 160066 2128
rect 401318 2116 401324 2128
rect 401376 2116 401382 2168
rect 179046 2048 179052 2100
rect 179104 2088 179110 2100
rect 479334 2088 479340 2100
rect 179104 2060 479340 2088
rect 179104 2048 179110 2060
rect 479334 2048 479340 2060
rect 479392 2048 479398 2100
<< via1 >>
rect 201500 702992 201552 703044
rect 202788 702992 202840 703044
rect 209136 700816 209188 700868
rect 218980 700816 219032 700868
rect 198004 700748 198056 700800
rect 235172 700748 235224 700800
rect 206284 700680 206336 700732
rect 267648 700680 267700 700732
rect 200764 700612 200816 700664
rect 283840 700612 283892 700664
rect 204904 700544 204956 700596
rect 300124 700544 300176 700596
rect 385684 700544 385736 700596
rect 462320 700544 462372 700596
rect 213184 700476 213236 700528
rect 332508 700476 332560 700528
rect 388444 700476 388496 700528
rect 397460 700476 397512 700528
rect 400864 700476 400916 700528
rect 478512 700476 478564 700528
rect 215944 700408 215996 700460
rect 348792 700408 348844 700460
rect 370504 700408 370556 700460
rect 494796 700408 494848 700460
rect 40500 700340 40552 700392
rect 41328 700340 41380 700392
rect 170312 700340 170364 700392
rect 196532 700340 196584 700392
rect 214564 700340 214616 700392
rect 364984 700340 365036 700392
rect 382924 700340 382976 700392
rect 527180 700340 527232 700392
rect 24308 700272 24360 700324
rect 33784 700272 33836 700324
rect 58808 700272 58860 700324
rect 72976 700272 73028 700324
rect 137836 700272 137888 700324
rect 146944 700272 146996 700324
rect 154120 700272 154172 700324
rect 196624 700272 196676 700324
rect 209044 700272 209096 700324
rect 559656 700272 559708 700324
rect 88340 699660 88392 699712
rect 89168 699660 89220 699712
rect 104900 699660 104952 699712
rect 105452 699660 105504 699712
rect 381544 696940 381596 696992
rect 580172 696940 580224 696992
rect 2780 683680 2832 683732
rect 4804 683680 4856 683732
rect 399484 683136 399536 683188
rect 580172 683136 580224 683188
rect 146944 677492 146996 677544
rect 153844 677492 153896 677544
rect 3516 670692 3568 670744
rect 35164 670692 35216 670744
rect 206376 670692 206428 670744
rect 580172 670692 580224 670744
rect 153844 661036 153896 661088
rect 159364 661036 159416 661088
rect 3424 656888 3476 656940
rect 15844 656888 15896 656940
rect 159364 652672 159416 652724
rect 162768 652672 162820 652724
rect 162768 648864 162820 648916
rect 166264 648864 166316 648916
rect 377404 643084 377456 643136
rect 580172 643084 580224 643136
rect 166264 639548 166316 639600
rect 175924 639548 175976 639600
rect 3424 632068 3476 632120
rect 14464 632068 14516 632120
rect 396724 630640 396776 630692
rect 580172 630640 580224 630692
rect 3148 618264 3200 618316
rect 36544 618264 36596 618316
rect 175924 617516 175976 617568
rect 186964 617516 187016 617568
rect 367744 616836 367796 616888
rect 580172 616836 580224 616888
rect 3240 605820 3292 605872
rect 22744 605820 22796 605872
rect 186964 597456 187016 597508
rect 189724 597456 189776 597508
rect 376024 590656 376076 590708
rect 579804 590656 579856 590708
rect 3332 579640 3384 579692
rect 11704 579640 11756 579692
rect 395344 576852 395396 576904
rect 580172 576852 580224 576904
rect 189724 566448 189776 566500
rect 196900 566448 196952 566500
rect 3424 565836 3476 565888
rect 39304 565836 39356 565888
rect 363604 563048 363656 563100
rect 579804 563048 579856 563100
rect 3424 553392 3476 553444
rect 25504 553392 25556 553444
rect 378784 536800 378836 536852
rect 580172 536800 580224 536852
rect 3424 527144 3476 527196
rect 17224 527144 17276 527196
rect 393964 524424 394016 524476
rect 580172 524424 580224 524476
rect 3424 514768 3476 514820
rect 43444 514768 43496 514820
rect 360844 510620 360896 510672
rect 580172 510620 580224 510672
rect 3056 500964 3108 501016
rect 29644 500964 29696 501016
rect 374644 484372 374696 484424
rect 580172 484372 580224 484424
rect 3424 474716 3476 474768
rect 18604 474716 18656 474768
rect 392584 470568 392636 470620
rect 579988 470568 580040 470620
rect 3240 462340 3292 462392
rect 47584 462340 47636 462392
rect 358084 456764 358136 456816
rect 580172 456764 580224 456816
rect 3148 448536 3200 448588
rect 32404 448536 32456 448588
rect 206468 434732 206520 434784
rect 216680 434732 216732 434784
rect 202236 433304 202288 433356
rect 216680 433304 216732 433356
rect 213276 432352 213328 432404
rect 216680 432352 216732 432404
rect 389824 430584 389876 430636
rect 580172 430584 580224 430636
rect 204996 429156 205048 429208
rect 216680 429156 216732 429208
rect 3424 422288 3476 422340
rect 21364 422288 21416 422340
rect 3148 409844 3200 409896
rect 50344 409844 50396 409896
rect 211804 409844 211856 409896
rect 216680 409844 216732 409896
rect 371884 404336 371936 404388
rect 580172 404336 580224 404388
rect 219716 403044 219768 403096
rect 219900 403044 219952 403096
rect 59360 400052 59412 400104
rect 217324 400052 217376 400104
rect 122748 399984 122800 400036
rect 209136 399984 209188 400036
rect 115756 399916 115808 399968
rect 213184 399916 213236 399968
rect 218980 399916 219032 399968
rect 227352 399916 227404 399968
rect 115664 399848 115716 399900
rect 215944 399848 215996 399900
rect 218612 399848 218664 399900
rect 226432 399848 226484 399900
rect 53472 399780 53524 399832
rect 199016 399780 199068 399832
rect 218428 399780 218480 399832
rect 226524 399780 226576 399832
rect 52276 399712 52328 399764
rect 217232 399712 217284 399764
rect 217508 399712 217560 399764
rect 233240 399712 233292 399764
rect 57796 399644 57848 399696
rect 172520 399644 172572 399696
rect 187608 399644 187660 399696
rect 357532 399644 357584 399696
rect 57888 399576 57940 399628
rect 232044 399576 232096 399628
rect 57704 399508 57756 399560
rect 233424 399508 233476 399560
rect 249156 399508 249208 399560
rect 359004 399508 359056 399560
rect 57336 399440 57388 399492
rect 233332 399440 233384 399492
rect 246304 399440 246356 399492
rect 359096 399440 359148 399492
rect 58808 399372 58860 399424
rect 125600 399372 125652 399424
rect 191748 399372 191800 399424
rect 206468 399372 206520 399424
rect 188988 399304 189040 399356
rect 202236 399304 202288 399356
rect 219532 398624 219584 398676
rect 224960 398624 225012 398676
rect 219624 398556 219676 398608
rect 224776 398556 224828 398608
rect 219440 398420 219492 398472
rect 224868 398420 224920 398472
rect 175188 398216 175240 398268
rect 211804 398216 211856 398268
rect 217692 398216 217744 398268
rect 227904 398284 227956 398336
rect 125508 398148 125560 398200
rect 196624 398148 196676 398200
rect 217600 398148 217652 398200
rect 227996 398216 228048 398268
rect 219716 398148 219768 398200
rect 227812 398148 227864 398200
rect 119988 398080 120040 398132
rect 198004 398080 198056 398132
rect 217784 398080 217836 398132
rect 220084 398080 220136 398132
rect 228088 398080 228140 398132
rect 228180 397944 228232 397996
rect 3424 397468 3476 397520
rect 146300 397468 146352 397520
rect 87696 397332 87748 397384
rect 229100 397332 229152 397384
rect 61476 397264 61528 397316
rect 265164 397264 265216 397316
rect 300124 397264 300176 397316
rect 308588 397264 308640 397316
rect 83280 397196 83332 397248
rect 225052 397196 225104 397248
rect 238024 397196 238076 397248
rect 239220 397196 239272 397248
rect 61752 397128 61804 397180
rect 273260 397128 273312 397180
rect 62764 397060 62816 397112
rect 278044 397060 278096 397112
rect 58440 396992 58492 397044
rect 113180 396992 113232 397044
rect 114468 396992 114520 397044
rect 137284 396992 137336 397044
rect 78312 396924 78364 396976
rect 170404 396924 170456 396976
rect 183468 396924 183520 396976
rect 228272 396924 228324 396976
rect 92296 396856 92348 396908
rect 189080 396856 189132 396908
rect 191104 396856 191156 396908
rect 236184 396856 236236 396908
rect 93492 396788 93544 396840
rect 193220 396788 193272 396840
rect 196624 396788 196676 396840
rect 241612 396788 241664 396840
rect 109776 396720 109828 396772
rect 231952 396720 232004 396772
rect 244924 396720 244976 396772
rect 247132 396720 247184 396772
rect 264244 396720 264296 396772
rect 265256 396720 265308 396772
rect 269764 396720 269816 396772
rect 272524 396720 272576 396772
rect 282184 396720 282236 396772
rect 283564 396720 283616 396772
rect 58532 396652 58584 396704
rect 103704 396652 103756 396704
rect 105912 396652 105964 396704
rect 231860 396652 231912 396704
rect 242256 396652 242308 396704
rect 101864 396584 101916 396636
rect 230572 396584 230624 396636
rect 242164 396584 242216 396636
rect 247684 396584 247736 396636
rect 253204 396652 253256 396704
rect 254492 396652 254544 396704
rect 262864 396652 262916 396704
rect 263876 396652 263928 396704
rect 284944 396652 284996 396704
rect 285956 396652 286008 396704
rect 307024 396652 307076 396704
rect 315764 396652 315816 396704
rect 274732 396584 274784 396636
rect 79968 396516 80020 396568
rect 98644 396516 98696 396568
rect 100116 396516 100168 396568
rect 230480 396516 230532 396568
rect 238116 396516 238168 396568
rect 273628 396516 273680 396568
rect 61660 396448 61712 396500
rect 88708 396448 88760 396500
rect 98920 396448 98972 396500
rect 229192 396448 229244 396500
rect 233976 396448 234028 396500
rect 271144 396448 271196 396500
rect 58808 396380 58860 396432
rect 86500 396380 86552 396432
rect 226984 396380 227036 396432
rect 263600 396380 263652 396432
rect 59912 396312 59964 396364
rect 80428 396312 80480 396364
rect 101588 396312 101640 396364
rect 112444 396312 112496 396364
rect 220084 396312 220136 396364
rect 310980 396312 311032 396364
rect 59544 396244 59596 396296
rect 252652 396244 252704 396296
rect 258724 396244 258776 396296
rect 342260 396244 342312 396296
rect 102876 396176 102928 396228
rect 107016 396176 107068 396228
rect 263600 396176 263652 396228
rect 276388 396176 276440 396228
rect 276664 396176 276716 396228
rect 298468 396176 298520 396228
rect 111616 396108 111668 396160
rect 119344 396108 119396 396160
rect 249064 396108 249116 396160
rect 262036 396108 262088 396160
rect 291844 396108 291896 396160
rect 300860 396108 300912 396160
rect 96528 396040 96580 396092
rect 106924 396040 106976 396092
rect 107200 396040 107252 396092
rect 116584 396040 116636 396092
rect 304264 396040 304316 396092
rect 313372 396040 313424 396092
rect 183192 395972 183244 396024
rect 187700 395972 187752 396024
rect 232504 395972 232556 396024
rect 250076 395972 250128 396024
rect 179328 395904 179380 395956
rect 244464 395904 244516 395956
rect 113640 395836 113692 395888
rect 194600 395836 194652 395888
rect 233884 395836 233936 395888
rect 256148 395836 256200 395888
rect 138480 395768 138532 395820
rect 228548 395768 228600 395820
rect 231124 395768 231176 395820
rect 260932 395768 260984 395820
rect 56324 395700 56376 395752
rect 118148 395700 118200 395752
rect 136456 395700 136508 395752
rect 228456 395700 228508 395752
rect 235264 395700 235316 395752
rect 273444 395700 273496 395752
rect 54668 395632 54720 395684
rect 150716 395632 150768 395684
rect 177948 395632 178000 395684
rect 253572 395632 253624 395684
rect 54852 395564 54904 395616
rect 98460 395564 98512 395616
rect 115848 395564 115900 395616
rect 222200 395564 222252 395616
rect 224684 395564 224736 395616
rect 263600 395564 263652 395616
rect 96436 395496 96488 395548
rect 229284 395496 229336 395548
rect 231216 395496 231268 395548
rect 293316 395496 293368 395548
rect 52368 395428 52420 395480
rect 242900 395428 242952 395480
rect 52184 395360 52236 395412
rect 248604 395360 248656 395412
rect 54760 395292 54812 395344
rect 290188 395292 290240 395344
rect 193312 393252 193364 393304
rect 196900 393320 196952 393372
rect 219072 392912 219124 392964
rect 219348 392912 219400 392964
rect 191380 390328 191432 390380
rect 193312 390328 193364 390380
rect 186320 387812 186372 387864
rect 191380 387812 191432 387864
rect 185676 385636 185728 385688
rect 186320 385636 186372 385688
rect 219072 383732 219124 383784
rect 219348 383664 219400 383716
rect 183560 379516 183612 379568
rect 185676 379516 185728 379568
rect 85396 378768 85448 378820
rect 232136 378768 232188 378820
rect 85396 378156 85448 378208
rect 580172 378156 580224 378208
rect 177304 374620 177356 374672
rect 183560 374620 183612 374672
rect 3424 371220 3476 371272
rect 149060 371220 149112 371272
rect 86868 364352 86920 364404
rect 579620 364352 579672 364404
rect 173440 360136 173492 360188
rect 177304 360204 177356 360256
rect 171784 358504 171836 358556
rect 173440 358504 173492 358556
rect 119896 358028 119948 358080
rect 223580 358028 223632 358080
rect 3148 357416 3200 357468
rect 150440 357416 150492 357468
rect 170496 352044 170548 352096
rect 171784 352044 171836 352096
rect 84108 351908 84160 351960
rect 580172 351908 580224 351960
rect 3332 345040 3384 345092
rect 149152 345040 149204 345092
rect 166724 340892 166776 340944
rect 170496 340892 170548 340944
rect 162860 338036 162912 338088
rect 166724 338104 166776 338156
rect 219072 335112 219124 335164
rect 219348 335112 219400 335164
rect 156604 331168 156656 331220
rect 162860 331236 162912 331288
rect 219072 325796 219124 325848
rect 219348 325796 219400 325848
rect 82636 324300 82688 324352
rect 580172 324300 580224 324352
rect 155224 320424 155276 320476
rect 156604 320424 156656 320476
rect 131028 319404 131080 319456
rect 228732 319404 228784 319456
rect 3424 318792 3476 318844
rect 151820 318792 151872 318844
rect 84016 311856 84068 311908
rect 579988 311856 580040 311908
rect 154488 305600 154540 305652
rect 228364 305600 228416 305652
rect 3240 304988 3292 305040
rect 153200 304988 153252 305040
rect 153844 301520 153896 301572
rect 155224 301520 155276 301572
rect 191656 301452 191708 301504
rect 342352 301452 342404 301504
rect 97816 300092 97868 300144
rect 376024 300092 376076 300144
rect 95056 298732 95108 298784
rect 378784 298732 378836 298784
rect 81348 298120 81400 298172
rect 580172 298120 580224 298172
rect 18604 297372 18656 297424
rect 142160 297372 142212 297424
rect 112996 294652 113048 294704
rect 412640 294652 412692 294704
rect 107476 294584 107528 294636
rect 542360 294584 542412 294636
rect 3424 292544 3476 292596
rect 153292 292544 153344 292596
rect 14464 290436 14516 290488
rect 133880 290436 133932 290488
rect 111616 284928 111668 284980
rect 429200 284928 429252 284980
rect 152832 276020 152884 276072
rect 153844 276020 153896 276072
rect 79968 271872 80020 271924
rect 580172 271872 580224 271924
rect 144828 269764 144880 269816
rect 213920 269764 213972 269816
rect 150532 269084 150584 269136
rect 152832 269084 152884 269136
rect 52092 268336 52144 268388
rect 258172 268336 258224 268388
rect 176568 267044 176620 267096
rect 191104 267044 191156 267096
rect 98644 266976 98696 267028
rect 176660 266976 176712 267028
rect 182088 266976 182140 267028
rect 204996 266976 205048 267028
rect 213184 266976 213236 267028
rect 266452 266976 266504 267028
rect 3056 266364 3108 266416
rect 154580 266364 154632 266416
rect 112444 266296 112496 266348
rect 204260 266296 204312 266348
rect 116584 266228 116636 266280
rect 211160 266228 211212 266280
rect 107016 266160 107068 266212
rect 207020 266160 207072 266212
rect 101956 266092 102008 266144
rect 225144 266092 225196 266144
rect 107384 266024 107436 266076
rect 232412 266024 232464 266076
rect 82728 265956 82780 266008
rect 233516 265956 233568 266008
rect 77208 265888 77260 265940
rect 232228 265888 232280 265940
rect 57152 265820 57204 265872
rect 213276 265820 213328 265872
rect 52000 265752 52052 265804
rect 259552 265752 259604 265804
rect 61568 265684 61620 265736
rect 278780 265684 278832 265736
rect 56232 265616 56284 265668
rect 325700 265616 325752 265668
rect 137284 265548 137336 265600
rect 219440 265548 219492 265600
rect 111524 265480 111576 265532
rect 191840 265480 191892 265532
rect 197268 265480 197320 265532
rect 276112 265480 276164 265532
rect 195888 265412 195940 265464
rect 253204 265412 253256 265464
rect 50344 264868 50396 264920
rect 147772 264868 147824 264920
rect 47584 264800 47636 264852
rect 144920 264800 144972 264852
rect 43444 264732 43496 264784
rect 142252 264732 142304 264784
rect 164148 264732 164200 264784
rect 229376 264732 229428 264784
rect 97908 264664 97960 264716
rect 197544 264664 197596 264716
rect 209688 264664 209740 264716
rect 262864 264664 262916 264716
rect 93768 264596 93820 264648
rect 228640 264596 228692 264648
rect 95148 264528 95200 264580
rect 230664 264528 230716 264580
rect 91008 264460 91060 264512
rect 232320 264460 232372 264512
rect 234068 264460 234120 264512
rect 256700 264460 256752 264512
rect 54484 264392 54536 264444
rect 280160 264392 280212 264444
rect 54392 264324 54444 264376
rect 295340 264324 295392 264376
rect 54300 264256 54352 264308
rect 305000 264256 305052 264308
rect 89536 264188 89588 264240
rect 580264 264188 580316 264240
rect 35164 264120 35216 264172
rect 132500 264120 132552 264172
rect 133788 264120 133840 264172
rect 208400 264120 208452 264172
rect 119344 264052 119396 264104
rect 215300 264052 215352 264104
rect 106924 263984 106976 264036
rect 197452 263984 197504 264036
rect 56048 263916 56100 263968
rect 140780 263916 140832 263968
rect 126888 263848 126940 263900
rect 201684 263848 201736 263900
rect 149244 263576 149296 263628
rect 150532 263576 150584 263628
rect 29644 263508 29696 263560
rect 140780 263508 140832 263560
rect 213828 263508 213880 263560
rect 291844 263508 291896 263560
rect 8208 263440 8260 263492
rect 128360 263440 128412 263492
rect 181996 263440 182048 263492
rect 196624 263440 196676 263492
rect 205548 263440 205600 263492
rect 287060 263440 287112 263492
rect 108856 263372 108908 263424
rect 230848 263372 230900 263424
rect 235356 263372 235408 263424
rect 358820 263372 358872 263424
rect 111708 263304 111760 263356
rect 388444 263304 388496 263356
rect 108856 263236 108908 263288
rect 385684 263236 385736 263288
rect 102048 263168 102100 263220
rect 396724 263168 396776 263220
rect 104716 263100 104768 263152
rect 399484 263100 399536 263152
rect 97908 263032 97960 263084
rect 395344 263032 395396 263084
rect 95148 262964 95200 263016
rect 393964 262964 394016 263016
rect 92388 262896 92440 262948
rect 392584 262896 392636 262948
rect 88248 262828 88300 262880
rect 389824 262828 389876 262880
rect 32404 262760 32456 262812
rect 143540 262760 143592 262812
rect 201408 262760 201460 262812
rect 259460 262760 259512 262812
rect 39304 262692 39356 262744
rect 138020 262692 138072 262744
rect 36544 262624 36596 262676
rect 135260 262624 135312 262676
rect 33784 262556 33836 262608
rect 129740 262556 129792 262608
rect 55956 262488 56008 262540
rect 147680 262488 147732 262540
rect 118516 262420 118568 262472
rect 200764 262420 200816 262472
rect 129648 262352 129700 262404
rect 205640 262352 205692 262404
rect 11704 262148 11756 262200
rect 136640 262148 136692 262200
rect 146944 262148 146996 262200
rect 149244 262148 149296 262200
rect 202788 262148 202840 262200
rect 284944 262148 284996 262200
rect 21364 262080 21416 262132
rect 146392 262080 146444 262132
rect 170404 262080 170456 262132
rect 173900 262080 173952 262132
rect 218980 262080 219032 262132
rect 307024 262080 307076 262132
rect 53196 262012 53248 262064
rect 198924 262012 198976 262064
rect 222108 262012 222160 262064
rect 317420 262012 317472 262064
rect 108764 261944 108816 261996
rect 370504 261944 370556 261996
rect 99288 261876 99340 261928
rect 367744 261876 367796 261928
rect 100668 261808 100720 261860
rect 377404 261808 377456 261860
rect 106096 261740 106148 261792
rect 382924 261740 382976 261792
rect 103428 261672 103480 261724
rect 381544 261672 381596 261724
rect 91008 261604 91060 261656
rect 374644 261604 374696 261656
rect 88156 261536 88208 261588
rect 371884 261536 371936 261588
rect 110328 261468 110380 261520
rect 400864 261468 400916 261520
rect 17224 261400 17276 261452
rect 139400 261400 139452 261452
rect 161388 261400 161440 261452
rect 228824 261400 228876 261452
rect 238208 261400 238260 261452
rect 270592 261400 270644 261452
rect 22744 261332 22796 261384
rect 135352 261332 135404 261384
rect 186228 261332 186280 261384
rect 226984 261332 227036 261384
rect 240876 261332 240928 261384
rect 266360 261332 266412 261384
rect 117136 261264 117188 261316
rect 226064 261264 226116 261316
rect 104624 261196 104676 261248
rect 209044 261196 209096 261248
rect 55864 261128 55916 261180
rect 155960 261128 156012 261180
rect 117136 261060 117188 261112
rect 204904 261060 204956 261112
rect 41328 260992 41380 261044
rect 128452 260992 128504 261044
rect 121276 260924 121328 260976
rect 201500 260924 201552 260976
rect 114468 260788 114520 260840
rect 214564 260788 214616 260840
rect 101956 260720 102008 260772
rect 206376 260720 206428 260772
rect 121368 260652 121420 260704
rect 226156 260652 226208 260704
rect 25504 260584 25556 260636
rect 138112 260584 138164 260636
rect 166908 260584 166960 260636
rect 228916 260584 228968 260636
rect 15844 260516 15896 260568
rect 131120 260516 131172 260568
rect 200028 260516 200080 260568
rect 282184 260516 282236 260568
rect 4804 260448 4856 260500
rect 131212 260448 131264 260500
rect 218612 260448 218664 260500
rect 304264 260448 304316 260500
rect 89628 260380 89680 260432
rect 225236 260380 225288 260432
rect 231308 260380 231360 260432
rect 320180 260380 320232 260432
rect 93768 260312 93820 260364
rect 360844 260312 360896 260364
rect 96528 260244 96580 260296
rect 363604 260244 363656 260296
rect 56140 260176 56192 260228
rect 89720 260176 89772 260228
rect 90916 260176 90968 260228
rect 358084 260176 358136 260228
rect 53288 260108 53340 260160
rect 358912 260108 358964 260160
rect 118424 260040 118476 260092
rect 206284 260040 206336 260092
rect 282000 245556 282052 245608
rect 580172 245556 580224 245608
rect 54576 225360 54628 225412
rect 57244 225360 57296 225412
rect 2780 215228 2832 215280
rect 4804 215228 4856 215280
rect 54668 195916 54720 195968
rect 57520 195916 57572 195968
rect 53380 192652 53432 192704
rect 57520 192652 57572 192704
rect 3148 188980 3200 189032
rect 17224 188980 17276 189032
rect 54944 187620 54996 187672
rect 57244 187620 57296 187672
rect 54300 182792 54352 182844
rect 57520 182792 57572 182844
rect 57520 175584 57572 175636
rect 59820 175584 59872 175636
rect 57428 175176 57480 175228
rect 58900 175176 58952 175228
rect 54392 169668 54444 169720
rect 57796 169668 57848 169720
rect 3332 162936 3384 162988
rect 7564 162936 7616 162988
rect 55036 162800 55088 162852
rect 57428 162800 57480 162852
rect 54760 160012 54812 160064
rect 57796 160012 57848 160064
rect 52000 157292 52052 157344
rect 57428 157292 57480 157344
rect 52092 153824 52144 153876
rect 57428 153824 57480 153876
rect 396724 153144 396776 153196
rect 579620 153144 579672 153196
rect 54484 151716 54536 151768
rect 57428 151716 57480 151768
rect 53564 144576 53616 144628
rect 57428 144576 57480 144628
rect 53656 142060 53708 142112
rect 57796 142060 57848 142112
rect 3332 137912 3384 137964
rect 18604 137912 18656 137964
rect 57612 137436 57664 137488
rect 57796 137436 57848 137488
rect 53748 136552 53800 136604
rect 57612 136552 57664 136604
rect 55128 126896 55180 126948
rect 57612 126896 57664 126948
rect 260104 126896 260156 126948
rect 580172 126896 580224 126948
rect 53196 121388 53248 121440
rect 57612 121388 57664 121440
rect 52184 113092 52236 113144
rect 57612 113092 57664 113144
rect 3148 111732 3200 111784
rect 11704 111732 11756 111784
rect 56508 108332 56560 108384
rect 57244 108332 57296 108384
rect 53472 105544 53524 105596
rect 57612 105544 57664 105596
rect 54852 103436 54904 103488
rect 57612 103436 57664 103488
rect 54576 100648 54628 100700
rect 57612 100648 57664 100700
rect 3240 97928 3292 97980
rect 25504 97928 25556 97980
rect 52276 88272 52328 88324
rect 57612 88272 57664 88324
rect 3332 85484 3384 85536
rect 21364 85484 21416 85536
rect 53288 82764 53340 82816
rect 57244 82764 57296 82816
rect 3332 71680 3384 71732
rect 14464 71680 14516 71732
rect 52368 70320 52420 70372
rect 57612 70320 57664 70372
rect 208124 59848 208176 59900
rect 223856 59848 223908 59900
rect 225420 59848 225472 59900
rect 226064 59848 226116 59900
rect 580172 59916 580224 59968
rect 214564 59780 214616 59832
rect 218060 59712 218112 59764
rect 212448 59644 212500 59696
rect 213828 59576 213880 59628
rect 232228 59576 232280 59628
rect 224132 59508 224184 59560
rect 226064 59508 226116 59560
rect 233332 59576 233384 59628
rect 238024 59576 238076 59628
rect 240140 59848 240192 59900
rect 240692 59848 240744 59900
rect 267832 59848 267884 59900
rect 251180 59780 251232 59832
rect 245660 59576 245712 59628
rect 237380 59508 237432 59560
rect 207296 59440 207348 59492
rect 205548 59372 205600 59424
rect 212448 59372 212500 59424
rect 223948 59372 224000 59424
rect 232228 59372 232280 59424
rect 56692 59304 56744 59356
rect 212908 59304 212960 59356
rect 216956 59304 217008 59356
rect 224776 59304 224828 59356
rect 232412 59440 232464 59492
rect 236000 59440 236052 59492
rect 232504 59372 232556 59424
rect 322940 59372 322992 59424
rect 233332 59304 233384 59356
rect 56600 59236 56652 59288
rect 203800 59236 203852 59288
rect 215760 59236 215812 59288
rect 218428 59168 218480 59220
rect 221004 59236 221056 59288
rect 267740 59236 267792 59288
rect 224960 59168 225012 59220
rect 262220 59100 262272 59152
rect 223396 59032 223448 59084
rect 225236 59032 225288 59084
rect 207572 58964 207624 59016
rect 227996 58964 228048 59016
rect 208216 58896 208268 58948
rect 227904 58896 227956 58948
rect 209320 58828 209372 58880
rect 222476 58828 222528 58880
rect 223764 58828 223816 58880
rect 228088 58828 228140 58880
rect 216404 58760 216456 58812
rect 229192 58760 229244 58812
rect 216680 58692 216732 58744
rect 224224 58692 224276 58744
rect 224408 58692 224460 58744
rect 228272 58692 228324 58744
rect 211988 58624 212040 58676
rect 264244 58624 264296 58676
rect 214932 58556 214984 58608
rect 140228 58488 140280 58540
rect 140688 58488 140740 58540
rect 217784 58488 217836 58540
rect 219440 58488 219492 58540
rect 222292 58556 222344 58608
rect 258724 58556 258776 58608
rect 224868 58488 224920 58540
rect 210792 58420 210844 58472
rect 222384 58420 222436 58472
rect 222476 58420 222528 58472
rect 229100 58420 229152 58472
rect 217508 58352 217560 58404
rect 249064 58352 249116 58404
rect 212540 58284 212592 58336
rect 222292 58284 222344 58336
rect 222384 58284 222436 58336
rect 228180 58284 228232 58336
rect 205824 58216 205876 58268
rect 223764 58216 223816 58268
rect 224224 58216 224276 58268
rect 230480 58216 230532 58268
rect 214012 58148 214064 58200
rect 221832 58148 221884 58200
rect 221924 58148 221976 58200
rect 231952 58148 232004 58200
rect 59268 57944 59320 57996
rect 61292 57944 61344 57996
rect 45468 57876 45520 57928
rect 64696 57944 64748 57996
rect 41328 57808 41380 57860
rect 64880 57808 64932 57860
rect 143172 58012 143224 58064
rect 149428 58012 149480 58064
rect 35808 57740 35860 57792
rect 68468 57740 68520 57792
rect 39948 57672 40000 57724
rect 61936 57672 61988 57724
rect 34428 57604 34480 57656
rect 62028 57604 62080 57656
rect 33048 57536 33100 57588
rect 67916 57672 67968 57724
rect 84568 57876 84620 57928
rect 92848 57876 92900 57928
rect 95056 57876 95108 57928
rect 102140 57944 102192 57996
rect 120356 57944 120408 57996
rect 128176 57944 128228 57996
rect 132868 57944 132920 57996
rect 140964 57944 141016 57996
rect 143264 57944 143316 57996
rect 143448 57944 143500 57996
rect 162216 58080 162268 58132
rect 172152 58080 172204 58132
rect 179236 58080 179288 58132
rect 204996 58080 205048 58132
rect 100576 57876 100628 57928
rect 159824 57876 159876 57928
rect 165804 57876 165856 57928
rect 165896 57876 165948 57928
rect 168564 57876 168616 57928
rect 219532 58080 219584 58132
rect 230572 58080 230624 58132
rect 219808 58012 219860 58064
rect 231860 58012 231912 58064
rect 225052 57944 225104 57996
rect 85396 57808 85448 57860
rect 70860 57740 70912 57792
rect 80428 57740 80480 57792
rect 83004 57740 83056 57792
rect 83740 57740 83792 57792
rect 83924 57740 83976 57792
rect 86316 57740 86368 57792
rect 62212 57604 62264 57656
rect 68192 57604 68244 57656
rect 73068 57672 73120 57724
rect 77852 57672 77904 57724
rect 81900 57672 81952 57724
rect 87604 57672 87656 57724
rect 73712 57604 73764 57656
rect 74724 57604 74776 57656
rect 75276 57604 75328 57656
rect 76656 57604 76708 57656
rect 78404 57604 78456 57656
rect 81072 57604 81124 57656
rect 81348 57604 81400 57656
rect 86592 57604 86644 57656
rect 86868 57604 86920 57656
rect 87420 57604 87472 57656
rect 88156 57604 88208 57656
rect 88616 57604 88668 57656
rect 89352 57604 89404 57656
rect 91284 57604 91336 57656
rect 92296 57604 92348 57656
rect 28908 57468 28960 57520
rect 66720 57536 66772 57588
rect 66904 57536 66956 57588
rect 70216 57536 70268 57588
rect 71688 57536 71740 57588
rect 77576 57536 77628 57588
rect 80152 57536 80204 57588
rect 81256 57536 81308 57588
rect 83372 57536 83424 57588
rect 84108 57536 84160 57588
rect 86040 57536 86092 57588
rect 86684 57536 86736 57588
rect 88340 57536 88392 57588
rect 89628 57536 89680 57588
rect 64880 57468 64932 57520
rect 26148 57400 26200 57452
rect 65984 57400 66036 57452
rect 66168 57468 66220 57520
rect 76104 57468 76156 57520
rect 69940 57400 69992 57452
rect 70216 57400 70268 57452
rect 77300 57468 77352 57520
rect 80796 57468 80848 57520
rect 81348 57468 81400 57520
rect 82820 57468 82872 57520
rect 83924 57468 83976 57520
rect 84292 57468 84344 57520
rect 85396 57468 85448 57520
rect 85672 57468 85724 57520
rect 86592 57468 86644 57520
rect 92756 57604 92808 57656
rect 93676 57604 93728 57656
rect 94136 57808 94188 57860
rect 96712 57808 96764 57860
rect 96804 57808 96856 57860
rect 143172 57808 143224 57860
rect 143264 57808 143316 57860
rect 148324 57808 148376 57860
rect 149244 57808 149296 57860
rect 156788 57808 156840 57860
rect 156880 57808 156932 57860
rect 157156 57808 157208 57860
rect 159180 57808 159232 57860
rect 166816 57808 166868 57860
rect 167000 57808 167052 57860
rect 168288 57808 168340 57860
rect 168840 57808 168892 57860
rect 169576 57808 169628 57860
rect 213184 57876 213236 57928
rect 216036 57876 216088 57928
rect 173716 57808 173768 57860
rect 175556 57808 175608 57860
rect 183008 57808 183060 57860
rect 183100 57808 183152 57860
rect 183376 57808 183428 57860
rect 185124 57808 185176 57860
rect 186044 57808 186096 57860
rect 186780 57808 186832 57860
rect 187516 57808 187568 57860
rect 188068 57808 188120 57860
rect 188896 57808 188948 57860
rect 189540 57808 189592 57860
rect 190276 57808 190328 57860
rect 191288 57808 191340 57860
rect 191564 57808 191616 57860
rect 192208 57808 192260 57860
rect 193036 57808 193088 57860
rect 193220 57808 193272 57860
rect 193864 57808 193916 57860
rect 195060 57808 195112 57860
rect 195888 57808 195940 57860
rect 196256 57808 196308 57860
rect 196992 57808 197044 57860
rect 197360 57808 197412 57860
rect 198280 57808 198332 57860
rect 198832 57808 198884 57860
rect 199844 57808 199896 57860
rect 201776 57808 201828 57860
rect 202512 57808 202564 57860
rect 202972 57808 203024 57860
rect 204168 57808 204220 57860
rect 208492 57808 208544 57860
rect 218060 57808 218112 57860
rect 95884 57740 95936 57792
rect 92848 57536 92900 57588
rect 94504 57536 94556 57588
rect 95608 57604 95660 57656
rect 96344 57604 96396 57656
rect 101496 57740 101548 57792
rect 162032 57740 162084 57792
rect 162216 57740 162268 57792
rect 164516 57740 164568 57792
rect 165896 57740 165948 57792
rect 166908 57740 166960 57792
rect 167092 57740 167144 57792
rect 168104 57740 168156 57792
rect 169392 57740 169444 57792
rect 169668 57740 169720 57792
rect 169852 57740 169904 57792
rect 170864 57740 170916 57792
rect 174176 57740 174228 57792
rect 101588 57672 101640 57724
rect 101772 57672 101824 57724
rect 102048 57672 102100 57724
rect 102324 57672 102376 57724
rect 171048 57672 171100 57724
rect 171140 57672 171192 57724
rect 172152 57672 172204 57724
rect 172888 57672 172940 57724
rect 173624 57672 173676 57724
rect 174084 57672 174136 57724
rect 175004 57672 175056 57724
rect 176660 57672 176712 57724
rect 177488 57672 177540 57724
rect 178132 57672 178184 57724
rect 179052 57672 179104 57724
rect 179236 57740 179288 57792
rect 200488 57740 200540 57792
rect 200580 57740 200632 57792
rect 201224 57740 201276 57792
rect 201684 57740 201736 57792
rect 202328 57740 202380 57792
rect 203248 57740 203300 57792
rect 204076 57740 204128 57792
rect 210884 57740 210936 57792
rect 220176 57740 220228 57792
rect 221280 57876 221332 57928
rect 225788 57876 225840 57928
rect 221832 57808 221884 57860
rect 222936 57808 222988 57860
rect 223028 57808 223080 57860
rect 228364 57808 228416 57860
rect 224316 57740 224368 57792
rect 213276 57672 213328 57724
rect 213368 57672 213420 57724
rect 215116 57672 215168 57724
rect 215208 57672 215260 57724
rect 223396 57672 223448 57724
rect 97080 57604 97132 57656
rect 97264 57536 97316 57588
rect 98552 57604 98604 57656
rect 99288 57604 99340 57656
rect 100024 57604 100076 57656
rect 100576 57604 100628 57656
rect 101128 57604 101180 57656
rect 101864 57604 101916 57656
rect 103244 57604 103296 57656
rect 172704 57604 172756 57656
rect 172796 57604 172848 57656
rect 173532 57604 173584 57656
rect 174636 57604 174688 57656
rect 175188 57604 175240 57656
rect 177028 57604 177080 57656
rect 177580 57604 177632 57656
rect 177672 57604 177724 57656
rect 177948 57604 178000 57656
rect 178776 57604 178828 57656
rect 179236 57604 179288 57656
rect 179604 57604 179656 57656
rect 180432 57604 180484 57656
rect 182272 57604 182324 57656
rect 183100 57604 183152 57656
rect 183928 57604 183980 57656
rect 184848 57604 184900 57656
rect 185032 57604 185084 57656
rect 185768 57604 185820 57656
rect 188620 57604 188672 57656
rect 188988 57604 189040 57656
rect 189356 57604 189408 57656
rect 190092 57604 190144 57656
rect 190368 57604 190420 57656
rect 216036 57604 216088 57656
rect 217232 57604 217284 57656
rect 223948 57604 224000 57656
rect 103060 57536 103112 57588
rect 104348 57536 104400 57588
rect 104716 57536 104768 57588
rect 106740 57536 106792 57588
rect 107476 57536 107528 57588
rect 108212 57536 108264 57588
rect 113732 57536 113784 57588
rect 113824 57536 113876 57588
rect 142528 57536 142580 57588
rect 142620 57536 142672 57588
rect 143448 57536 143500 57588
rect 143540 57536 143592 57588
rect 77208 57400 77260 57452
rect 78680 57400 78732 57452
rect 81624 57400 81676 57452
rect 82728 57400 82780 57452
rect 83096 57400 83148 57452
rect 93124 57400 93176 57452
rect 93860 57468 93912 57520
rect 95056 57468 95108 57520
rect 95332 57468 95384 57520
rect 96436 57468 96488 57520
rect 96712 57468 96764 57520
rect 100760 57468 100812 57520
rect 100852 57468 100904 57520
rect 101956 57468 102008 57520
rect 102140 57468 102192 57520
rect 133052 57468 133104 57520
rect 133236 57468 133288 57520
rect 133696 57468 133748 57520
rect 134156 57468 134208 57520
rect 134892 57468 134944 57520
rect 135904 57468 135956 57520
rect 136364 57468 136416 57520
rect 136456 57468 136508 57520
rect 137192 57468 137244 57520
rect 138112 57468 138164 57520
rect 139124 57468 139176 57520
rect 139952 57468 140004 57520
rect 140780 57468 140832 57520
rect 141148 57468 141200 57520
rect 141976 57468 142028 57520
rect 142252 57468 142304 57520
rect 144184 57468 144236 57520
rect 144276 57468 144328 57520
rect 144828 57468 144880 57520
rect 145196 57468 145248 57520
rect 146116 57468 146168 57520
rect 146668 57536 146720 57588
rect 147496 57536 147548 57588
rect 147680 57536 147732 57588
rect 152188 57536 152240 57588
rect 152464 57536 152516 57588
rect 222936 57536 222988 57588
rect 223028 57536 223080 57588
rect 225880 57536 225932 57588
rect 147312 57468 147364 57520
rect 148048 57468 148100 57520
rect 148968 57468 149020 57520
rect 150256 57468 150308 57520
rect 214564 57468 214616 57520
rect 215116 57468 215168 57520
rect 216772 57468 216824 57520
rect 219440 57468 219492 57520
rect 226156 57468 226208 57520
rect 101404 57400 101456 57452
rect 101588 57400 101640 57452
rect 113824 57400 113876 57452
rect 113916 57400 113968 57452
rect 118608 57400 118660 57452
rect 118792 57400 118844 57452
rect 128268 57400 128320 57452
rect 128544 57400 128596 57452
rect 129648 57400 129700 57452
rect 130752 57400 130804 57452
rect 130936 57400 130988 57452
rect 131120 57400 131172 57452
rect 132040 57400 132092 57452
rect 132776 57400 132828 57452
rect 133788 57400 133840 57452
rect 134432 57400 134484 57452
rect 134984 57400 135036 57452
rect 135628 57400 135680 57452
rect 136548 57400 136600 57452
rect 136732 57400 136784 57452
rect 137836 57400 137888 57452
rect 139400 57400 139452 57452
rect 140596 57400 140648 57452
rect 140964 57400 141016 57452
rect 222384 57400 222436 57452
rect 27528 57332 27580 57384
rect 66444 57332 66496 57384
rect 67548 57332 67600 57384
rect 76380 57332 76432 57384
rect 87144 57332 87196 57384
rect 93952 57332 94004 57384
rect 94596 57332 94648 57384
rect 103612 57332 103664 57384
rect 103796 57332 103848 57384
rect 104532 57332 104584 57384
rect 105820 57332 105872 57384
rect 117320 57332 117372 57384
rect 118976 57332 119028 57384
rect 201776 57332 201828 57384
rect 202052 57332 202104 57384
rect 202788 57332 202840 57384
rect 203984 57332 204036 57384
rect 208492 57332 208544 57384
rect 210240 57332 210292 57384
rect 214380 57332 214432 57384
rect 214472 57332 214524 57384
rect 225328 57332 225380 57384
rect 6828 57264 6880 57316
rect 59268 57264 59320 57316
rect 59452 57264 59504 57316
rect 60464 57264 60516 57316
rect 62028 57264 62080 57316
rect 75184 57264 75236 57316
rect 82176 57264 82228 57316
rect 90180 57264 90232 57316
rect 91836 57264 91888 57316
rect 118516 57264 118568 57316
rect 120448 57264 120500 57316
rect 121184 57264 121236 57316
rect 122840 57264 122892 57316
rect 123300 57264 123352 57316
rect 124404 57264 124456 57316
rect 125048 57264 125100 57316
rect 125692 57264 125744 57316
rect 126612 57264 126664 57316
rect 127072 57264 127124 57316
rect 127992 57264 128044 57316
rect 128176 57264 128228 57316
rect 129832 57264 129884 57316
rect 130016 57264 130068 57316
rect 131028 57264 131080 57316
rect 131488 57264 131540 57316
rect 132132 57264 132184 57316
rect 132500 57264 132552 57316
rect 223028 57264 223080 57316
rect 24768 57196 24820 57248
rect 65892 57196 65944 57248
rect 68928 57196 68980 57248
rect 76472 57196 76524 57248
rect 83740 57196 83792 57248
rect 96712 57196 96764 57248
rect 43444 57128 43496 57180
rect 61844 57128 61896 57180
rect 61936 57128 61988 57180
rect 64880 57128 64932 57180
rect 65248 57128 65300 57180
rect 46848 57060 46900 57112
rect 68652 57128 68704 57180
rect 74080 57128 74132 57180
rect 89812 57128 89864 57180
rect 104164 57196 104216 57248
rect 104992 57196 105044 57248
rect 108212 57196 108264 57248
rect 108304 57196 108356 57248
rect 147680 57196 147732 57248
rect 147956 57196 148008 57248
rect 151820 57196 151872 57248
rect 155408 57196 155460 57248
rect 166448 57196 166500 57248
rect 166816 57196 166868 57248
rect 401600 57196 401652 57248
rect 103520 57128 103572 57180
rect 143264 57128 143316 57180
rect 143540 57128 143592 57180
rect 144644 57128 144696 57180
rect 144828 57128 144880 57180
rect 146300 57128 146352 57180
rect 146392 57128 146444 57180
rect 152464 57128 152516 57180
rect 49608 56992 49660 57044
rect 63776 56992 63828 57044
rect 74356 57060 74408 57112
rect 96160 57060 96212 57112
rect 96528 57060 96580 57112
rect 98276 57060 98328 57112
rect 99012 57060 99064 57112
rect 99104 57060 99156 57112
rect 48228 56924 48280 56976
rect 71412 56992 71464 57044
rect 79876 56992 79928 57044
rect 80428 56992 80480 57044
rect 88892 56992 88944 57044
rect 102876 56992 102928 57044
rect 71504 56924 71556 56976
rect 74816 56924 74868 56976
rect 75000 56924 75052 56976
rect 93952 56924 94004 56976
rect 102784 56924 102836 56976
rect 103704 57060 103756 57112
rect 104808 57060 104860 57112
rect 105176 57060 105228 57112
rect 156144 57128 156196 57180
rect 153660 57060 153712 57112
rect 154488 57060 154540 57112
rect 156328 57060 156380 57112
rect 210884 57128 210936 57180
rect 212264 57128 212316 57180
rect 162032 57060 162084 57112
rect 168564 57060 168616 57112
rect 168656 57060 168708 57112
rect 213368 57060 213420 57112
rect 213736 57128 213788 57180
rect 215392 57060 215444 57112
rect 215484 57060 215536 57112
rect 216588 57060 216640 57112
rect 216772 57128 216824 57180
rect 222016 57060 222068 57112
rect 222200 57128 222252 57180
rect 300124 57128 300176 57180
rect 224132 57060 224184 57112
rect 103060 56992 103112 57044
rect 132684 56992 132736 57044
rect 132868 56992 132920 57044
rect 142160 56992 142212 57044
rect 142252 56992 142304 57044
rect 133788 56924 133840 56976
rect 53748 56856 53800 56908
rect 65156 56856 65208 56908
rect 65524 56856 65576 56908
rect 71780 56856 71832 56908
rect 76564 56856 76616 56908
rect 78128 56856 78180 56908
rect 93308 56856 93360 56908
rect 135444 56924 135496 56976
rect 137008 56924 137060 56976
rect 141332 56924 141384 56976
rect 141424 56924 141476 56976
rect 146944 56924 146996 56976
rect 147312 56924 147364 56976
rect 150256 56924 150308 56976
rect 150440 56924 150492 56976
rect 151544 56924 151596 56976
rect 151912 56924 151964 56976
rect 153108 56924 153160 56976
rect 153384 56924 153436 56976
rect 154212 56924 154264 56976
rect 154580 56924 154632 56976
rect 155868 56924 155920 56976
rect 155960 56924 156012 56976
rect 157064 56924 157116 56976
rect 161572 56992 161624 57044
rect 166356 56992 166408 57044
rect 166908 56992 166960 57044
rect 162768 56924 162820 56976
rect 163320 56924 163372 56976
rect 166816 56924 166868 56976
rect 167184 56924 167236 56976
rect 213552 56924 213604 56976
rect 214564 56992 214616 57044
rect 220268 56992 220320 57044
rect 220728 56992 220780 57044
rect 302240 56992 302292 57044
rect 215944 56924 215996 56976
rect 216588 56924 216640 56976
rect 277492 56924 277544 56976
rect 133972 56856 134024 56908
rect 134708 56856 134760 56908
rect 134800 56856 134852 56908
rect 138664 56856 138716 56908
rect 138756 56856 138808 56908
rect 142068 56856 142120 56908
rect 53656 56788 53708 56840
rect 63408 56788 63460 56840
rect 65616 56788 65668 56840
rect 72884 56788 72936 56840
rect 89168 56788 89220 56840
rect 89536 56788 89588 56840
rect 90732 56788 90784 56840
rect 91008 56788 91060 56840
rect 91560 56788 91612 56840
rect 94596 56788 94648 56840
rect 94688 56788 94740 56840
rect 99104 56788 99156 56840
rect 99748 56788 99800 56840
rect 105176 56788 105228 56840
rect 105268 56788 105320 56840
rect 106188 56788 106240 56840
rect 107844 56788 107896 56840
rect 108764 56788 108816 56840
rect 110236 56788 110288 56840
rect 113640 56788 113692 56840
rect 113732 56788 113784 56840
rect 132500 56788 132552 56840
rect 132684 56788 132736 56840
rect 142528 56856 142580 56908
rect 144920 56856 144972 56908
rect 145104 56856 145156 56908
rect 146576 56788 146628 56840
rect 146668 56788 146720 56840
rect 156052 56788 156104 56840
rect 180892 56856 180944 56908
rect 180984 56856 181036 56908
rect 181904 56856 181956 56908
rect 182548 56856 182600 56908
rect 183284 56856 183336 56908
rect 186320 56856 186372 56908
rect 187240 56856 187292 56908
rect 190736 56856 190788 56908
rect 191656 56856 191708 56908
rect 191840 56856 191892 56908
rect 193036 56856 193088 56908
rect 193588 56856 193640 56908
rect 194232 56856 194284 56908
rect 194600 56856 194652 56908
rect 195704 56856 195756 56908
rect 198280 56856 198332 56908
rect 198556 56856 198608 56908
rect 198740 56856 198792 56908
rect 200028 56856 200080 56908
rect 201776 56856 201828 56908
rect 203524 56856 203576 56908
rect 204720 56856 204772 56908
rect 55128 56720 55180 56772
rect 64788 56720 64840 56772
rect 65340 56720 65392 56772
rect 73160 56720 73212 56772
rect 84844 56720 84896 56772
rect 86224 56720 86276 56772
rect 98828 56720 98880 56772
rect 99196 56720 99248 56772
rect 99380 56720 99432 56772
rect 100668 56720 100720 56772
rect 100760 56720 100812 56772
rect 103060 56720 103112 56772
rect 103612 56720 103664 56772
rect 105544 56720 105596 56772
rect 106372 56720 106424 56772
rect 107568 56720 107620 56772
rect 107660 56720 107712 56772
rect 108488 56720 108540 56772
rect 59268 56652 59320 56704
rect 57244 56584 57296 56636
rect 64696 56584 64748 56636
rect 65248 56584 65300 56636
rect 64880 56516 64932 56568
rect 69664 56652 69716 56704
rect 70308 56652 70360 56704
rect 76932 56652 76984 56704
rect 90088 56652 90140 56704
rect 91008 56652 91060 56704
rect 98000 56652 98052 56704
rect 99104 56652 99156 56704
rect 102600 56652 102652 56704
rect 103336 56652 103388 56704
rect 104072 56652 104124 56704
rect 64788 56448 64840 56500
rect 73436 56584 73488 56636
rect 97632 56584 97684 56636
rect 108304 56584 108356 56636
rect 113916 56720 113968 56772
rect 114100 56720 114152 56772
rect 118608 56720 118660 56772
rect 118700 56720 118752 56772
rect 119804 56720 119856 56772
rect 120080 56720 120132 56772
rect 120724 56720 120776 56772
rect 123300 56720 123352 56772
rect 123944 56720 123996 56772
rect 124588 56720 124640 56772
rect 125416 56720 125468 56772
rect 125600 56720 125652 56772
rect 126244 56720 126296 56772
rect 126336 56720 126388 56772
rect 129740 56720 129792 56772
rect 129832 56720 129884 56772
rect 130384 56720 130436 56772
rect 131212 56720 131264 56772
rect 132408 56720 132460 56772
rect 133788 56720 133840 56772
rect 136732 56720 136784 56772
rect 136824 56720 136876 56772
rect 138020 56720 138072 56772
rect 138480 56720 138532 56772
rect 139124 56720 139176 56772
rect 139216 56720 139268 56772
rect 142068 56720 142120 56772
rect 110788 56652 110840 56704
rect 109316 56584 109368 56636
rect 110328 56584 110380 56636
rect 110512 56584 110564 56636
rect 111616 56584 111668 56636
rect 112260 56584 112312 56636
rect 112996 56584 113048 56636
rect 113456 56652 113508 56704
rect 114376 56652 114428 56704
rect 115204 56652 115256 56704
rect 115756 56652 115808 56704
rect 116032 56652 116084 56704
rect 117136 56652 117188 56704
rect 146852 56720 146904 56772
rect 146944 56720 146996 56772
rect 162952 56720 163004 56772
rect 164056 56720 164108 56772
rect 165620 56720 165672 56772
rect 166724 56720 166776 56772
rect 166816 56720 166868 56772
rect 167184 56720 167236 56772
rect 168380 56720 168432 56772
rect 169116 56720 169168 56772
rect 170312 56720 170364 56772
rect 171048 56720 171100 56772
rect 171416 56720 171468 56772
rect 172336 56720 172388 56772
rect 172704 56788 172756 56840
rect 174912 56788 174964 56840
rect 175280 56788 175332 56840
rect 176384 56788 176436 56840
rect 175740 56720 175792 56772
rect 175832 56720 175884 56772
rect 176568 56720 176620 56772
rect 114192 56584 114244 56636
rect 114468 56584 114520 56636
rect 114836 56584 114888 56636
rect 115572 56584 115624 56636
rect 116860 56584 116912 56636
rect 116952 56584 117004 56636
rect 117228 56584 117280 56636
rect 113640 56448 113692 56500
rect 142252 56652 142304 56704
rect 147772 56652 147824 56704
rect 147864 56652 147916 56704
rect 148784 56652 148836 56704
rect 149612 56652 149664 56704
rect 150256 56652 150308 56704
rect 151084 56652 151136 56704
rect 151636 56652 151688 56704
rect 152832 56652 152884 56704
rect 153016 56652 153068 56704
rect 153936 56652 153988 56704
rect 154396 56652 154448 56704
rect 154856 56652 154908 56704
rect 155776 56652 155828 56704
rect 156788 56652 156840 56704
rect 170404 56652 170456 56704
rect 173716 56652 173768 56704
rect 204812 56788 204864 56840
rect 205272 56856 205324 56908
rect 213828 56856 213880 56908
rect 214748 56856 214800 56908
rect 229468 56856 229520 56908
rect 209872 56788 209924 56840
rect 213460 56788 213512 56840
rect 176752 56720 176804 56772
rect 180708 56720 180760 56772
rect 180892 56720 180944 56772
rect 182916 56720 182968 56772
rect 183008 56720 183060 56772
rect 190368 56720 190420 56772
rect 193312 56720 193364 56772
rect 194416 56720 194468 56772
rect 197728 56720 197780 56772
rect 198556 56720 198608 56772
rect 200488 56720 200540 56772
rect 179880 56652 179932 56704
rect 180524 56652 180576 56704
rect 180800 56652 180852 56704
rect 204720 56652 204772 56704
rect 206468 56720 206520 56772
rect 214472 56720 214524 56772
rect 214656 56720 214708 56772
rect 216312 56720 216364 56772
rect 216496 56788 216548 56840
rect 221924 56788 221976 56840
rect 222016 56788 222068 56840
rect 226248 56788 226300 56840
rect 225696 56720 225748 56772
rect 208400 56652 208452 56704
rect 208492 56652 208544 56704
rect 214748 56652 214800 56704
rect 215392 56652 215444 56704
rect 221832 56652 221884 56704
rect 221924 56652 221976 56704
rect 225972 56652 226024 56704
rect 117320 56380 117372 56432
rect 142160 56584 142212 56636
rect 118516 56516 118568 56568
rect 120724 56516 120776 56568
rect 128268 56516 128320 56568
rect 129832 56516 129884 56568
rect 139860 56448 139912 56500
rect 156696 56584 156748 56636
rect 158076 56584 158128 56636
rect 158628 56584 158680 56636
rect 158904 56584 158956 56636
rect 160008 56584 160060 56636
rect 160928 56584 160980 56636
rect 161388 56584 161440 56636
rect 162124 56584 162176 56636
rect 162676 56584 162728 56636
rect 162768 56584 162820 56636
rect 163872 56584 163924 56636
rect 164148 56584 164200 56636
rect 164608 56584 164660 56636
rect 164700 56584 164752 56636
rect 165436 56584 165488 56636
rect 166540 56584 166592 56636
rect 166816 56584 166868 56636
rect 166448 56516 166500 56568
rect 219624 56584 219676 56636
rect 219900 56584 219952 56636
rect 276664 56584 276716 56636
rect 174912 56516 174964 56568
rect 175280 56516 175332 56568
rect 182916 56516 182968 56568
rect 184204 56516 184256 56568
rect 184388 56516 184440 56568
rect 450544 56516 450596 56568
rect 180248 56448 180300 56500
rect 447784 56448 447836 56500
rect 142068 56380 142120 56432
rect 142620 56380 142672 56432
rect 175740 56380 175792 56432
rect 178132 56380 178184 56432
rect 182088 56380 182140 56432
rect 454684 56380 454736 56432
rect 182824 56312 182876 56364
rect 461584 56312 461636 56364
rect 178408 56244 178460 56296
rect 479524 56244 479576 56296
rect 74816 56176 74868 56228
rect 75644 56176 75696 56228
rect 181076 56176 181128 56228
rect 184388 56176 184440 56228
rect 184572 56176 184624 56228
rect 468484 56176 468536 56228
rect 179328 56108 179380 56160
rect 483020 56108 483072 56160
rect 183744 56040 183796 56092
rect 500960 56040 501012 56092
rect 185492 55972 185544 56024
rect 507860 55972 507912 56024
rect 129740 55904 129792 55956
rect 178040 55904 178092 55956
rect 189264 55904 189316 55956
rect 519544 55904 519596 55956
rect 55772 55836 55824 55888
rect 580356 55836 580408 55888
rect 112812 55768 112864 55820
rect 167368 55768 167420 55820
rect 434720 55768 434772 55820
rect 63500 55564 63552 55616
rect 64236 55564 64288 55616
rect 63684 55496 63736 55548
rect 64512 55496 64564 55548
rect 127900 55700 127952 55752
rect 128176 55700 128228 55752
rect 152372 55700 152424 55752
rect 152832 55700 152884 55752
rect 163596 55700 163648 55752
rect 417424 55700 417476 55752
rect 116308 55632 116360 55684
rect 227720 55632 227772 55684
rect 114560 55564 114612 55616
rect 220820 55564 220872 55616
rect 213920 55496 213972 55548
rect 111064 55428 111116 55480
rect 207020 55428 207072 55480
rect 111984 55360 112036 55412
rect 209780 55360 209832 55412
rect 112720 55292 112772 55344
rect 112904 55292 112956 55344
rect 158260 55292 158312 55344
rect 158536 55292 158588 55344
rect 137100 55156 137152 55208
rect 313280 55156 313332 55208
rect 138296 55088 138348 55140
rect 316040 55088 316092 55140
rect 138112 55020 138164 55072
rect 320180 55020 320232 55072
rect 140780 54952 140832 55004
rect 324320 54952 324372 55004
rect 140872 54884 140924 54936
rect 327080 54884 327132 54936
rect 157616 54816 157668 54868
rect 158536 54816 158588 54868
rect 160100 54816 160152 54868
rect 405740 54816 405792 54868
rect 161848 54748 161900 54800
rect 412640 54748 412692 54800
rect 166172 54680 166224 54732
rect 430580 54680 430632 54732
rect 60648 54612 60700 54664
rect 75000 54612 75052 54664
rect 167000 54612 167052 54664
rect 438860 54612 438912 54664
rect 50988 54544 51040 54596
rect 71872 54544 71924 54596
rect 185032 54544 185084 54596
rect 475384 54544 475436 54596
rect 38568 54476 38620 54528
rect 69388 54476 69440 54528
rect 189356 54476 189408 54528
rect 526444 54476 526496 54528
rect 137192 54408 137244 54460
rect 309140 54408 309192 54460
rect 133972 54340 134024 54392
rect 302240 54340 302292 54392
rect 131120 54272 131172 54324
rect 132316 54272 132368 54324
rect 132776 54272 132828 54324
rect 299480 54272 299532 54324
rect 129740 54204 129792 54256
rect 218060 54204 218112 54256
rect 161388 53728 161440 53780
rect 407764 53728 407816 53780
rect 162584 53660 162636 53712
rect 414664 53660 414716 53712
rect 164424 53592 164476 53644
rect 421564 53592 421616 53644
rect 186780 53524 186832 53576
rect 443644 53524 443696 53576
rect 165344 53456 165396 53508
rect 425704 53456 425756 53508
rect 171508 53388 171560 53440
rect 452660 53388 452712 53440
rect 183928 53320 183980 53372
rect 472624 53320 472676 53372
rect 183836 53252 183888 53304
rect 502340 53252 502392 53304
rect 186596 53184 186648 53236
rect 512644 53184 512696 53236
rect 188160 53116 188212 53168
rect 520280 53116 520332 53168
rect 190828 53048 190880 53100
rect 530584 53048 530636 53100
rect 119252 52980 119304 53032
rect 240140 52980 240192 53032
rect 116584 52912 116636 52964
rect 229100 52912 229152 52964
rect 115848 52844 115900 52896
rect 226340 52844 226392 52896
rect 123484 52776 123536 52828
rect 233240 52776 233292 52828
rect 142896 52708 142948 52760
rect 236000 52708 236052 52760
rect 156144 52640 156196 52692
rect 160192 52640 160244 52692
rect 121920 52368 121972 52420
rect 251180 52368 251232 52420
rect 122748 52300 122800 52352
rect 253940 52300 253992 52352
rect 142804 52232 142856 52284
rect 335360 52232 335412 52284
rect 143724 52164 143776 52216
rect 339500 52164 339552 52216
rect 143540 52096 143592 52148
rect 342260 52096 342312 52148
rect 145472 52028 145524 52080
rect 346400 52028 346452 52080
rect 148140 51960 148192 52012
rect 357532 51960 357584 52012
rect 149888 51892 149940 51944
rect 364340 51892 364392 51944
rect 168380 51824 168432 51876
rect 436744 51824 436796 51876
rect 192116 51756 192168 51808
rect 535460 51756 535512 51808
rect 193220 51688 193272 51740
rect 542360 51688 542412 51740
rect 143908 51620 143960 51672
rect 247040 51620 247092 51672
rect 177120 51348 177172 51400
rect 177948 51348 178000 51400
rect 172796 51008 172848 51060
rect 432604 51008 432656 51060
rect 169760 50940 169812 50992
rect 445760 50940 445812 50992
rect 169852 50872 169904 50924
rect 448520 50872 448572 50924
rect 172612 50804 172664 50856
rect 456800 50804 456852 50856
rect 174268 50736 174320 50788
rect 463700 50736 463752 50788
rect 196440 50668 196492 50720
rect 533344 50668 533396 50720
rect 194600 50600 194652 50652
rect 537484 50600 537536 50652
rect 197544 50532 197596 50584
rect 544384 50532 544436 50584
rect 194692 50464 194744 50516
rect 199200 50396 199252 50448
rect 200028 50464 200080 50516
rect 539600 50464 539652 50516
rect 106372 50328 106424 50380
rect 107568 50328 107620 50380
rect 107660 50328 107712 50380
rect 108948 50328 109000 50380
rect 109040 50328 109092 50380
rect 110144 50328 110196 50380
rect 130108 50328 130160 50380
rect 130936 50328 130988 50380
rect 135260 50328 135312 50380
rect 136456 50328 136508 50380
rect 187700 50328 187752 50380
rect 188804 50328 188856 50380
rect 196072 50328 196124 50380
rect 197176 50328 197228 50380
rect 198740 50328 198792 50380
rect 199752 50328 199804 50380
rect 546500 50396 546552 50448
rect 564440 50328 564492 50380
rect 147680 50260 147732 50312
rect 360200 50260 360252 50312
rect 137928 50192 137980 50244
rect 280160 50192 280212 50244
rect 192208 50124 192260 50176
rect 200028 50124 200080 50176
rect 200120 50124 200172 50176
rect 201316 50124 201368 50176
rect 201684 50124 201736 50176
rect 202604 50124 202656 50176
rect 201592 50056 201644 50108
rect 202696 50056 202748 50108
rect 151820 49308 151872 49360
rect 291200 49308 291252 49360
rect 178132 49240 178184 49292
rect 329840 49240 329892 49292
rect 156696 49172 156748 49224
rect 322940 49172 322992 49224
rect 141332 49104 141384 49156
rect 311900 49104 311952 49156
rect 156052 49036 156104 49088
rect 340880 49036 340932 49088
rect 197360 48968 197412 49020
rect 560300 48968 560352 49020
rect 242348 46860 242400 46912
rect 579988 46860 580040 46912
rect 124404 46316 124456 46368
rect 125508 46316 125560 46368
rect 124588 46248 124640 46300
rect 125324 46248 125376 46300
rect 125784 46248 125836 46300
rect 126888 46248 126940 46300
rect 126980 46248 127032 46300
rect 128268 46248 128320 46300
rect 118884 46180 118936 46232
rect 119896 46180 119948 46232
rect 120080 46180 120132 46232
rect 121368 46180 121420 46232
rect 122840 46180 122892 46232
rect 124128 46180 124180 46232
rect 124496 46180 124548 46232
rect 125232 46180 125284 46232
rect 125600 46180 125652 46232
rect 126704 46180 126756 46232
rect 127072 46180 127124 46232
rect 128084 46180 128136 46232
rect 124312 46112 124364 46164
rect 125416 46112 125468 46164
rect 119344 45364 119396 45416
rect 119712 45364 119764 45416
rect 2872 33056 2924 33108
rect 15844 33056 15896 33108
rect 130384 24080 130436 24132
rect 242900 24080 242952 24132
rect 3424 20612 3476 20664
rect 29644 20612 29696 20664
rect 55680 20612 55732 20664
rect 580080 20612 580132 20664
rect 204904 20068 204956 20120
rect 440240 20068 440292 20120
rect 209044 20000 209096 20052
rect 454040 20000 454092 20052
rect 216036 19932 216088 19984
rect 467840 19932 467892 19984
rect 115664 18844 115716 18896
rect 224960 18844 225012 18896
rect 164884 18776 164936 18828
rect 318800 18776 318852 18828
rect 160744 18708 160796 18760
rect 325700 18708 325752 18760
rect 170404 18640 170456 18692
rect 361580 18640 361632 18692
rect 213276 18572 213328 18624
rect 460940 18572 460992 18624
rect 126520 17892 126572 17944
rect 269120 17892 269172 17944
rect 127900 17824 127952 17876
rect 273260 17824 273312 17876
rect 127992 17756 128044 17808
rect 276020 17756 276072 17808
rect 130752 17688 130804 17740
rect 287060 17688 287112 17740
rect 184204 17620 184256 17672
rect 343640 17620 343692 17672
rect 133604 17552 133656 17604
rect 298100 17552 298152 17604
rect 134984 17484 135036 17536
rect 300860 17484 300912 17536
rect 136272 17416 136324 17468
rect 307760 17416 307812 17468
rect 137744 17348 137796 17400
rect 316132 17348 316184 17400
rect 144184 17280 144236 17332
rect 332600 17280 332652 17332
rect 141884 17212 141936 17264
rect 332692 17212 332744 17264
rect 126612 17144 126664 17196
rect 266360 17144 266412 17196
rect 125140 17076 125192 17128
rect 262220 17076 262272 17128
rect 119804 16532 119856 16584
rect 238116 16532 238168 16584
rect 119712 16464 119764 16516
rect 241704 16464 241756 16516
rect 121184 16396 121236 16448
rect 245200 16396 245252 16448
rect 121276 16328 121328 16380
rect 248788 16328 248840 16380
rect 122564 16260 122616 16312
rect 252376 16260 252428 16312
rect 123852 16192 123904 16244
rect 255872 16192 255924 16244
rect 123944 16124 123996 16176
rect 259460 16124 259512 16176
rect 199752 16056 199804 16108
rect 568028 16056 568080 16108
rect 201132 15988 201184 16040
rect 571524 15988 571576 16040
rect 202512 15920 202564 15972
rect 575112 15920 575164 15972
rect 90732 15852 90784 15904
rect 123576 15852 123628 15904
rect 202420 15852 202472 15904
rect 578608 15852 578660 15904
rect 118516 15784 118568 15836
rect 234620 15784 234672 15836
rect 117044 15716 117096 15768
rect 231032 15716 231084 15768
rect 117136 15648 117188 15700
rect 227536 15648 227588 15700
rect 115756 15580 115808 15632
rect 223948 15580 224000 15632
rect 114284 15512 114336 15564
rect 219992 15512 220044 15564
rect 114376 15444 114428 15496
rect 216864 15444 216916 15496
rect 112904 15376 112956 15428
rect 213092 15376 213144 15428
rect 111524 15308 111576 15360
rect 209872 15308 209924 15360
rect 183284 15104 183336 15156
rect 497096 15104 497148 15156
rect 183192 15036 183244 15088
rect 500592 15036 500644 15088
rect 184572 14968 184624 15020
rect 504180 14968 504232 15020
rect 186044 14900 186096 14952
rect 507676 14900 507728 14952
rect 186136 14832 186188 14884
rect 511264 14832 511316 14884
rect 187424 14764 187476 14816
rect 514760 14764 514812 14816
rect 188804 14696 188856 14748
rect 518348 14696 518400 14748
rect 188712 14628 188764 14680
rect 521844 14628 521896 14680
rect 190276 14560 190328 14612
rect 525432 14560 525484 14612
rect 190184 14492 190236 14544
rect 529020 14492 529072 14544
rect 191564 14424 191616 14476
rect 532516 14424 532568 14476
rect 181996 14356 182048 14408
rect 493508 14356 493560 14408
rect 181904 14288 181956 14340
rect 489920 14288 489972 14340
rect 180524 14220 180576 14272
rect 486424 14220 486476 14272
rect 179144 14152 179196 14204
rect 481640 14152 481692 14204
rect 177672 14084 177724 14136
rect 478144 14084 478196 14136
rect 177580 14016 177632 14068
rect 473360 14016 473412 14068
rect 176476 13948 176528 14000
rect 471060 13948 471112 14000
rect 176384 13880 176436 13932
rect 467472 13880 467524 13932
rect 158352 13744 158404 13796
rect 396540 13744 396592 13796
rect 158260 13676 158312 13728
rect 398840 13676 398892 13728
rect 159916 13608 159968 13660
rect 403624 13608 403676 13660
rect 161020 13540 161072 13592
rect 407212 13540 407264 13592
rect 161204 13472 161256 13524
rect 410800 13472 410852 13524
rect 162676 13404 162728 13456
rect 414296 13404 414348 13456
rect 164056 13336 164108 13388
rect 417424 13336 417476 13388
rect 163964 13268 164016 13320
rect 421380 13268 421432 13320
rect 165436 13200 165488 13252
rect 423772 13200 423824 13252
rect 166724 13132 166776 13184
rect 428464 13132 428516 13184
rect 166816 13064 166868 13116
rect 432052 13064 432104 13116
rect 156972 12996 157024 13048
rect 393044 12996 393096 13048
rect 157064 12928 157116 12980
rect 389456 12928 389508 12980
rect 155592 12860 155644 12912
rect 385960 12860 386012 12912
rect 154304 12792 154356 12844
rect 382372 12792 382424 12844
rect 154212 12724 154264 12776
rect 378876 12724 378928 12776
rect 152740 12656 152792 12708
rect 374000 12656 374052 12708
rect 151360 12588 151412 12640
rect 368204 12588 368256 12640
rect 132224 12384 132276 12436
rect 293684 12384 293736 12436
rect 133696 12316 133748 12368
rect 297272 12316 297324 12368
rect 134892 12248 134944 12300
rect 299572 12248 299624 12300
rect 135076 12180 135128 12232
rect 304356 12180 304408 12232
rect 136364 12112 136416 12164
rect 307944 12112 307996 12164
rect 137836 12044 137888 12096
rect 311440 12044 311492 12096
rect 137652 11976 137704 12028
rect 315028 11976 315080 12028
rect 139124 11908 139176 11960
rect 318524 11908 318576 11960
rect 140596 11840 140648 11892
rect 322112 11840 322164 11892
rect 140688 11772 140740 11824
rect 325608 11772 325660 11824
rect 141976 11704 142028 11756
rect 329196 11704 329248 11756
rect 132132 11636 132184 11688
rect 290188 11636 290240 11688
rect 130844 11568 130896 11620
rect 286600 11568 286652 11620
rect 129464 11500 129516 11552
rect 279516 11500 279568 11552
rect 128084 11432 128136 11484
rect 276112 11432 276164 11484
rect 126704 11364 126756 11416
rect 268844 11364 268896 11416
rect 125324 11296 125376 11348
rect 265348 11296 265400 11348
rect 125232 11228 125284 11280
rect 261760 11228 261812 11280
rect 124036 11160 124088 11212
rect 258264 11160 258316 11212
rect 209780 11092 209832 11144
rect 210976 11092 211028 11144
rect 194232 10956 194284 11008
rect 541992 10956 542044 11008
rect 106004 10888 106056 10940
rect 184940 10888 184992 10940
rect 194324 10888 194376 10940
rect 545488 10888 545540 10940
rect 107200 10820 107252 10872
rect 188528 10820 188580 10872
rect 195796 10820 195848 10872
rect 547880 10820 547932 10872
rect 107292 10752 107344 10804
rect 190828 10752 190880 10804
rect 196992 10752 197044 10804
rect 552664 10752 552716 10804
rect 107384 10684 107436 10736
rect 192024 10684 192076 10736
rect 197084 10684 197136 10736
rect 556160 10684 556212 10736
rect 108764 10616 108816 10668
rect 193220 10616 193272 10668
rect 198464 10616 198516 10668
rect 559748 10616 559800 10668
rect 108672 10548 108724 10600
rect 195612 10548 195664 10600
rect 199844 10548 199896 10600
rect 563244 10548 563296 10600
rect 108856 10480 108908 10532
rect 197912 10480 197964 10532
rect 199936 10480 199988 10532
rect 566832 10480 566884 10532
rect 110144 10412 110196 10464
rect 199108 10412 199160 10464
rect 201224 10412 201276 10464
rect 570328 10412 570380 10464
rect 110236 10344 110288 10396
rect 202696 10344 202748 10396
rect 202880 10344 202932 10396
rect 572720 10344 572772 10396
rect 110052 10276 110104 10328
rect 201592 10276 201644 10328
rect 202512 10276 202564 10328
rect 577412 10276 577464 10328
rect 192944 10208 192996 10260
rect 538404 10208 538456 10260
rect 193036 10140 193088 10192
rect 534908 10140 534960 10192
rect 115572 10072 115624 10124
rect 222752 10072 222804 10124
rect 114468 10004 114520 10056
rect 219256 10004 219308 10056
rect 112812 9936 112864 9988
rect 215668 9936 215720 9988
rect 112996 9868 113048 9920
rect 212172 9868 212224 9920
rect 111432 9800 111484 9852
rect 208584 9800 208636 9852
rect 111616 9732 111668 9784
rect 205088 9732 205140 9784
rect 175096 9596 175148 9648
rect 466276 9596 466328 9648
rect 176568 9528 176620 9580
rect 469864 9528 469916 9580
rect 177764 9460 177816 9512
rect 473452 9460 473504 9512
rect 177948 9392 178000 9444
rect 475752 9392 475804 9444
rect 98920 9324 98972 9376
rect 158904 9324 158956 9376
rect 177856 9324 177908 9376
rect 476948 9324 477000 9376
rect 100484 9256 100536 9308
rect 163688 9256 163740 9308
rect 179236 9256 179288 9308
rect 481732 9256 481784 9308
rect 101864 9188 101916 9240
rect 167184 9188 167236 9240
rect 180432 9188 180484 9240
rect 485228 9188 485280 9240
rect 101772 9120 101824 9172
rect 170772 9120 170824 9172
rect 180616 9120 180668 9172
rect 488816 9120 488868 9172
rect 103336 9052 103388 9104
rect 174268 9052 174320 9104
rect 181812 9052 181864 9104
rect 492312 9052 492364 9104
rect 86224 8984 86276 9036
rect 101036 8984 101088 9036
rect 104440 8984 104492 9036
rect 177856 8984 177908 9036
rect 183100 8984 183152 9036
rect 495900 8984 495952 9036
rect 86592 8916 86644 8968
rect 104532 8916 104584 8968
rect 104624 8916 104676 8968
rect 181444 8916 181496 8968
rect 183376 8916 183428 8968
rect 499396 8916 499448 8968
rect 175004 8848 175056 8900
rect 462780 8848 462832 8900
rect 173716 8780 173768 8832
rect 459192 8780 459244 8832
rect 172244 8712 172296 8764
rect 455696 8712 455748 8764
rect 172336 8644 172388 8696
rect 452108 8644 452160 8696
rect 170956 8576 171008 8628
rect 448612 8576 448664 8628
rect 169484 8508 169536 8560
rect 445024 8508 445076 8560
rect 169576 8440 169628 8492
rect 441528 8440 441580 8492
rect 168196 8372 168248 8424
rect 437940 8372 437992 8424
rect 93124 8304 93176 8356
rect 93952 8304 94004 8356
rect 168104 8304 168156 8356
rect 434444 8304 434496 8356
rect 150256 8236 150308 8288
rect 363512 8236 363564 8288
rect 151544 8168 151596 8220
rect 367008 8168 367060 8220
rect 151452 8100 151504 8152
rect 370596 8100 370648 8152
rect 152832 8032 152884 8084
rect 374092 8032 374144 8084
rect 93584 7964 93636 8016
rect 134156 7964 134208 8016
rect 152924 7964 152976 8016
rect 377680 7964 377732 8016
rect 95056 7896 95108 7948
rect 137652 7896 137704 7948
rect 154396 7896 154448 7948
rect 381176 7896 381228 7948
rect 95148 7828 95200 7880
rect 141240 7828 141292 7880
rect 155776 7828 155828 7880
rect 384764 7828 384816 7880
rect 96344 7760 96396 7812
rect 144736 7760 144788 7812
rect 155684 7760 155736 7812
rect 388260 7760 388312 7812
rect 96252 7692 96304 7744
rect 148232 7692 148284 7744
rect 157156 7692 157208 7744
rect 391848 7692 391900 7744
rect 97908 7624 97960 7676
rect 151820 7624 151872 7676
rect 158536 7624 158588 7676
rect 395344 7624 395396 7676
rect 99012 7556 99064 7608
rect 155408 7556 155460 7608
rect 158444 7556 158496 7608
rect 398932 7556 398984 7608
rect 148876 7488 148928 7540
rect 359924 7488 359976 7540
rect 148784 7420 148836 7472
rect 356336 7420 356388 7472
rect 147312 7352 147364 7404
rect 352840 7352 352892 7404
rect 146116 7284 146168 7336
rect 345756 7284 345808 7336
rect 144828 7216 144880 7268
rect 342168 7216 342220 7268
rect 143356 7148 143408 7200
rect 338672 7148 338724 7200
rect 143448 7080 143500 7132
rect 335084 7080 335136 7132
rect 141792 7012 141844 7064
rect 331588 7012 331640 7064
rect 3424 6808 3476 6860
rect 22744 6808 22796 6860
rect 125508 6808 125560 6860
rect 264152 6808 264204 6860
rect 126888 6740 126940 6792
rect 267740 6740 267792 6792
rect 126796 6672 126848 6724
rect 271236 6672 271288 6724
rect 128176 6604 128228 6656
rect 274824 6604 274876 6656
rect 129648 6536 129700 6588
rect 278320 6536 278372 6588
rect 129556 6468 129608 6520
rect 281908 6468 281960 6520
rect 130936 6400 130988 6452
rect 285404 6400 285456 6452
rect 132408 6332 132460 6384
rect 288992 6332 289044 6384
rect 132316 6264 132368 6316
rect 292580 6264 292632 6316
rect 105544 6196 105596 6248
rect 128176 6196 128228 6248
rect 133512 6196 133564 6248
rect 296076 6196 296128 6248
rect 92204 6128 92256 6180
rect 130568 6128 130620 6180
rect 151636 6128 151688 6180
rect 369400 6128 369452 6180
rect 125416 6060 125468 6112
rect 260656 6060 260708 6112
rect 124128 5992 124180 6044
rect 257068 5992 257120 6044
rect 122656 5924 122708 5976
rect 253480 5924 253532 5976
rect 122380 5856 122432 5908
rect 249984 5856 250036 5908
rect 121368 5788 121420 5840
rect 246396 5788 246448 5840
rect 119620 5720 119672 5772
rect 242992 5720 243044 5772
rect 119896 5652 119948 5704
rect 239312 5652 239364 5704
rect 118608 5584 118660 5636
rect 235816 5584 235868 5636
rect 116952 5516 117004 5568
rect 232228 5516 232280 5568
rect 276020 5516 276072 5568
rect 277124 5516 277176 5568
rect 299572 5516 299624 5568
rect 300768 5516 300820 5568
rect 101956 5448 102008 5500
rect 166080 5448 166132 5500
rect 191472 5448 191524 5500
rect 533712 5448 533764 5500
rect 102048 5380 102100 5432
rect 169576 5380 169628 5432
rect 192760 5380 192812 5432
rect 537208 5380 537260 5432
rect 103428 5312 103480 5364
rect 173164 5312 173216 5364
rect 194416 5312 194468 5364
rect 540796 5312 540848 5364
rect 104808 5244 104860 5296
rect 176660 5244 176712 5296
rect 196900 5244 196952 5296
rect 204904 5244 204956 5296
rect 204996 5244 205048 5296
rect 544292 5244 544344 5296
rect 104716 5176 104768 5228
rect 180248 5176 180300 5228
rect 195888 5176 195940 5228
rect 547972 5176 548024 5228
rect 106188 5108 106240 5160
rect 183744 5108 183796 5160
rect 187240 5108 187292 5160
rect 195336 5108 195388 5160
rect 197176 5108 197228 5160
rect 551468 5108 551520 5160
rect 106096 5040 106148 5092
rect 187332 5040 187384 5092
rect 107476 4972 107528 5024
rect 189724 4972 189776 5024
rect 200304 5040 200356 5092
rect 201316 5040 201368 5092
rect 204812 5040 204864 5092
rect 204904 5040 204956 5092
rect 554964 5040 555016 5092
rect 107568 4904 107620 4956
rect 193312 4904 193364 4956
rect 108948 4836 109000 4888
rect 193864 4836 193916 4888
rect 110328 4768 110380 4820
rect 198556 4972 198608 5024
rect 558552 4972 558604 5024
rect 194140 4904 194192 4956
rect 194048 4836 194100 4888
rect 196808 4836 196860 4888
rect 198280 4904 198332 4956
rect 562048 4904 562100 4956
rect 204720 4836 204772 4888
rect 204996 4836 205048 4888
rect 569132 4836 569184 4888
rect 195060 4768 195112 4820
rect 203892 4768 203944 4820
rect 204168 4768 204220 4820
rect 581000 4768 581052 4820
rect 100576 4700 100628 4752
rect 162492 4700 162544 4752
rect 191656 4700 191708 4752
rect 530124 4700 530176 4752
rect 99196 4632 99248 4684
rect 157800 4632 157852 4684
rect 190092 4632 190144 4684
rect 526628 4632 526680 4684
rect 96528 4564 96580 4616
rect 147128 4564 147180 4616
rect 147220 4564 147272 4616
rect 195060 4564 195112 4616
rect 195152 4564 195204 4616
rect 523040 4564 523092 4616
rect 99104 4496 99156 4548
rect 154212 4496 154264 4548
rect 188896 4496 188948 4548
rect 519544 4496 519596 4548
rect 96436 4428 96488 4480
rect 143540 4428 143592 4480
rect 146944 4428 146996 4480
rect 182548 4428 182600 4480
rect 188620 4428 188672 4480
rect 195152 4428 195204 4480
rect 93768 4360 93820 4412
rect 136456 4360 136508 4412
rect 142804 4360 142856 4412
rect 186136 4360 186188 4412
rect 187516 4360 187568 4412
rect 515956 4428 516008 4480
rect 195336 4360 195388 4412
rect 512460 4360 512512 4412
rect 93676 4292 93728 4344
rect 132960 4292 133012 4344
rect 173808 4292 173860 4344
rect 458088 4292 458140 4344
rect 92296 4224 92348 4276
rect 126980 4224 127032 4276
rect 172152 4224 172204 4276
rect 450912 4224 450964 4276
rect 99288 4156 99340 4208
rect 21824 4088 21876 4140
rect 24216 4088 24268 4140
rect 24768 4088 24820 4140
rect 27712 4088 27764 4140
rect 28908 4088 28960 4140
rect 29000 4088 29052 4140
rect 65156 4088 65208 4140
rect 84016 4088 84068 4140
rect 96252 4088 96304 4140
rect 97264 4088 97316 4140
rect 103336 4088 103388 4140
rect 171048 4156 171100 4208
rect 447416 4156 447468 4208
rect 156604 4088 156656 4140
rect 220176 4088 220228 4140
rect 390652 4088 390704 4140
rect 436744 4088 436796 4140
rect 442632 4088 442684 4140
rect 479524 4088 479576 4140
rect 480536 4088 480588 4140
rect 65064 4020 65116 4072
rect 85396 4020 85448 4072
rect 94412 4020 94464 4072
rect 94504 4020 94556 4072
rect 99840 4020 99892 4072
rect 100668 4020 100720 4072
rect 160100 4020 160152 4072
rect 215944 4020 215996 4072
rect 404820 4020 404872 4072
rect 26884 3952 26936 4004
rect 63684 3952 63736 4004
rect 88248 3952 88300 4004
rect 114008 3952 114060 4004
rect 146208 3952 146260 4004
rect 348056 3952 348108 4004
rect 475384 3952 475436 4004
rect 510068 3952 510120 4004
rect 18236 3884 18288 3936
rect 63500 3884 63552 3936
rect 89628 3884 89680 3936
rect 115204 3884 115256 3936
rect 147496 3884 147548 3936
rect 351644 3884 351696 3936
rect 472624 3884 472676 3936
rect 506480 3884 506532 3936
rect 20628 3816 20680 3868
rect 64972 3816 65024 3868
rect 89536 3816 89588 3868
rect 118792 3816 118844 3868
rect 147404 3816 147456 3868
rect 354036 3816 354088 3868
rect 468484 3816 468536 3868
rect 505376 3816 505428 3868
rect 15936 3748 15988 3800
rect 55680 3748 55732 3800
rect 55772 3748 55824 3800
rect 61016 3748 61068 3800
rect 89352 3748 89404 3800
rect 116400 3748 116452 3800
rect 147588 3748 147640 3800
rect 355232 3748 355284 3800
rect 421564 3748 421616 3800
rect 423680 3748 423732 3800
rect 432604 3748 432656 3800
rect 460388 3748 460440 3800
rect 461676 3748 461728 3800
rect 498200 3748 498252 3800
rect 12256 3680 12308 3732
rect 60004 3680 60056 3732
rect 60832 3680 60884 3732
rect 74908 3680 74960 3732
rect 81164 3680 81216 3732
rect 85672 3680 85724 3732
rect 89444 3680 89496 3732
rect 119896 3680 119948 3732
rect 120724 3680 120776 3732
rect 129372 3680 129424 3732
rect 148600 3680 148652 3732
rect 358728 3680 358780 3732
rect 447784 3680 447836 3732
rect 7656 3612 7708 3664
rect 55772 3612 55824 3664
rect 5264 3544 5316 3596
rect 60740 3612 60792 3664
rect 2872 3476 2924 3528
rect 59452 3544 59504 3596
rect 59728 3544 59780 3596
rect 63868 3544 63920 3596
rect 64328 3544 64380 3596
rect 74816 3612 74868 3664
rect 91008 3612 91060 3664
rect 122288 3612 122340 3664
rect 150348 3612 150400 3664
rect 365812 3612 365864 3664
rect 443644 3612 443696 3664
rect 69112 3544 69164 3596
rect 70216 3544 70268 3596
rect 73804 3544 73856 3596
rect 76564 3544 76616 3596
rect 77392 3544 77444 3596
rect 78772 3544 78824 3596
rect 82728 3544 82780 3596
rect 87972 3544 88024 3596
rect 90824 3544 90876 3596
rect 123484 3544 123536 3596
rect 153016 3544 153068 3596
rect 153108 3544 153160 3596
rect 372896 3544 372948 3596
rect 374000 3544 374052 3596
rect 375288 3544 375340 3596
rect 56048 3476 56100 3528
rect 57152 3476 57204 3528
rect 58440 3476 58492 3528
rect 59268 3476 59320 3528
rect 59636 3476 59688 3528
rect 60648 3476 60700 3528
rect 63224 3476 63276 3528
rect 74724 3476 74776 3528
rect 76196 3476 76248 3528
rect 77208 3476 77260 3528
rect 79140 3476 79192 3528
rect 79692 3476 79744 3528
rect 81348 3476 81400 3528
rect 84476 3476 84528 3528
rect 87604 3476 87656 3528
rect 89168 3476 89220 3528
rect 90916 3476 90968 3528
rect 124680 3476 124732 3528
rect 137284 3476 137336 3528
rect 140044 3476 140096 3528
rect 376484 3476 376536 3528
rect 398840 3476 398892 3528
rect 400128 3476 400180 3528
rect 414664 3476 414716 3528
rect 416688 3476 416740 3528
rect 423772 3476 423824 3528
rect 424968 3476 425020 3528
rect 425704 3476 425756 3528
rect 427268 3476 427320 3528
rect 448520 3476 448572 3528
rect 449808 3476 449860 3528
rect 454684 3680 454736 3732
rect 494704 3680 494756 3732
rect 450544 3612 450596 3664
rect 491116 3612 491168 3664
rect 537484 3612 537536 3664
rect 550272 3612 550324 3664
rect 481548 3544 481600 3596
rect 481640 3544 481692 3596
rect 482836 3544 482888 3596
rect 517152 3544 517204 3596
rect 544384 3544 544436 3596
rect 557356 3544 557408 3596
rect 512644 3476 512696 3528
rect 513564 3476 513616 3528
rect 526444 3476 526496 3528
rect 527824 3476 527876 3528
rect 530584 3476 530636 3528
rect 531320 3476 531372 3528
rect 533344 3476 533396 3528
rect 553768 3476 553820 3528
rect 572720 3476 572772 3528
rect 573916 3476 573968 3528
rect 1676 3408 1728 3460
rect 59544 3408 59596 3460
rect 65524 3408 65576 3460
rect 66168 3408 66220 3460
rect 66720 3408 66772 3460
rect 67548 3408 67600 3460
rect 67916 3408 67968 3460
rect 68928 3408 68980 3460
rect 72608 3408 72660 3460
rect 73068 3408 73120 3460
rect 82636 3408 82688 3460
rect 91560 3408 91612 3460
rect 92388 3408 92440 3460
rect 131764 3408 131816 3460
rect 148324 3408 148376 3460
rect 150624 3408 150676 3460
rect 154488 3408 154540 3460
rect 379980 3408 380032 3460
rect 429844 3408 429896 3460
rect 583392 3408 583444 3460
rect 8760 3340 8812 3392
rect 9588 3340 9640 3392
rect 9956 3340 10008 3392
rect 10968 3340 11020 3392
rect 11152 3340 11204 3392
rect 12348 3340 12400 3392
rect 17040 3340 17092 3392
rect 17868 3340 17920 3392
rect 23020 3340 23072 3392
rect 29000 3340 29052 3392
rect 32404 3340 32456 3392
rect 33048 3340 33100 3392
rect 33600 3340 33652 3392
rect 34428 3340 34480 3392
rect 19432 3272 19484 3324
rect 26884 3272 26936 3324
rect 28908 3272 28960 3324
rect 66352 3340 66404 3392
rect 88064 3340 88116 3392
rect 112812 3340 112864 3392
rect 136548 3340 136600 3392
rect 306748 3340 306800 3392
rect 307760 3340 307812 3392
rect 309048 3340 309100 3392
rect 316040 3340 316092 3392
rect 317328 3340 317380 3392
rect 332600 3340 332652 3392
rect 333888 3340 333940 3392
rect 347044 3340 347096 3392
rect 349252 3340 349304 3392
rect 473360 3340 473412 3392
rect 474556 3340 474608 3392
rect 481548 3340 481600 3392
rect 487620 3340 487672 3392
rect 547880 3340 547932 3392
rect 549076 3340 549128 3392
rect 34796 3272 34848 3324
rect 35808 3272 35860 3324
rect 40684 3272 40736 3324
rect 41328 3272 41380 3324
rect 41880 3272 41932 3324
rect 43444 3272 43496 3324
rect 44272 3272 44324 3324
rect 45376 3272 45428 3324
rect 45468 3272 45520 3324
rect 66536 3272 66588 3324
rect 88156 3272 88208 3324
rect 111616 3272 111668 3324
rect 136364 3272 136416 3324
rect 305552 3272 305604 3324
rect 31300 3204 31352 3256
rect 67824 3204 67876 3256
rect 86776 3204 86828 3256
rect 109316 3204 109368 3256
rect 193220 3204 193272 3256
rect 194416 3204 194468 3256
rect 203524 3204 203576 3256
rect 206192 3204 206244 3256
rect 220084 3204 220136 3256
rect 387156 3204 387208 3256
rect 30104 3136 30156 3188
rect 45376 3136 45428 3188
rect 26516 3068 26568 3120
rect 27528 3068 27580 3120
rect 37188 3068 37240 3120
rect 69204 3136 69256 3188
rect 86868 3136 86920 3188
rect 108120 3136 108172 3188
rect 123576 3136 123628 3188
rect 125876 3136 125928 3188
rect 131028 3136 131080 3188
rect 284300 3136 284352 3188
rect 48964 3068 49016 3120
rect 49608 3068 49660 3120
rect 50160 3068 50212 3120
rect 50988 3068 51040 3120
rect 52552 3068 52604 3120
rect 53656 3068 53708 3120
rect 25320 3000 25372 3052
rect 26148 3000 26200 3052
rect 35992 3000 36044 3052
rect 68008 3068 68060 3120
rect 86684 3068 86736 3120
rect 105728 3068 105780 3120
rect 128268 3068 128320 3120
rect 272432 3068 272484 3120
rect 417516 3068 417568 3120
rect 420184 3068 420236 3120
rect 53840 3000 53892 3052
rect 70584 3000 70636 3052
rect 75000 3000 75052 3052
rect 76656 3000 76708 3052
rect 85488 3000 85540 3052
rect 102232 3000 102284 3052
rect 104164 3000 104216 3052
rect 121092 3000 121144 3052
rect 222936 3000 222988 3052
rect 350448 3000 350500 3052
rect 407764 3000 407816 3052
rect 409604 3000 409656 3052
rect 45468 2932 45520 2984
rect 70676 2932 70728 2984
rect 84108 2932 84160 2984
rect 95148 2932 95200 2984
rect 102876 2932 102928 2984
rect 117596 2932 117648 2984
rect 220268 2932 220320 2984
rect 337476 2932 337528 2984
rect 368480 2932 368532 2984
rect 371700 2932 371752 2984
rect 51356 2864 51408 2916
rect 72056 2864 72108 2916
rect 81256 2864 81308 2916
rect 82084 2864 82136 2916
rect 83924 2864 83976 2916
rect 92756 2864 92808 2916
rect 94412 2864 94464 2916
rect 98644 2864 98696 2916
rect 102784 2864 102836 2916
rect 110512 2864 110564 2916
rect 222844 2864 222896 2916
rect 294880 2864 294932 2916
rect 519636 2864 519688 2916
rect 524236 2864 524288 2916
rect 43076 2796 43128 2848
rect 53840 2796 53892 2848
rect 57244 2796 57296 2848
rect 68284 2796 68336 2848
rect 81072 2796 81124 2848
rect 86868 2796 86920 2848
rect 101404 2796 101456 2848
rect 106924 2796 106976 2848
rect 223028 2796 223080 2848
rect 283104 2796 283156 2848
rect 242900 2728 242952 2780
rect 244096 2728 244148 2780
rect 160008 2116 160060 2168
rect 401324 2116 401376 2168
rect 179052 2048 179104 2100
rect 479340 2048 479392 2100
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 412652 703582 413508 703610
rect 8128 702434 8156 703520
rect 8128 702406 8248 702434
rect 2778 684312 2834 684321
rect 2778 684247 2834 684256
rect 2792 683738 2820 684247
rect 2780 683732 2832 683738
rect 2780 683674 2832 683680
rect 4804 683732 4856 683738
rect 4804 683674 4856 683680
rect 3514 671256 3570 671265
rect 3514 671191 3570 671200
rect 3528 670750 3556 671191
rect 3516 670744 3568 670750
rect 3516 670686 3568 670692
rect 3422 658200 3478 658209
rect 3422 658135 3478 658144
rect 3436 656946 3464 658135
rect 3424 656940 3476 656946
rect 3424 656882 3476 656888
rect 3424 632120 3476 632126
rect 3422 632088 3424 632097
rect 3476 632088 3478 632097
rect 3422 632023 3478 632032
rect 3146 619168 3202 619177
rect 3146 619103 3202 619112
rect 3160 618322 3188 619103
rect 3148 618316 3200 618322
rect 3148 618258 3200 618264
rect 3238 606112 3294 606121
rect 3238 606047 3294 606056
rect 3252 605878 3280 606047
rect 3240 605872 3292 605878
rect 3240 605814 3292 605820
rect 3330 580000 3386 580009
rect 3330 579935 3386 579944
rect 3344 579698 3372 579935
rect 3332 579692 3384 579698
rect 3332 579634 3384 579640
rect 3422 566944 3478 566953
rect 3422 566879 3478 566888
rect 3436 565894 3464 566879
rect 3424 565888 3476 565894
rect 3424 565830 3476 565836
rect 3422 553888 3478 553897
rect 3422 553823 3478 553832
rect 3436 553450 3464 553823
rect 3424 553444 3476 553450
rect 3424 553386 3476 553392
rect 3422 527912 3478 527921
rect 3422 527847 3478 527856
rect 3436 527202 3464 527847
rect 3424 527196 3476 527202
rect 3424 527138 3476 527144
rect 3422 514856 3478 514865
rect 3422 514791 3424 514800
rect 3476 514791 3478 514800
rect 3424 514762 3476 514768
rect 3054 501800 3110 501809
rect 3054 501735 3110 501744
rect 3068 501022 3096 501735
rect 3056 501016 3108 501022
rect 3056 500958 3108 500964
rect 3422 475688 3478 475697
rect 3422 475623 3478 475632
rect 3436 474774 3464 475623
rect 3424 474768 3476 474774
rect 3424 474710 3476 474716
rect 3238 462632 3294 462641
rect 3238 462567 3294 462576
rect 3252 462398 3280 462567
rect 3240 462392 3292 462398
rect 3240 462334 3292 462340
rect 3146 449576 3202 449585
rect 3146 449511 3202 449520
rect 3160 448594 3188 449511
rect 3148 448588 3200 448594
rect 3148 448530 3200 448536
rect 3422 423600 3478 423609
rect 3422 423535 3478 423544
rect 3436 422346 3464 423535
rect 3424 422340 3476 422346
rect 3424 422282 3476 422288
rect 3146 410544 3202 410553
rect 3146 410479 3202 410488
rect 3160 409902 3188 410479
rect 3148 409896 3200 409902
rect 3148 409838 3200 409844
rect 3424 397520 3476 397526
rect 3422 397488 3424 397497
rect 3476 397488 3478 397497
rect 3422 397423 3478 397432
rect 3422 371376 3478 371385
rect 3422 371311 3478 371320
rect 3436 371278 3464 371311
rect 3424 371272 3476 371278
rect 3424 371214 3476 371220
rect 3146 358456 3202 358465
rect 3146 358391 3202 358400
rect 3160 357474 3188 358391
rect 3148 357468 3200 357474
rect 3148 357410 3200 357416
rect 3330 345400 3386 345409
rect 3330 345335 3386 345344
rect 3344 345098 3372 345335
rect 3332 345092 3384 345098
rect 3332 345034 3384 345040
rect 3422 319288 3478 319297
rect 3422 319223 3478 319232
rect 3436 318850 3464 319223
rect 3424 318844 3476 318850
rect 3424 318786 3476 318792
rect 3238 306232 3294 306241
rect 3238 306167 3294 306176
rect 3252 305046 3280 306167
rect 3240 305040 3292 305046
rect 3240 304982 3292 304988
rect 3422 293176 3478 293185
rect 3422 293111 3478 293120
rect 3436 292602 3464 293111
rect 3424 292596 3476 292602
rect 3424 292538 3476 292544
rect 3054 267200 3110 267209
rect 3054 267135 3110 267144
rect 3068 266422 3096 267135
rect 3056 266416 3108 266422
rect 3056 266358 3108 266364
rect 4816 260506 4844 683674
rect 8220 263498 8248 702406
rect 24320 700330 24348 703520
rect 40512 700398 40540 703520
rect 40500 700392 40552 700398
rect 40500 700334 40552 700340
rect 41328 700392 41380 700398
rect 41328 700334 41380 700340
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 33784 700324 33836 700330
rect 33784 700266 33836 700272
rect 15844 656940 15896 656946
rect 15844 656882 15896 656888
rect 14464 632120 14516 632126
rect 14464 632062 14516 632068
rect 11704 579692 11756 579698
rect 11704 579634 11756 579640
rect 8208 263492 8260 263498
rect 8208 263434 8260 263440
rect 11716 262206 11744 579634
rect 14476 290494 14504 632062
rect 14464 290488 14516 290494
rect 14464 290430 14516 290436
rect 11704 262200 11756 262206
rect 11704 262142 11756 262148
rect 15856 260574 15884 656882
rect 22744 605872 22796 605878
rect 22744 605814 22796 605820
rect 17224 527196 17276 527202
rect 17224 527138 17276 527144
rect 17236 261458 17264 527138
rect 18604 474768 18656 474774
rect 18604 474710 18656 474716
rect 18616 297430 18644 474710
rect 21364 422340 21416 422346
rect 21364 422282 21416 422288
rect 18604 297424 18656 297430
rect 18604 297366 18656 297372
rect 21376 262138 21404 422282
rect 21364 262132 21416 262138
rect 21364 262074 21416 262080
rect 17224 261452 17276 261458
rect 17224 261394 17276 261400
rect 22756 261390 22784 605814
rect 25504 553444 25556 553450
rect 25504 553386 25556 553392
rect 22744 261384 22796 261390
rect 22744 261326 22796 261332
rect 25516 260642 25544 553386
rect 29644 501016 29696 501022
rect 29644 500958 29696 500964
rect 29656 263566 29684 500958
rect 32404 448588 32456 448594
rect 32404 448530 32456 448536
rect 29644 263560 29696 263566
rect 29644 263502 29696 263508
rect 32416 262818 32444 448530
rect 32404 262812 32456 262818
rect 32404 262754 32456 262760
rect 33796 262614 33824 700266
rect 35164 670744 35216 670750
rect 35164 670686 35216 670692
rect 35176 264178 35204 670686
rect 36544 618316 36596 618322
rect 36544 618258 36596 618264
rect 35164 264172 35216 264178
rect 35164 264114 35216 264120
rect 36556 262682 36584 618258
rect 39304 565888 39356 565894
rect 39304 565830 39356 565836
rect 39316 262750 39344 565830
rect 39304 262744 39356 262750
rect 39304 262686 39356 262692
rect 36544 262676 36596 262682
rect 36544 262618 36596 262624
rect 33784 262608 33836 262614
rect 33784 262550 33836 262556
rect 41340 261050 41368 700334
rect 72988 700330 73016 703520
rect 58808 700324 58860 700330
rect 58808 700266 58860 700272
rect 72976 700324 73028 700330
rect 72976 700266 73028 700272
rect 43444 514820 43496 514826
rect 43444 514762 43496 514768
rect 43456 264790 43484 514762
rect 58714 489968 58770 489977
rect 58714 489903 58770 489912
rect 53654 488880 53710 488889
rect 53654 488815 53710 488824
rect 53562 484800 53618 484809
rect 53562 484735 53618 484744
rect 53378 484664 53434 484673
rect 53378 484599 53434 484608
rect 47584 462392 47636 462398
rect 47584 462334 47636 462340
rect 47596 264858 47624 462334
rect 50344 409896 50396 409902
rect 50344 409838 50396 409844
rect 50356 264926 50384 409838
rect 52276 399764 52328 399770
rect 52276 399706 52328 399712
rect 52184 395412 52236 395418
rect 52184 395354 52236 395360
rect 52092 268388 52144 268394
rect 52092 268330 52144 268336
rect 52000 265804 52052 265810
rect 52000 265746 52052 265752
rect 50344 264920 50396 264926
rect 50344 264862 50396 264868
rect 47584 264852 47636 264858
rect 47584 264794 47636 264800
rect 43444 264784 43496 264790
rect 43444 264726 43496 264732
rect 41328 261044 41380 261050
rect 41328 260986 41380 260992
rect 25504 260636 25556 260642
rect 25504 260578 25556 260584
rect 15844 260568 15896 260574
rect 15844 260510 15896 260516
rect 4804 260500 4856 260506
rect 4804 260442 4856 260448
rect 3422 254144 3478 254153
rect 3422 254079 3478 254088
rect 3436 249121 3464 254079
rect 3422 249112 3478 249121
rect 3422 249047 3478 249056
rect 4066 241088 4122 241097
rect 4122 241046 4200 241074
rect 4066 241023 4122 241032
rect 4172 235249 4200 241046
rect 4158 235240 4214 235249
rect 4158 235175 4214 235184
rect 21362 233744 21418 233753
rect 21362 233679 21418 233688
rect 18602 233608 18658 233617
rect 18602 233543 18658 233552
rect 14462 231976 14518 231985
rect 14462 231911 14518 231920
rect 11702 231160 11758 231169
rect 11702 231095 11758 231104
rect 7562 231024 7618 231033
rect 7562 230959 7618 230968
rect 4802 230888 4858 230897
rect 4802 230823 4858 230832
rect 3606 228576 3662 228585
rect 3606 228511 3662 228520
rect 3422 228304 3478 228313
rect 3422 228239 3478 228248
rect 2780 215280 2832 215286
rect 2780 215222 2832 215228
rect 2792 214985 2820 215222
rect 2778 214976 2834 214985
rect 2778 214911 2834 214920
rect 3148 189032 3200 189038
rect 3148 188974 3200 188980
rect 3160 188873 3188 188974
rect 3146 188864 3202 188873
rect 3146 188799 3202 188808
rect 3332 162988 3384 162994
rect 3332 162930 3384 162936
rect 3344 162897 3372 162930
rect 3330 162888 3386 162897
rect 3330 162823 3386 162832
rect 3332 137964 3384 137970
rect 3332 137906 3384 137912
rect 3344 136785 3372 137906
rect 3330 136776 3386 136785
rect 3330 136711 3386 136720
rect 3148 111784 3200 111790
rect 3148 111726 3200 111732
rect 3160 110673 3188 111726
rect 3146 110664 3202 110673
rect 3146 110599 3202 110608
rect 3240 97980 3292 97986
rect 3240 97922 3292 97928
rect 3252 97617 3280 97922
rect 3238 97608 3294 97617
rect 3238 97543 3294 97552
rect 3332 85536 3384 85542
rect 3332 85478 3384 85484
rect 3344 84697 3372 85478
rect 3330 84688 3386 84697
rect 3330 84623 3386 84632
rect 3332 71732 3384 71738
rect 3332 71674 3384 71680
rect 3344 71641 3372 71674
rect 3330 71632 3386 71641
rect 3330 71567 3386 71576
rect 3436 45529 3464 228239
rect 3514 227080 3570 227089
rect 3514 227015 3570 227024
rect 3528 58585 3556 227015
rect 3620 201929 3648 228511
rect 3698 227216 3754 227225
rect 3698 227151 3754 227160
rect 3606 201920 3662 201929
rect 3606 201855 3662 201864
rect 3712 149841 3740 227151
rect 4816 215286 4844 230823
rect 4804 215280 4856 215286
rect 4804 215222 4856 215228
rect 7576 162994 7604 230959
rect 7564 162988 7616 162994
rect 7564 162930 7616 162936
rect 3698 149832 3754 149841
rect 3698 149767 3754 149776
rect 11716 111790 11744 231095
rect 11704 111784 11756 111790
rect 11704 111726 11756 111732
rect 14476 71738 14504 231911
rect 15842 230752 15898 230761
rect 15842 230687 15898 230696
rect 14464 71732 14516 71738
rect 14464 71674 14516 71680
rect 3514 58576 3570 58585
rect 3514 58511 3570 58520
rect 12346 57624 12402 57633
rect 12346 57559 12402 57568
rect 10966 57488 11022 57497
rect 10966 57423 11022 57432
rect 9586 57352 9642 57361
rect 6828 57316 6880 57322
rect 9586 57287 9642 57296
rect 6828 57258 6880 57264
rect 4066 57216 4122 57225
rect 4066 57151 4122 57160
rect 3422 45520 3478 45529
rect 3422 45455 3478 45464
rect 2872 33108 2924 33114
rect 2872 33050 2924 33056
rect 2884 32473 2912 33050
rect 2870 32464 2926 32473
rect 2870 32399 2926 32408
rect 3424 20664 3476 20670
rect 3424 20606 3476 20612
rect 3436 19417 3464 20606
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 3424 6860 3476 6866
rect 3424 6802 3476 6808
rect 3436 6497 3464 6802
rect 3422 6488 3478 6497
rect 3422 6423 3478 6432
rect 2872 3528 2924 3534
rect 2872 3470 2924 3476
rect 1676 3460 1728 3466
rect 1676 3402 1728 3408
rect 570 3360 626 3369
rect 570 3295 626 3304
rect 584 480 612 3295
rect 1688 480 1716 3402
rect 2884 480 2912 3470
rect 4080 480 4108 57151
rect 6840 6914 6868 57258
rect 6472 6886 6868 6914
rect 5264 3596 5316 3602
rect 5264 3538 5316 3544
rect 5276 480 5304 3538
rect 6472 480 6500 6886
rect 7656 3664 7708 3670
rect 7656 3606 7708 3612
rect 7668 480 7696 3606
rect 9600 3398 9628 57287
rect 10980 3398 11008 57423
rect 12256 3732 12308 3738
rect 12256 3674 12308 3680
rect 8760 3392 8812 3398
rect 8760 3334 8812 3340
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9956 3392 10008 3398
rect 9956 3334 10008 3340
rect 10968 3392 11020 3398
rect 10968 3334 11020 3340
rect 11152 3392 11204 3398
rect 11152 3334 11204 3340
rect 8772 480 8800 3334
rect 9968 480 9996 3334
rect 11164 480 11192 3334
rect 12268 1850 12296 3674
rect 12360 3398 12388 57559
rect 15106 57080 15162 57089
rect 15106 57015 15162 57024
rect 13726 56944 13782 56953
rect 13726 56879 13782 56888
rect 13740 6914 13768 56879
rect 15120 6914 15148 57015
rect 15856 33114 15884 230687
rect 17222 226808 17278 226817
rect 17222 226743 17278 226752
rect 17236 189038 17264 226743
rect 17224 189032 17276 189038
rect 17224 188974 17276 188980
rect 18616 137970 18644 233543
rect 18604 137964 18656 137970
rect 18604 137906 18656 137912
rect 21376 85542 21404 233679
rect 25502 229528 25558 229537
rect 25502 229463 25558 229472
rect 22742 228440 22798 228449
rect 22742 228375 22798 228384
rect 21364 85536 21416 85542
rect 21364 85478 21416 85484
rect 17866 56808 17922 56817
rect 17866 56743 17922 56752
rect 15844 33108 15896 33114
rect 15844 33050 15896 33056
rect 13556 6886 13768 6914
rect 14752 6886 15148 6914
rect 12348 3392 12400 3398
rect 12348 3334 12400 3340
rect 12268 1822 12388 1850
rect 12360 480 12388 1822
rect 13556 480 13584 6886
rect 14752 480 14780 6886
rect 15936 3800 15988 3806
rect 15936 3742 15988 3748
rect 15948 480 15976 3742
rect 17880 3398 17908 56743
rect 22756 6866 22784 228375
rect 25516 97986 25544 229463
rect 29642 229392 29698 229401
rect 29642 229327 29698 229336
rect 25504 97980 25556 97986
rect 25504 97922 25556 97928
rect 28908 57520 28960 57526
rect 28908 57462 28960 57468
rect 26148 57452 26200 57458
rect 26148 57394 26200 57400
rect 24768 57248 24820 57254
rect 24768 57190 24820 57196
rect 22744 6860 22796 6866
rect 22744 6802 22796 6808
rect 24780 4146 24808 57190
rect 21824 4140 21876 4146
rect 21824 4082 21876 4088
rect 24216 4140 24268 4146
rect 24216 4082 24268 4088
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 18236 3936 18288 3942
rect 18236 3878 18288 3884
rect 17040 3392 17092 3398
rect 17040 3334 17092 3340
rect 17868 3392 17920 3398
rect 17868 3334 17920 3340
rect 17052 480 17080 3334
rect 18248 480 18276 3878
rect 20628 3868 20680 3874
rect 20628 3810 20680 3816
rect 19432 3324 19484 3330
rect 19432 3266 19484 3272
rect 19444 480 19472 3266
rect 20640 480 20668 3810
rect 21836 480 21864 4082
rect 23020 3392 23072 3398
rect 23020 3334 23072 3340
rect 23032 480 23060 3334
rect 24228 480 24256 4082
rect 26160 3058 26188 57394
rect 27528 57384 27580 57390
rect 27528 57326 27580 57332
rect 26884 4004 26936 4010
rect 26884 3946 26936 3952
rect 26896 3330 26924 3946
rect 26884 3324 26936 3330
rect 26884 3266 26936 3272
rect 27540 3126 27568 57326
rect 28920 4146 28948 57462
rect 29656 20670 29684 229327
rect 52012 157350 52040 265746
rect 52000 157344 52052 157350
rect 52000 157286 52052 157292
rect 52104 153882 52132 268330
rect 52092 153876 52144 153882
rect 52092 153818 52144 153824
rect 52196 113150 52224 395354
rect 52184 113144 52236 113150
rect 52184 113086 52236 113092
rect 52288 88330 52316 399706
rect 52368 395480 52420 395486
rect 52368 395422 52420 395428
rect 52276 88324 52328 88330
rect 52276 88266 52328 88272
rect 52380 70378 52408 395422
rect 53196 262064 53248 262070
rect 53196 262006 53248 262012
rect 53208 121446 53236 262006
rect 53288 260160 53340 260166
rect 53288 260102 53340 260108
rect 53196 121440 53248 121446
rect 53196 121382 53248 121388
rect 53300 82822 53328 260102
rect 53392 192710 53420 484599
rect 53472 399832 53524 399838
rect 53472 399774 53524 399780
rect 53380 192704 53432 192710
rect 53380 192646 53432 192652
rect 53484 105602 53512 399774
rect 53576 144634 53604 484735
rect 53564 144628 53616 144634
rect 53564 144570 53616 144576
rect 53668 142118 53696 488815
rect 55034 487928 55090 487937
rect 55034 487863 55090 487872
rect 54942 487520 54998 487529
rect 54942 487455 54998 487464
rect 53746 487248 53802 487257
rect 53746 487183 53802 487192
rect 53656 142112 53708 142118
rect 53656 142054 53708 142060
rect 53760 136610 53788 487183
rect 54668 395684 54720 395690
rect 54668 395626 54720 395632
rect 54484 264444 54536 264450
rect 54484 264386 54536 264392
rect 54392 264376 54444 264382
rect 54392 264318 54444 264324
rect 54300 264308 54352 264314
rect 54300 264250 54352 264256
rect 54312 182850 54340 264250
rect 54300 182844 54352 182850
rect 54300 182786 54352 182792
rect 54404 169726 54432 264318
rect 54392 169720 54444 169726
rect 54392 169662 54444 169668
rect 54496 151774 54524 264386
rect 54576 225412 54628 225418
rect 54576 225354 54628 225360
rect 54484 151768 54536 151774
rect 54484 151710 54536 151716
rect 53748 136604 53800 136610
rect 53748 136546 53800 136552
rect 53472 105596 53524 105602
rect 53472 105538 53524 105544
rect 54588 100706 54616 225354
rect 54680 195974 54708 395626
rect 54852 395616 54904 395622
rect 54852 395558 54904 395564
rect 54760 395344 54812 395350
rect 54760 395286 54812 395292
rect 54668 195968 54720 195974
rect 54668 195910 54720 195916
rect 54772 160070 54800 395286
rect 54760 160064 54812 160070
rect 54760 160006 54812 160012
rect 54864 103494 54892 395558
rect 54956 187678 54984 487455
rect 54944 187672 54996 187678
rect 54944 187614 54996 187620
rect 55048 162858 55076 487863
rect 56874 487384 56930 487393
rect 56874 487319 56930 487328
rect 56506 486024 56562 486033
rect 56506 485959 56562 485968
rect 55126 484936 55182 484945
rect 55126 484871 55182 484880
rect 55036 162852 55088 162858
rect 55036 162794 55088 162800
rect 55140 126954 55168 484871
rect 56414 483984 56470 483993
rect 56414 483919 56470 483928
rect 56324 395752 56376 395758
rect 56324 395694 56376 395700
rect 56232 265668 56284 265674
rect 56232 265610 56284 265616
rect 56048 263968 56100 263974
rect 56048 263910 56100 263916
rect 55956 262540 56008 262546
rect 55956 262482 56008 262488
rect 55864 261180 55916 261186
rect 55864 261122 55916 261128
rect 55678 226536 55734 226545
rect 55678 226471 55734 226480
rect 55128 126948 55180 126954
rect 55128 126890 55180 126896
rect 54852 103488 54904 103494
rect 54852 103430 54904 103436
rect 54576 100700 54628 100706
rect 54576 100642 54628 100648
rect 53288 82816 53340 82822
rect 53288 82758 53340 82764
rect 52368 70372 52420 70378
rect 52368 70314 52420 70320
rect 45468 57928 45520 57934
rect 45468 57870 45520 57876
rect 41328 57860 41380 57866
rect 41328 57802 41380 57808
rect 35808 57792 35860 57798
rect 35808 57734 35860 57740
rect 34428 57656 34480 57662
rect 34428 57598 34480 57604
rect 33048 57588 33100 57594
rect 33048 57530 33100 57536
rect 29644 20664 29696 20670
rect 29644 20606 29696 20612
rect 27712 4140 27764 4146
rect 27712 4082 27764 4088
rect 28908 4140 28960 4146
rect 28908 4082 28960 4088
rect 29000 4140 29052 4146
rect 29000 4082 29052 4088
rect 26516 3120 26568 3126
rect 26516 3062 26568 3068
rect 27528 3120 27580 3126
rect 27528 3062 27580 3068
rect 25320 3052 25372 3058
rect 25320 2994 25372 3000
rect 26148 3052 26200 3058
rect 26148 2994 26200 3000
rect 25332 480 25360 2994
rect 26528 480 26556 3062
rect 27724 480 27752 4082
rect 29012 3398 29040 4082
rect 33060 3398 33088 57530
rect 34440 3398 34468 57598
rect 29000 3392 29052 3398
rect 29000 3334 29052 3340
rect 32404 3392 32456 3398
rect 32404 3334 32456 3340
rect 33048 3392 33100 3398
rect 33048 3334 33100 3340
rect 33600 3392 33652 3398
rect 33600 3334 33652 3340
rect 34428 3392 34480 3398
rect 34428 3334 34480 3340
rect 28908 3324 28960 3330
rect 28908 3266 28960 3272
rect 28920 480 28948 3266
rect 31300 3256 31352 3262
rect 31300 3198 31352 3204
rect 30104 3188 30156 3194
rect 30104 3130 30156 3136
rect 30116 480 30144 3130
rect 31312 480 31340 3198
rect 32416 480 32444 3334
rect 33612 480 33640 3334
rect 35820 3330 35848 57734
rect 39948 57724 40000 57730
rect 39948 57666 40000 57672
rect 38568 54528 38620 54534
rect 38568 54470 38620 54476
rect 38580 6914 38608 54470
rect 39960 6914 39988 57666
rect 38396 6886 38608 6914
rect 39592 6886 39988 6914
rect 34796 3324 34848 3330
rect 34796 3266 34848 3272
rect 35808 3324 35860 3330
rect 35808 3266 35860 3272
rect 34808 480 34836 3266
rect 37188 3120 37240 3126
rect 37188 3062 37240 3068
rect 35992 3052 36044 3058
rect 35992 2994 36044 3000
rect 36004 480 36032 2994
rect 37200 480 37228 3062
rect 38396 480 38424 6886
rect 39592 480 39620 6886
rect 41340 3330 41368 57802
rect 43444 57180 43496 57186
rect 43444 57122 43496 57128
rect 43456 3330 43484 57122
rect 45480 6914 45508 57870
rect 46848 57112 46900 57118
rect 46848 57054 46900 57060
rect 46860 6914 46888 57054
rect 49608 57044 49660 57050
rect 49608 56986 49660 56992
rect 48228 56976 48280 56982
rect 48228 56918 48280 56924
rect 48240 6914 48268 56918
rect 45388 6886 45508 6914
rect 46676 6886 46888 6914
rect 47872 6886 48268 6914
rect 45388 3330 45416 6886
rect 40684 3324 40736 3330
rect 40684 3266 40736 3272
rect 41328 3324 41380 3330
rect 41328 3266 41380 3272
rect 41880 3324 41932 3330
rect 41880 3266 41932 3272
rect 43444 3324 43496 3330
rect 43444 3266 43496 3272
rect 44272 3324 44324 3330
rect 44272 3266 44324 3272
rect 45376 3324 45428 3330
rect 45376 3266 45428 3272
rect 45468 3324 45520 3330
rect 45468 3266 45520 3272
rect 40696 480 40724 3266
rect 41892 480 41920 3266
rect 43076 2848 43128 2854
rect 43076 2790 43128 2796
rect 43088 480 43116 2790
rect 44284 480 44312 3266
rect 45480 3210 45508 3266
rect 45388 3194 45508 3210
rect 45376 3188 45508 3194
rect 45428 3182 45508 3188
rect 45376 3130 45428 3136
rect 45468 2984 45520 2990
rect 45468 2926 45520 2932
rect 45480 480 45508 2926
rect 46676 480 46704 6886
rect 47872 480 47900 6886
rect 49620 3126 49648 56986
rect 53748 56908 53800 56914
rect 53748 56850 53800 56856
rect 53656 56840 53708 56846
rect 53656 56782 53708 56788
rect 50988 54596 51040 54602
rect 50988 54538 51040 54544
rect 51000 3126 51028 54538
rect 53668 3126 53696 56782
rect 48964 3120 49016 3126
rect 48964 3062 49016 3068
rect 49608 3120 49660 3126
rect 49608 3062 49660 3068
rect 50160 3120 50212 3126
rect 50160 3062 50212 3068
rect 50988 3120 51040 3126
rect 50988 3062 51040 3068
rect 52552 3120 52604 3126
rect 52552 3062 52604 3068
rect 53656 3120 53708 3126
rect 53656 3062 53708 3068
rect 48976 480 49004 3062
rect 50172 480 50200 3062
rect 51356 2916 51408 2922
rect 51356 2858 51408 2864
rect 51368 480 51396 2858
rect 52564 480 52592 3062
rect 53760 480 53788 56850
rect 55128 56772 55180 56778
rect 55128 56714 55180 56720
rect 55140 6914 55168 56714
rect 55692 20670 55720 226471
rect 55770 226400 55826 226409
rect 55770 226335 55826 226344
rect 55784 55894 55812 226335
rect 55876 207369 55904 261122
rect 55862 207360 55918 207369
rect 55862 207295 55918 207304
rect 55968 189553 55996 262482
rect 55954 189544 56010 189553
rect 55954 189479 56010 189488
rect 56060 177585 56088 263910
rect 56140 260228 56192 260234
rect 56140 260170 56192 260176
rect 56046 177576 56102 177585
rect 56046 177511 56102 177520
rect 56152 73273 56180 260170
rect 56244 222329 56272 265610
rect 56230 222320 56286 222329
rect 56230 222255 56286 222264
rect 56336 147801 56364 395694
rect 56428 216345 56456 483919
rect 56414 216336 56470 216345
rect 56414 216271 56470 216280
rect 56322 147792 56378 147801
rect 56322 147727 56378 147736
rect 56520 108390 56548 485959
rect 56690 435432 56746 435441
rect 56690 435367 56746 435376
rect 56598 407552 56654 407561
rect 56598 407487 56654 407496
rect 56508 108384 56560 108390
rect 56508 108326 56560 108332
rect 56138 73264 56194 73273
rect 56138 73199 56194 73208
rect 56612 59294 56640 407487
rect 56704 59362 56732 435367
rect 56782 225992 56838 226001
rect 56782 225927 56838 225936
rect 56796 171601 56824 225927
rect 56782 171592 56838 171601
rect 56782 171527 56838 171536
rect 56888 64297 56916 487319
rect 58622 485072 58678 485081
rect 58622 485007 58678 485016
rect 57518 484256 57574 484265
rect 57518 484191 57574 484200
rect 57426 432440 57482 432449
rect 57426 432375 57482 432384
rect 57334 430672 57390 430681
rect 57334 430607 57390 430616
rect 57242 429448 57298 429457
rect 57242 429383 57298 429392
rect 57152 265872 57204 265878
rect 57152 265814 57204 265820
rect 57058 237960 57114 237969
rect 57058 237895 57114 237904
rect 57072 109041 57100 237895
rect 57164 118017 57192 265814
rect 57256 225418 57284 429383
rect 57348 399498 57376 430607
rect 57336 399492 57388 399498
rect 57336 399434 57388 399440
rect 57334 239456 57390 239465
rect 57334 239391 57390 239400
rect 57244 225412 57296 225418
rect 57244 225354 57296 225360
rect 57244 187672 57296 187678
rect 57244 187614 57296 187620
rect 57256 186561 57284 187614
rect 57242 186552 57298 186561
rect 57242 186487 57298 186496
rect 57150 118008 57206 118017
rect 57150 117943 57206 117952
rect 57058 109032 57114 109041
rect 57058 108967 57114 108976
rect 57244 108384 57296 108390
rect 57244 108326 57296 108332
rect 57256 84194 57284 108326
rect 57164 84166 57284 84194
rect 57164 79257 57192 84166
rect 57244 82816 57296 82822
rect 57244 82758 57296 82764
rect 57256 82249 57284 82758
rect 57242 82240 57298 82249
rect 57242 82175 57298 82184
rect 57150 79248 57206 79257
rect 57150 79183 57206 79192
rect 56874 64288 56930 64297
rect 56874 64223 56930 64232
rect 57348 61441 57376 239391
rect 57440 175234 57468 432375
rect 57532 210361 57560 484191
rect 57610 436384 57666 436393
rect 57610 436319 57666 436328
rect 57518 210352 57574 210361
rect 57518 210287 57574 210296
rect 57520 195968 57572 195974
rect 57520 195910 57572 195916
rect 57532 195401 57560 195910
rect 57518 195392 57574 195401
rect 57518 195327 57574 195336
rect 57520 192704 57572 192710
rect 57520 192646 57572 192652
rect 57532 192545 57560 192646
rect 57518 192536 57574 192545
rect 57518 192471 57574 192480
rect 57518 183560 57574 183569
rect 57518 183495 57574 183504
rect 57532 182850 57560 183495
rect 57520 182844 57572 182850
rect 57520 182786 57572 182792
rect 57520 175636 57572 175642
rect 57520 175578 57572 175584
rect 57428 175228 57480 175234
rect 57428 175170 57480 175176
rect 57428 162852 57480 162858
rect 57428 162794 57480 162800
rect 57440 162625 57468 162794
rect 57426 162616 57482 162625
rect 57426 162551 57482 162560
rect 57428 157344 57480 157350
rect 57428 157286 57480 157292
rect 57440 156777 57468 157286
rect 57426 156768 57482 156777
rect 57426 156703 57482 156712
rect 57428 153876 57480 153882
rect 57428 153818 57480 153824
rect 57440 153785 57468 153818
rect 57426 153776 57482 153785
rect 57426 153711 57482 153720
rect 57428 151768 57480 151774
rect 57428 151710 57480 151716
rect 57440 150793 57468 151710
rect 57426 150784 57482 150793
rect 57426 150719 57482 150728
rect 57426 144800 57482 144809
rect 57426 144735 57482 144744
rect 57440 144634 57468 144735
rect 57428 144628 57480 144634
rect 57428 144570 57480 144576
rect 57532 91225 57560 175578
rect 57624 137494 57652 436319
rect 57702 433392 57758 433401
rect 57702 433327 57758 433336
rect 57716 399566 57744 433327
rect 57886 427952 57942 427961
rect 57886 427887 57942 427896
rect 57794 410000 57850 410009
rect 57794 409935 57850 409944
rect 57808 399702 57836 409935
rect 57796 399696 57848 399702
rect 57796 399638 57848 399644
rect 57900 399634 57928 427887
rect 57888 399628 57940 399634
rect 57888 399570 57940 399576
rect 57704 399560 57756 399566
rect 57704 399502 57756 399508
rect 58440 397044 58492 397050
rect 58440 396986 58492 396992
rect 58346 242176 58402 242185
rect 58346 242111 58402 242120
rect 58254 236600 58310 236609
rect 58254 236535 58310 236544
rect 58162 232656 58218 232665
rect 58162 232591 58218 232600
rect 57794 227760 57850 227769
rect 57794 227695 57850 227704
rect 57702 226264 57758 226273
rect 57702 226199 57758 226208
rect 57612 137488 57664 137494
rect 57612 137430 57664 137436
rect 57612 136604 57664 136610
rect 57612 136546 57664 136552
rect 57624 135833 57652 136546
rect 57610 135824 57666 135833
rect 57610 135759 57666 135768
rect 57610 126984 57666 126993
rect 57610 126919 57612 126928
rect 57664 126919 57666 126928
rect 57612 126890 57664 126896
rect 57612 121440 57664 121446
rect 57612 121382 57664 121388
rect 57624 121009 57652 121382
rect 57610 121000 57666 121009
rect 57610 120935 57666 120944
rect 57716 115025 57744 226199
rect 57808 219337 57836 227695
rect 57886 226128 57942 226137
rect 57886 226063 57942 226072
rect 57794 219328 57850 219337
rect 57794 219263 57850 219272
rect 57900 198393 57928 226063
rect 57886 198384 57942 198393
rect 57886 198319 57942 198328
rect 57796 169720 57848 169726
rect 57796 169662 57848 169668
rect 57808 168609 57836 169662
rect 57794 168600 57850 168609
rect 57794 168535 57850 168544
rect 57796 160064 57848 160070
rect 57796 160006 57848 160012
rect 57808 159769 57836 160006
rect 57794 159760 57850 159769
rect 57794 159695 57850 159704
rect 57796 142112 57848 142118
rect 57796 142054 57848 142060
rect 57808 141817 57836 142054
rect 57794 141808 57850 141817
rect 57794 141743 57850 141752
rect 57796 137488 57848 137494
rect 57796 137430 57848 137436
rect 57808 132841 57836 137430
rect 57794 132832 57850 132841
rect 57794 132767 57850 132776
rect 58176 129849 58204 232591
rect 58162 129840 58218 129849
rect 58162 129775 58218 129784
rect 57702 115016 57758 115025
rect 57702 114951 57758 114960
rect 57612 113144 57664 113150
rect 57612 113086 57664 113092
rect 57624 112033 57652 113086
rect 57610 112024 57666 112033
rect 57610 111959 57666 111968
rect 57610 106040 57666 106049
rect 57610 105975 57666 105984
rect 57624 105602 57652 105975
rect 57612 105596 57664 105602
rect 57612 105538 57664 105544
rect 57612 103488 57664 103494
rect 57612 103430 57664 103436
rect 57624 103057 57652 103430
rect 57610 103048 57666 103057
rect 57610 102983 57666 102992
rect 57612 100700 57664 100706
rect 57612 100642 57664 100648
rect 57624 100065 57652 100642
rect 57610 100056 57666 100065
rect 57610 99991 57666 100000
rect 58268 94217 58296 236535
rect 58254 94208 58310 94217
rect 58254 94143 58310 94152
rect 57518 91216 57574 91225
rect 57518 91151 57574 91160
rect 57612 88324 57664 88330
rect 57612 88266 57664 88272
rect 57624 88233 57652 88266
rect 57610 88224 57666 88233
rect 57610 88159 57666 88168
rect 58360 85241 58388 242111
rect 58452 201385 58480 396986
rect 58532 396704 58584 396710
rect 58532 396646 58584 396652
rect 58438 201376 58494 201385
rect 58438 201311 58494 201320
rect 58544 165617 58572 396646
rect 58636 232801 58664 485007
rect 58622 232792 58678 232801
rect 58622 232727 58678 232736
rect 58622 227352 58678 227361
rect 58622 227287 58678 227296
rect 58530 165608 58586 165617
rect 58530 165543 58586 165552
rect 58346 85232 58402 85241
rect 58346 85167 58402 85176
rect 57612 70372 57664 70378
rect 57612 70314 57664 70320
rect 57624 70281 57652 70314
rect 57610 70272 57666 70281
rect 57610 70207 57666 70216
rect 57334 61432 57390 61441
rect 57334 61367 57390 61376
rect 56692 59356 56744 59362
rect 56692 59298 56744 59304
rect 56600 59288 56652 59294
rect 56600 59230 56652 59236
rect 56506 57760 56562 57769
rect 56506 57695 56562 57704
rect 56520 57361 56548 57695
rect 56506 57352 56562 57361
rect 56506 57287 56562 57296
rect 58636 57089 58664 227287
rect 58728 204377 58756 489903
rect 58820 399430 58848 700266
rect 89180 699718 89208 703520
rect 105464 699718 105492 703520
rect 137848 700330 137876 703520
rect 154132 700330 154160 703520
rect 170324 700398 170352 703520
rect 202800 703050 202828 703520
rect 201500 703044 201552 703050
rect 201500 702986 201552 702992
rect 202788 703044 202840 703050
rect 202788 702986 202840 702992
rect 198004 700800 198056 700806
rect 198004 700742 198056 700748
rect 170312 700392 170364 700398
rect 170312 700334 170364 700340
rect 196532 700392 196584 700398
rect 196532 700334 196584 700340
rect 137836 700324 137888 700330
rect 137836 700266 137888 700272
rect 146944 700324 146996 700330
rect 146944 700266 146996 700272
rect 154120 700324 154172 700330
rect 154120 700266 154172 700272
rect 88340 699712 88392 699718
rect 88340 699654 88392 699660
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 104900 699712 104952 699718
rect 104900 699654 104952 699660
rect 105452 699712 105504 699718
rect 105452 699654 105504 699660
rect 59082 490104 59138 490113
rect 59082 490039 59138 490048
rect 58990 488744 59046 488753
rect 58990 488679 59046 488688
rect 58898 488608 58954 488617
rect 58898 488543 58954 488552
rect 58808 399424 58860 399430
rect 58808 399366 58860 399372
rect 58808 396432 58860 396438
rect 58808 396374 58860 396380
rect 58714 204368 58770 204377
rect 58714 204303 58770 204312
rect 58820 97073 58848 396374
rect 58912 180577 58940 488543
rect 58898 180568 58954 180577
rect 58898 180503 58954 180512
rect 58900 175228 58952 175234
rect 58900 175170 58952 175176
rect 58806 97064 58862 97073
rect 58806 96999 58862 97008
rect 58912 57905 58940 175170
rect 59004 174593 59032 488679
rect 58990 174584 59046 174593
rect 58990 174519 59046 174528
rect 59096 124001 59124 490039
rect 59174 489016 59230 489025
rect 59174 488951 59230 488960
rect 59082 123992 59138 124001
rect 59082 123927 59138 123936
rect 59188 76265 59216 488951
rect 88352 485217 88380 699654
rect 103978 491464 104034 491473
rect 103978 491399 104034 491408
rect 101678 491328 101734 491337
rect 101678 491263 101734 491272
rect 99194 487792 99250 487801
rect 99194 487727 99250 487736
rect 99208 486033 99236 487727
rect 101692 486577 101720 491263
rect 103992 486577 104020 491399
rect 101678 486568 101734 486577
rect 101678 486503 101734 486512
rect 103978 486568 104034 486577
rect 103978 486503 104034 486512
rect 99194 486024 99250 486033
rect 99194 485959 99250 485968
rect 60002 485208 60058 485217
rect 60002 485143 60058 485152
rect 88338 485208 88394 485217
rect 88338 485143 88394 485152
rect 59266 484528 59322 484537
rect 59266 484463 59322 484472
rect 59174 76256 59230 76265
rect 59174 76191 59230 76200
rect 59280 67289 59308 484463
rect 59450 484120 59506 484129
rect 59450 484055 59506 484064
rect 59358 408232 59414 408241
rect 59358 408167 59414 408176
rect 59372 400110 59400 408167
rect 59360 400104 59412 400110
rect 59360 400046 59412 400052
rect 59372 74534 59400 400046
rect 59464 213353 59492 484055
rect 59912 396364 59964 396370
rect 59912 396306 59964 396312
rect 59544 396296 59596 396302
rect 59544 396238 59596 396244
rect 59450 213344 59506 213353
rect 59450 213279 59506 213288
rect 59556 138825 59584 396238
rect 59924 180794 59952 396306
rect 60016 229945 60044 485143
rect 104912 485081 104940 699654
rect 146956 677550 146984 700266
rect 146944 677544 146996 677550
rect 146944 677486 146996 677492
rect 153844 677544 153896 677550
rect 153844 677486 153896 677492
rect 153856 661094 153884 677486
rect 153844 661088 153896 661094
rect 153844 661030 153896 661036
rect 159364 661088 159416 661094
rect 159364 661030 159416 661036
rect 159376 652730 159404 661030
rect 159364 652724 159416 652730
rect 159364 652666 159416 652672
rect 162768 652724 162820 652730
rect 162768 652666 162820 652672
rect 162780 648922 162808 652666
rect 162768 648916 162820 648922
rect 162768 648858 162820 648864
rect 166264 648916 166316 648922
rect 166264 648858 166316 648864
rect 166276 639606 166304 648858
rect 166264 639600 166316 639606
rect 166264 639542 166316 639548
rect 175924 639600 175976 639606
rect 175924 639542 175976 639548
rect 175936 617574 175964 639542
rect 175924 617568 175976 617574
rect 175924 617510 175976 617516
rect 186964 617568 187016 617574
rect 186964 617510 187016 617516
rect 186976 597514 187004 617510
rect 186964 597508 187016 597514
rect 186964 597450 187016 597456
rect 189724 597508 189776 597514
rect 189724 597450 189776 597456
rect 189736 566506 189764 597450
rect 189724 566500 189776 566506
rect 189724 566442 189776 566448
rect 108762 490240 108818 490249
rect 108762 490175 108818 490184
rect 108776 486577 108804 490175
rect 178314 489016 178370 489025
rect 178314 488951 178370 488960
rect 130842 487928 130898 487937
rect 130842 487863 130898 487872
rect 126334 487656 126390 487665
rect 126334 487591 126390 487600
rect 126348 486713 126376 487591
rect 130856 486713 130884 487863
rect 126334 486704 126390 486713
rect 126334 486639 126390 486648
rect 130842 486704 130898 486713
rect 130842 486639 130898 486648
rect 108762 486568 108818 486577
rect 108762 486503 108818 486512
rect 178328 485625 178356 488951
rect 178314 485616 178370 485625
rect 178314 485551 178370 485560
rect 104898 485072 104954 485081
rect 104898 485007 104954 485016
rect 122748 400036 122800 400042
rect 122748 399978 122800 399984
rect 115756 399968 115808 399974
rect 115756 399910 115808 399916
rect 115664 399900 115716 399906
rect 115664 399842 115716 399848
rect 85394 398168 85450 398177
rect 85394 398103 85450 398112
rect 113638 398168 113694 398177
rect 113638 398103 113694 398112
rect 78310 397352 78366 397361
rect 61476 397316 61528 397322
rect 78310 397287 78366 397296
rect 79966 397352 80022 397361
rect 79966 397287 80022 397296
rect 80426 397352 80482 397361
rect 80426 397287 80482 397296
rect 83278 397352 83334 397361
rect 83278 397287 83334 397296
rect 61476 397258 61528 397264
rect 60002 229936 60058 229945
rect 60002 229871 60058 229880
rect 61488 229094 61516 397258
rect 61752 397180 61804 397186
rect 61752 397122 61804 397128
rect 61660 396500 61712 396506
rect 61660 396442 61712 396448
rect 61568 265736 61620 265742
rect 61568 265678 61620 265684
rect 61120 229066 61516 229094
rect 61120 226681 61148 229066
rect 61580 227066 61608 265678
rect 61672 229094 61700 396442
rect 61764 248414 61792 397122
rect 62764 397112 62816 397118
rect 62764 397054 62816 397060
rect 61764 248386 61976 248414
rect 61672 229066 61792 229094
rect 61212 227038 61608 227066
rect 61106 226672 61162 226681
rect 61106 226607 61162 226616
rect 60186 226400 60242 226409
rect 60242 226358 60490 226386
rect 60186 226335 60242 226344
rect 61106 226264 61162 226273
rect 61212 226250 61240 227038
rect 61290 226944 61346 226953
rect 61290 226879 61346 226888
rect 61304 226794 61332 226879
rect 61304 226766 61410 226794
rect 61764 226409 61792 229066
rect 61750 226400 61806 226409
rect 61750 226335 61806 226344
rect 61948 226273 61976 248386
rect 62776 227769 62804 397054
rect 78324 396982 78352 397287
rect 78312 396976 78364 396982
rect 78312 396918 78364 396924
rect 77206 396808 77262 396817
rect 77206 396743 77262 396752
rect 75918 396672 75974 396681
rect 75918 396607 75974 396616
rect 73618 234696 73674 234705
rect 73618 234631 73674 234640
rect 67546 233472 67602 233481
rect 67546 233407 67602 233416
rect 64786 233336 64842 233345
rect 64786 233271 64842 233280
rect 63406 230344 63462 230353
rect 63406 230279 63462 230288
rect 62762 227760 62818 227769
rect 62762 227695 62818 227704
rect 63420 226780 63448 230279
rect 64800 226794 64828 233271
rect 66350 229256 66406 229265
rect 66350 229191 66406 229200
rect 65338 227896 65394 227905
rect 65338 227831 65394 227840
rect 64354 226766 64828 226794
rect 65352 226780 65380 227831
rect 66364 226780 66392 229191
rect 67560 226794 67588 233407
rect 72698 232112 72754 232121
rect 72698 232047 72754 232056
rect 69294 230616 69350 230625
rect 69294 230551 69350 230560
rect 67390 226766 67588 226794
rect 69308 226780 69336 230551
rect 70306 229664 70362 229673
rect 70306 229599 70362 229608
rect 70320 228585 70348 229599
rect 70306 228576 70362 228585
rect 70306 228511 70362 228520
rect 71226 228032 71282 228041
rect 71226 227967 71282 227976
rect 70306 227760 70362 227769
rect 70306 227695 70362 227704
rect 70320 226780 70348 227695
rect 71240 226780 71268 227967
rect 72712 226794 72740 232047
rect 73632 226794 73660 234631
rect 74538 229800 74594 229809
rect 74538 229735 74594 229744
rect 74262 228168 74318 228177
rect 74262 228103 74318 228112
rect 72266 226766 72740 226794
rect 73278 226766 73660 226794
rect 74276 226780 74304 228103
rect 74552 227225 74580 229735
rect 75932 227361 75960 396607
rect 77220 265946 77248 396743
rect 79980 396574 80008 397287
rect 79968 396568 80020 396574
rect 79968 396510 80020 396516
rect 80440 396370 80468 397287
rect 83292 397254 83320 397287
rect 83280 397248 83332 397254
rect 83280 397190 83332 397196
rect 82726 396808 82782 396817
rect 82726 396743 82782 396752
rect 80428 396364 80480 396370
rect 80428 396306 80480 396312
rect 82636 324352 82688 324358
rect 82636 324294 82688 324300
rect 81348 298172 81400 298178
rect 81348 298114 81400 298120
rect 79968 271924 80020 271930
rect 79968 271866 80020 271872
rect 77208 265940 77260 265946
rect 77208 265882 77260 265888
rect 78586 247072 78642 247081
rect 78586 247007 78642 247016
rect 76562 234832 76618 234841
rect 76562 234767 76618 234776
rect 75918 227352 75974 227361
rect 75918 227287 75974 227296
rect 74538 227216 74594 227225
rect 74538 227151 74594 227160
rect 76576 226794 76604 234767
rect 78600 226794 78628 247007
rect 79980 229094 80008 271866
rect 80610 236328 80666 236337
rect 80610 236263 80666 236272
rect 79520 229066 80008 229094
rect 79520 226794 79548 229066
rect 80624 226794 80652 236263
rect 81360 226794 81388 298114
rect 82648 229094 82676 324294
rect 82740 266014 82768 396743
rect 85408 378826 85436 398103
rect 87696 397384 87748 397390
rect 86498 397352 86554 397361
rect 86498 397287 86554 397296
rect 87694 397352 87696 397361
rect 87748 397352 87750 397361
rect 87694 397287 87750 397296
rect 88706 397352 88762 397361
rect 88706 397287 88762 397296
rect 92294 397352 92350 397361
rect 92294 397287 92350 397296
rect 93490 397352 93546 397361
rect 93490 397287 93546 397296
rect 96526 397352 96582 397361
rect 96526 397287 96582 397296
rect 98918 397352 98974 397361
rect 98918 397287 98974 397296
rect 100114 397352 100170 397361
rect 100114 397287 100170 397296
rect 101586 397352 101642 397361
rect 101586 397287 101642 397296
rect 101862 397352 101918 397361
rect 101862 397287 101918 397296
rect 102874 397352 102930 397361
rect 102874 397287 102930 397296
rect 103702 397352 103758 397361
rect 103702 397287 103758 397296
rect 105910 397352 105966 397361
rect 105910 397287 105966 397296
rect 107198 397352 107254 397361
rect 107198 397287 107254 397296
rect 109774 397352 109830 397361
rect 109774 397287 109830 397296
rect 111614 397352 111670 397361
rect 111614 397287 111670 397296
rect 85486 396808 85542 396817
rect 85486 396743 85542 396752
rect 85396 378820 85448 378826
rect 85396 378762 85448 378768
rect 85396 378208 85448 378214
rect 85396 378150 85448 378156
rect 84108 351960 84160 351966
rect 84108 351902 84160 351908
rect 84016 311908 84068 311914
rect 84016 311850 84068 311856
rect 82728 266008 82780 266014
rect 82728 265950 82780 265956
rect 84028 229094 84056 311850
rect 82464 229066 82676 229094
rect 83568 229066 84056 229094
rect 82464 226794 82492 229066
rect 83568 226794 83596 229066
rect 76222 226766 76604 226794
rect 78246 226766 78628 226794
rect 79166 226766 79548 226794
rect 80178 226766 80652 226794
rect 81190 226766 81388 226794
rect 82110 226766 82492 226794
rect 83122 226766 83596 226794
rect 84120 226780 84148 351902
rect 85408 226794 85436 378150
rect 85500 232529 85528 396743
rect 86512 396438 86540 397287
rect 88720 396506 88748 397287
rect 92308 396914 92336 397287
rect 92296 396908 92348 396914
rect 92296 396850 92348 396856
rect 93504 396846 93532 397287
rect 96434 397216 96490 397225
rect 96434 397151 96490 397160
rect 93492 396840 93544 396846
rect 89626 396808 89682 396817
rect 89626 396743 89682 396752
rect 91006 396808 91062 396817
rect 93492 396782 93544 396788
rect 93766 396808 93822 396817
rect 91006 396743 91062 396752
rect 93766 396743 93822 396752
rect 95146 396808 95202 396817
rect 95146 396743 95202 396752
rect 88708 396500 88760 396506
rect 88708 396442 88760 396448
rect 86500 396432 86552 396438
rect 86500 396374 86552 396380
rect 86868 364404 86920 364410
rect 86868 364346 86920 364352
rect 86222 257952 86278 257961
rect 86222 257887 86278 257896
rect 86236 236337 86264 257887
rect 86222 236328 86278 236337
rect 86222 236263 86278 236272
rect 85486 232520 85542 232529
rect 85486 232455 85542 232464
rect 86880 229094 86908 364346
rect 89536 264240 89588 264246
rect 89536 264182 89588 264188
rect 88248 262880 88300 262886
rect 88248 262822 88300 262828
rect 88156 261588 88208 261594
rect 88156 261530 88208 261536
rect 88168 229094 88196 261530
rect 86512 229066 86908 229094
rect 87432 229066 88196 229094
rect 86512 226794 86540 229066
rect 87432 226794 87460 229066
rect 88260 226794 88288 262822
rect 89548 229094 89576 264182
rect 89640 260438 89668 396743
rect 89718 396672 89774 396681
rect 89718 396607 89774 396616
rect 89628 260432 89680 260438
rect 89628 260374 89680 260380
rect 89732 260234 89760 396607
rect 91020 264518 91048 396743
rect 91098 396672 91154 396681
rect 91098 396607 91154 396616
rect 91008 264512 91060 264518
rect 91008 264454 91060 264460
rect 91008 261656 91060 261662
rect 91008 261598 91060 261604
rect 89720 260228 89772 260234
rect 89720 260170 89772 260176
rect 90916 260228 90968 260234
rect 90916 260170 90968 260176
rect 90928 229094 90956 260170
rect 89456 229066 89576 229094
rect 90376 229066 90956 229094
rect 89456 226794 89484 229066
rect 90376 226794 90404 229066
rect 85146 226766 85436 226794
rect 86066 226766 86540 226794
rect 87078 226766 87460 226794
rect 88090 226766 88288 226794
rect 89102 226766 89484 226794
rect 90022 226766 90404 226794
rect 91020 226780 91048 261598
rect 91112 232665 91140 396607
rect 93780 264654 93808 396743
rect 95056 298784 95108 298790
rect 95056 298726 95108 298732
rect 93768 264648 93820 264654
rect 93768 264590 93820 264596
rect 92388 262948 92440 262954
rect 92388 262890 92440 262896
rect 91098 232656 91154 232665
rect 91098 232591 91154 232600
rect 92400 226794 92428 262890
rect 93768 260364 93820 260370
rect 93768 260306 93820 260312
rect 93780 229094 93808 260306
rect 95068 229094 95096 298726
rect 95160 264586 95188 396743
rect 96448 395554 96476 397151
rect 96540 396098 96568 397287
rect 98458 397216 98514 397225
rect 98458 397151 98514 397160
rect 97906 396808 97962 396817
rect 97906 396743 97962 396752
rect 96528 396092 96580 396098
rect 96528 396034 96580 396040
rect 96436 395548 96488 395554
rect 96436 395490 96488 395496
rect 97816 300144 97868 300150
rect 97816 300086 97868 300092
rect 95148 264580 95200 264586
rect 95148 264522 95200 264528
rect 95148 263016 95200 263022
rect 95148 262958 95200 262964
rect 93320 229066 93808 229094
rect 94424 229066 95096 229094
rect 93320 226794 93348 229066
rect 94424 226794 94452 229066
rect 95160 226794 95188 262958
rect 96528 260296 96580 260302
rect 96528 260238 96580 260244
rect 96540 229094 96568 260238
rect 97828 229094 97856 300086
rect 97920 264722 97948 396743
rect 98472 395622 98500 397151
rect 98644 396568 98696 396574
rect 98644 396510 98696 396516
rect 98460 395616 98512 395622
rect 98460 395558 98512 395564
rect 98656 267034 98684 396510
rect 98932 396506 98960 397287
rect 100128 396574 100156 397287
rect 100116 396568 100168 396574
rect 100116 396510 100168 396516
rect 98920 396500 98972 396506
rect 98920 396442 98972 396448
rect 101600 396370 101628 397287
rect 101876 396642 101904 397287
rect 101954 396808 102010 396817
rect 101954 396743 102010 396752
rect 101864 396636 101916 396642
rect 101864 396578 101916 396584
rect 101588 396364 101640 396370
rect 101588 396306 101640 396312
rect 98644 267028 98696 267034
rect 98644 266970 98696 266976
rect 101968 266150 101996 396743
rect 102888 396234 102916 397287
rect 103716 396710 103744 397287
rect 104806 397216 104862 397225
rect 104806 397151 104862 397160
rect 103704 396704 103756 396710
rect 103704 396646 103756 396652
rect 102876 396228 102928 396234
rect 102876 396170 102928 396176
rect 101956 266144 102008 266150
rect 101956 266086 102008 266092
rect 97908 264716 97960 264722
rect 97908 264658 97960 264664
rect 102048 263220 102100 263226
rect 102048 263162 102100 263168
rect 97908 263084 97960 263090
rect 97908 263026 97960 263032
rect 96448 229066 96568 229094
rect 97368 229066 97856 229094
rect 96448 226794 96476 229066
rect 97368 226794 97396 229066
rect 92046 226766 92428 226794
rect 92966 226766 93348 226794
rect 93978 226766 94452 226794
rect 94990 226766 95188 226794
rect 96002 226766 96476 226794
rect 96922 226766 97396 226794
rect 97920 226780 97948 263026
rect 99288 261928 99340 261934
rect 99288 261870 99340 261876
rect 99300 226794 99328 261870
rect 100668 261860 100720 261866
rect 100668 261802 100720 261808
rect 100680 229094 100708 261802
rect 101956 260772 102008 260778
rect 101956 260714 102008 260720
rect 101126 233880 101182 233889
rect 101126 233815 101182 233824
rect 100312 229066 100708 229094
rect 100312 226794 100340 229066
rect 101140 226794 101168 233815
rect 101968 226794 101996 260714
rect 102060 233889 102088 263162
rect 104716 263152 104768 263158
rect 104716 263094 104768 263100
rect 103428 261724 103480 261730
rect 103428 261666 103480 261672
rect 102046 233880 102102 233889
rect 102046 233815 102102 233824
rect 103440 229094 103468 261666
rect 104624 261248 104676 261254
rect 104624 261190 104676 261196
rect 104070 233880 104126 233889
rect 104070 233815 104126 233824
rect 103256 229066 103468 229094
rect 103256 226794 103284 229066
rect 104084 226794 104112 233815
rect 98946 226766 99328 226794
rect 99866 226766 100340 226794
rect 100878 226766 101168 226794
rect 101890 226766 101996 226794
rect 102902 226766 103284 226794
rect 103822 226766 104112 226794
rect 104636 226794 104664 261190
rect 104728 233889 104756 263094
rect 104820 238105 104848 397151
rect 105924 396710 105952 397287
rect 106002 396808 106058 396817
rect 106002 396743 106058 396752
rect 105912 396704 105964 396710
rect 105912 396646 105964 396652
rect 104806 238096 104862 238105
rect 104806 238031 104862 238040
rect 104714 233880 104770 233889
rect 104714 233815 104770 233824
rect 106016 232665 106044 396743
rect 107016 396228 107068 396234
rect 107016 396170 107068 396176
rect 106924 396092 106976 396098
rect 106924 396034 106976 396040
rect 106936 264042 106964 396034
rect 107028 266218 107056 396170
rect 107212 396098 107240 397287
rect 107382 396808 107438 396817
rect 107382 396743 107438 396752
rect 108854 396808 108910 396817
rect 109788 396778 109816 397287
rect 111522 396808 111578 396817
rect 108854 396743 108910 396752
rect 109776 396772 109828 396778
rect 107200 396092 107252 396098
rect 107200 396034 107252 396040
rect 107016 266212 107068 266218
rect 107016 266154 107068 266160
rect 107396 266082 107424 396743
rect 107476 294636 107528 294642
rect 107476 294578 107528 294584
rect 107384 266076 107436 266082
rect 107384 266018 107436 266024
rect 106924 264036 106976 264042
rect 106924 263978 106976 263984
rect 106096 261792 106148 261798
rect 106096 261734 106148 261740
rect 106002 232656 106058 232665
rect 106002 232591 106058 232600
rect 106108 226794 106136 261734
rect 107488 229094 107516 294578
rect 108868 263430 108896 396743
rect 111522 396743 111578 396752
rect 109776 396714 109828 396720
rect 108946 396672 109002 396681
rect 108946 396607 109002 396616
rect 108856 263424 108908 263430
rect 108856 263366 108908 263372
rect 108856 263288 108908 263294
rect 108856 263230 108908 263236
rect 108764 261996 108816 262002
rect 108764 261938 108816 261944
rect 108776 229094 108804 261938
rect 107304 229066 107516 229094
rect 108224 229066 108804 229094
rect 107304 226794 107332 229066
rect 108224 226794 108252 229066
rect 108868 226794 108896 263230
rect 108960 244905 108988 396607
rect 111536 265538 111564 396743
rect 111628 396166 111656 397287
rect 113178 397216 113234 397225
rect 113178 397151 113234 397160
rect 113192 397050 113220 397151
rect 113180 397044 113232 397050
rect 113180 396986 113232 396992
rect 113086 396808 113142 396817
rect 113086 396743 113142 396752
rect 112444 396364 112496 396370
rect 112444 396306 112496 396312
rect 111616 396160 111668 396166
rect 111616 396102 111668 396108
rect 111616 284980 111668 284986
rect 111616 284922 111668 284928
rect 111524 265532 111576 265538
rect 111524 265474 111576 265480
rect 110328 261520 110380 261526
rect 110328 261462 110380 261468
rect 108946 244896 109002 244905
rect 108946 244831 109002 244840
rect 110340 229094 110368 261462
rect 111628 229094 111656 284922
rect 112456 266354 112484 396306
rect 112996 294704 113048 294710
rect 112996 294646 113048 294652
rect 112444 266348 112496 266354
rect 112444 266290 112496 266296
rect 111708 263356 111760 263362
rect 111708 263298 111760 263304
rect 110248 229066 110368 229094
rect 111168 229066 111656 229094
rect 110248 226794 110276 229066
rect 111168 226794 111196 229066
rect 104636 226766 104834 226794
rect 105846 226766 106136 226794
rect 106858 226766 107332 226794
rect 107778 226766 108252 226794
rect 108790 226766 108896 226794
rect 109802 226766 110276 226794
rect 110722 226766 111196 226794
rect 111720 226780 111748 263298
rect 113008 226794 113036 294646
rect 113100 243545 113128 396743
rect 113652 395894 113680 398103
rect 114466 397352 114522 397361
rect 114466 397287 114522 397296
rect 114480 397050 114508 397287
rect 114468 397044 114520 397050
rect 114468 396986 114520 396992
rect 113640 395888 113692 395894
rect 113640 395830 113692 395836
rect 115676 393314 115704 399842
rect 115768 395434 115796 399910
rect 119988 398132 120040 398138
rect 119988 398074 120040 398080
rect 115846 397352 115902 397361
rect 115846 397287 115902 397296
rect 118146 397352 118202 397361
rect 118146 397287 118202 397296
rect 115860 395622 115888 397287
rect 117226 396808 117282 396817
rect 117226 396743 117282 396752
rect 117134 396672 117190 396681
rect 117134 396607 117190 396616
rect 116584 396092 116636 396098
rect 116584 396034 116636 396040
rect 115848 395616 115900 395622
rect 115848 395558 115900 395564
rect 115768 395406 115888 395434
rect 115676 393286 115796 393314
rect 114468 260840 114520 260846
rect 114468 260782 114520 260788
rect 113086 243536 113142 243545
rect 113086 243471 113142 243480
rect 114480 229094 114508 260782
rect 114926 233880 114982 233889
rect 114926 233815 114982 233824
rect 114112 229066 114508 229094
rect 114112 226794 114140 229066
rect 114940 226794 114968 233815
rect 115768 226794 115796 393286
rect 115860 233889 115888 395406
rect 116596 266286 116624 396034
rect 116584 266280 116636 266286
rect 116584 266222 116636 266228
rect 117148 261322 117176 396607
rect 117136 261316 117188 261322
rect 117136 261258 117188 261264
rect 117136 261112 117188 261118
rect 117136 261054 117188 261060
rect 115846 233880 115902 233889
rect 115846 233815 115902 233824
rect 117148 229094 117176 261054
rect 117240 242321 117268 396743
rect 118160 395758 118188 397287
rect 118606 396808 118662 396817
rect 118606 396743 118662 396752
rect 119894 396808 119950 396817
rect 119894 396743 119950 396752
rect 118148 395752 118200 395758
rect 118148 395694 118200 395700
rect 118516 262472 118568 262478
rect 118516 262414 118568 262420
rect 118424 260092 118476 260098
rect 118424 260034 118476 260040
rect 117226 242312 117282 242321
rect 117226 242247 117282 242256
rect 118436 229094 118464 260034
rect 117056 229066 117176 229094
rect 118160 229066 118464 229094
rect 117056 226794 117084 229066
rect 118160 226794 118188 229066
rect 112746 226766 113036 226794
rect 113758 226766 114140 226794
rect 114678 226766 114968 226794
rect 115690 226766 115796 226794
rect 116702 226766 117084 226794
rect 117714 226766 118188 226794
rect 118528 226794 118556 262414
rect 118620 249257 118648 396743
rect 119344 396160 119396 396166
rect 119344 396102 119396 396108
rect 119356 264110 119384 396102
rect 119908 358086 119936 396743
rect 119896 358080 119948 358086
rect 119896 358022 119948 358028
rect 119344 264104 119396 264110
rect 119344 264046 119396 264052
rect 118606 249248 118662 249257
rect 118606 249183 118662 249192
rect 120000 226794 120028 398074
rect 121366 396808 121422 396817
rect 121366 396743 121422 396752
rect 121276 260976 121328 260982
rect 121276 260918 121328 260924
rect 121288 229094 121316 260918
rect 121380 260710 121408 396743
rect 121368 260704 121420 260710
rect 121368 260646 121420 260652
rect 122760 238754 122788 399978
rect 172520 399696 172572 399702
rect 172520 399638 172572 399644
rect 187608 399696 187660 399702
rect 187608 399638 187660 399644
rect 125600 399424 125652 399430
rect 125600 399366 125652 399372
rect 125508 398200 125560 398206
rect 125508 398142 125560 398148
rect 124126 396808 124182 396817
rect 124126 396743 124182 396752
rect 124140 250481 124168 396743
rect 124126 250472 124182 250481
rect 124126 250407 124182 250416
rect 124126 240816 124182 240825
rect 124126 240751 124182 240760
rect 121104 229066 121316 229094
rect 121932 238726 122788 238754
rect 121104 226794 121132 229066
rect 121932 226794 121960 238726
rect 122654 236736 122710 236745
rect 122654 236671 122710 236680
rect 122668 226794 122696 236671
rect 124140 229094 124168 240751
rect 125520 238754 125548 398142
rect 125612 248414 125640 399366
rect 146300 397520 146352 397526
rect 146300 397462 146352 397468
rect 136454 397352 136510 397361
rect 136454 397287 136510 397296
rect 138478 397352 138534 397361
rect 138478 397287 138534 397296
rect 126886 396808 126942 396817
rect 126886 396743 126942 396752
rect 129646 396808 129702 396817
rect 129646 396743 129702 396752
rect 131026 396808 131082 396817
rect 131026 396743 131082 396752
rect 133786 396808 133842 396817
rect 133786 396743 133842 396752
rect 126900 263906 126928 396743
rect 126888 263900 126940 263906
rect 126888 263842 126940 263848
rect 128360 263492 128412 263498
rect 128360 263434 128412 263440
rect 125612 248386 126192 248414
rect 124048 229066 124168 229094
rect 124968 238726 125548 238754
rect 124048 226794 124076 229066
rect 124968 226794 124996 238726
rect 125138 232792 125194 232801
rect 125138 232727 125194 232736
rect 118528 226766 118634 226794
rect 119646 226766 120028 226794
rect 120658 226766 121132 226794
rect 121578 226766 121960 226794
rect 122590 226766 122696 226794
rect 123602 226766 124076 226794
rect 124614 226766 124996 226794
rect 125152 226794 125180 232727
rect 126164 226794 126192 248386
rect 128372 230489 128400 263434
rect 129660 262410 129688 396743
rect 131040 319462 131068 396743
rect 131028 319456 131080 319462
rect 131028 319398 131080 319404
rect 133800 264178 133828 396743
rect 136468 395758 136496 397287
rect 137284 397044 137336 397050
rect 137284 396986 137336 396992
rect 136456 395752 136508 395758
rect 136456 395694 136508 395700
rect 133880 290488 133932 290494
rect 133880 290430 133932 290436
rect 132500 264172 132552 264178
rect 132500 264114 132552 264120
rect 133788 264172 133840 264178
rect 133788 264114 133840 264120
rect 129740 262608 129792 262614
rect 129740 262550 129792 262556
rect 129648 262404 129700 262410
rect 129648 262346 129700 262352
rect 128452 261044 128504 261050
rect 128452 260986 128504 260992
rect 128358 230480 128414 230489
rect 128358 230415 128414 230424
rect 127530 229936 127586 229945
rect 127530 229871 127586 229880
rect 125152 226766 125534 226794
rect 126164 226766 126546 226794
rect 127544 226780 127572 229871
rect 128464 226780 128492 260986
rect 129752 248414 129780 262550
rect 131120 260568 131172 260574
rect 131120 260510 131172 260516
rect 129752 248386 130056 248414
rect 129186 230480 129242 230489
rect 129186 230415 129242 230424
rect 129200 226794 129228 230415
rect 130028 226794 130056 248386
rect 131132 230489 131160 260510
rect 131212 260500 131264 260506
rect 131212 260442 131264 260448
rect 131118 230480 131174 230489
rect 131118 230415 131174 230424
rect 131224 226794 131252 260442
rect 132512 248414 132540 264114
rect 133892 248414 133920 290430
rect 137296 265606 137324 396986
rect 138492 395826 138520 397287
rect 140778 396808 140834 396817
rect 140778 396743 140834 396752
rect 144826 396808 144882 396817
rect 144826 396743 144882 396752
rect 146206 396808 146262 396817
rect 146206 396743 146262 396752
rect 138480 395820 138532 395826
rect 138480 395762 138532 395768
rect 137284 265600 137336 265606
rect 137284 265542 137336 265548
rect 140792 263974 140820 396743
rect 142160 297424 142212 297430
rect 142160 297366 142212 297372
rect 140780 263968 140832 263974
rect 140780 263910 140832 263916
rect 140780 263560 140832 263566
rect 140780 263502 140832 263508
rect 138020 262744 138072 262750
rect 138020 262686 138072 262692
rect 135260 262676 135312 262682
rect 135260 262618 135312 262624
rect 132512 248386 133000 248414
rect 133892 248386 134104 248414
rect 132130 230480 132186 230489
rect 132130 230415 132186 230424
rect 132144 226794 132172 230415
rect 132972 226794 133000 248386
rect 134076 226794 134104 248386
rect 135272 230489 135300 262618
rect 136640 262200 136692 262206
rect 136640 262142 136692 262148
rect 135352 261384 135404 261390
rect 135352 261326 135404 261332
rect 135364 234614 135392 261326
rect 136652 248414 136680 262142
rect 136652 248386 137048 248414
rect 135364 234586 135484 234614
rect 135258 230480 135314 230489
rect 135258 230415 135314 230424
rect 129200 226766 129490 226794
rect 130028 226766 130502 226794
rect 131224 226766 131514 226794
rect 132144 226766 132434 226794
rect 132972 226766 133446 226794
rect 134076 226766 134458 226794
rect 135456 226780 135484 234586
rect 135994 230480 136050 230489
rect 135994 230415 136050 230424
rect 136008 226794 136036 230415
rect 137020 226794 137048 248386
rect 138032 230489 138060 262686
rect 139400 261452 139452 261458
rect 139400 261394 139452 261400
rect 138112 260636 138164 260642
rect 138112 260578 138164 260584
rect 138018 230480 138074 230489
rect 138018 230415 138074 230424
rect 138124 226794 138152 260578
rect 139412 248414 139440 261394
rect 140792 248414 140820 263502
rect 141422 255912 141478 255921
rect 141422 255847 141478 255856
rect 139412 248386 139992 248414
rect 140792 248386 140912 248414
rect 138202 245712 138258 245721
rect 138202 245647 138258 245656
rect 138216 240825 138244 245647
rect 138202 240816 138258 240825
rect 138202 240751 138258 240760
rect 138938 230480 138994 230489
rect 138938 230415 138994 230424
rect 138952 226794 138980 230415
rect 139964 226794 139992 248386
rect 140884 226794 140912 248386
rect 141436 245721 141464 255847
rect 141422 245712 141478 245721
rect 141422 245647 141478 245656
rect 142172 230489 142200 297366
rect 144840 269822 144868 396743
rect 144828 269816 144880 269822
rect 144828 269758 144880 269764
rect 144920 264852 144972 264858
rect 144920 264794 144972 264800
rect 142252 264784 142304 264790
rect 142252 264726 142304 264732
rect 142158 230480 142214 230489
rect 142158 230415 142214 230424
rect 142264 226794 142292 264726
rect 143540 262812 143592 262818
rect 143540 262754 143592 262760
rect 143552 248414 143580 262754
rect 143552 248386 143856 248414
rect 142986 230480 143042 230489
rect 142986 230415 143042 230424
rect 143000 226794 143028 230415
rect 143828 226794 143856 248386
rect 144932 226794 144960 264794
rect 146220 232801 146248 396743
rect 146206 232792 146262 232801
rect 146206 232727 146262 232736
rect 146312 230489 146340 397462
rect 150714 397352 150770 397361
rect 150714 397287 150770 397296
rect 147678 396808 147734 396817
rect 147678 396743 147734 396752
rect 147692 262546 147720 396743
rect 150728 395690 150756 397287
rect 170404 396976 170456 396982
rect 170404 396918 170456 396924
rect 154486 396808 154542 396817
rect 154486 396743 154542 396752
rect 155958 396808 156014 396817
rect 155958 396743 156014 396752
rect 158626 396808 158682 396817
rect 158626 396743 158682 396752
rect 161386 396808 161442 396817
rect 161386 396743 161442 396752
rect 164146 396808 164202 396817
rect 164146 396743 164202 396752
rect 166906 396808 166962 396817
rect 166906 396743 166962 396752
rect 150716 395684 150768 395690
rect 150716 395626 150768 395632
rect 149060 371272 149112 371278
rect 149060 371214 149112 371220
rect 147772 264920 147824 264926
rect 147772 264862 147824 264868
rect 147680 262540 147732 262546
rect 147680 262482 147732 262488
rect 146944 262200 146996 262206
rect 146944 262142 146996 262148
rect 146392 262132 146444 262138
rect 146392 262074 146444 262080
rect 146404 234614 146432 262074
rect 146956 255921 146984 262142
rect 146942 255912 146998 255921
rect 146942 255847 146998 255856
rect 147784 248414 147812 264862
rect 147784 248386 147904 248414
rect 146404 234586 146524 234614
rect 146298 230480 146354 230489
rect 146298 230415 146354 230424
rect 146496 226794 146524 234586
rect 146850 230480 146906 230489
rect 146850 230415 146906 230424
rect 136008 226766 136390 226794
rect 137020 226766 137402 226794
rect 138124 226766 138414 226794
rect 138952 226766 139334 226794
rect 139964 226766 140346 226794
rect 140884 226766 141358 226794
rect 142264 226766 142370 226794
rect 143000 226766 143290 226794
rect 143828 226766 144302 226794
rect 144932 226766 145314 226794
rect 146326 226766 146524 226794
rect 146864 226794 146892 230415
rect 147876 226794 147904 248386
rect 149072 226794 149100 371214
rect 150440 357468 150492 357474
rect 150440 357410 150492 357416
rect 149152 345092 149204 345098
rect 149152 345034 149204 345040
rect 149164 248414 149192 345034
rect 149244 263628 149296 263634
rect 149244 263570 149296 263576
rect 149256 262206 149284 263570
rect 149244 262200 149296 262206
rect 149244 262142 149296 262148
rect 150452 248414 150480 357410
rect 151820 318844 151872 318850
rect 151820 318786 151872 318792
rect 150532 269136 150584 269142
rect 150532 269078 150584 269084
rect 150544 263634 150572 269078
rect 150532 263628 150584 263634
rect 150532 263570 150584 263576
rect 149164 248386 149744 248414
rect 150452 248386 150848 248414
rect 149716 226794 149744 248386
rect 150820 226794 150848 248386
rect 151832 226794 151860 318786
rect 154500 305658 154528 396743
rect 155224 320476 155276 320482
rect 155224 320418 155276 320424
rect 154488 305652 154540 305658
rect 154488 305594 154540 305600
rect 153200 305040 153252 305046
rect 153200 304982 153252 304988
rect 152832 276072 152884 276078
rect 152832 276014 152884 276020
rect 152844 269142 152872 276014
rect 152832 269136 152884 269142
rect 152832 269078 152884 269084
rect 153212 230489 153240 304982
rect 155236 301578 155264 320418
rect 153844 301572 153896 301578
rect 153844 301514 153896 301520
rect 155224 301572 155276 301578
rect 155224 301514 155276 301520
rect 153292 292596 153344 292602
rect 153292 292538 153344 292544
rect 153198 230480 153254 230489
rect 153198 230415 153254 230424
rect 153304 226794 153332 292538
rect 153856 276078 153884 301514
rect 153844 276072 153896 276078
rect 153844 276014 153896 276020
rect 154580 266416 154632 266422
rect 154580 266358 154632 266364
rect 154592 248414 154620 266358
rect 155972 261186 156000 396743
rect 156604 331220 156656 331226
rect 156604 331162 156656 331168
rect 156616 320482 156644 331162
rect 156604 320476 156656 320482
rect 156604 320418 156656 320424
rect 155960 261180 156012 261186
rect 155960 261122 156012 261128
rect 155958 249112 156014 249121
rect 155958 249047 156014 249056
rect 155972 248414 156000 249047
rect 154592 248386 154712 248414
rect 155972 248386 156828 248414
rect 153842 230480 153898 230489
rect 153842 230415 153898 230424
rect 146864 226766 147246 226794
rect 147876 226766 148258 226794
rect 149072 226766 149270 226794
rect 149716 226766 150190 226794
rect 150820 226766 151202 226794
rect 151832 226766 152214 226794
rect 153226 226766 153332 226794
rect 153856 226794 153884 230415
rect 154684 226794 154712 248386
rect 156050 235240 156106 235249
rect 156050 235175 156106 235184
rect 156064 226794 156092 235175
rect 156800 226794 156828 248386
rect 158640 240825 158668 396743
rect 161400 261458 161428 396743
rect 162860 338088 162912 338094
rect 162860 338030 162912 338036
rect 162872 331294 162900 338030
rect 162860 331288 162912 331294
rect 162860 331230 162912 331236
rect 164160 264790 164188 396743
rect 166724 340944 166776 340950
rect 166724 340886 166776 340892
rect 166736 338162 166764 340886
rect 166724 338156 166776 338162
rect 166724 338098 166776 338104
rect 164148 264784 164200 264790
rect 164148 264726 164200 264732
rect 161388 261452 161440 261458
rect 161388 261394 161440 261400
rect 166920 260642 166948 396743
rect 170416 262138 170444 396918
rect 171784 358556 171836 358562
rect 171784 358498 171836 358504
rect 171796 352102 171824 358498
rect 170496 352096 170548 352102
rect 170496 352038 170548 352044
rect 171784 352096 171836 352102
rect 171784 352038 171836 352044
rect 170508 340950 170536 352038
rect 170496 340944 170548 340950
rect 170496 340886 170548 340892
rect 170404 262132 170456 262138
rect 170404 262074 170456 262080
rect 166908 260636 166960 260642
rect 166908 260578 166960 260584
rect 158626 240816 158682 240825
rect 158626 240751 158682 240760
rect 164606 233744 164662 233753
rect 164606 233679 164662 233688
rect 161662 233608 161718 233617
rect 161662 233543 161718 233552
rect 161018 231024 161074 231033
rect 161018 230959 161074 230968
rect 158074 230888 158130 230897
rect 158074 230823 158130 230832
rect 153856 226766 154146 226794
rect 154684 226766 155158 226794
rect 156064 226766 156170 226794
rect 156800 226766 157182 226794
rect 158088 226780 158116 230823
rect 160190 229800 160246 229809
rect 160190 229735 160246 229744
rect 160098 229664 160154 229673
rect 160098 229599 160154 229608
rect 160112 228313 160140 229599
rect 160098 228304 160154 228313
rect 160098 228239 160154 228248
rect 158810 226808 158866 226817
rect 160204 226794 160232 229735
rect 158866 226766 159114 226794
rect 160126 226766 160232 226794
rect 161032 226780 161060 230959
rect 161676 226794 161704 233543
rect 164054 231160 164110 231169
rect 164054 231095 164110 231104
rect 163042 229936 163098 229945
rect 163042 229871 163098 229880
rect 161676 226766 162058 226794
rect 163056 226780 163084 229871
rect 164068 226780 164096 231095
rect 164620 226794 164648 233679
rect 166998 231976 167054 231985
rect 166998 231911 167054 231920
rect 165986 229528 166042 229537
rect 165986 229463 166042 229472
rect 164620 226766 165002 226794
rect 166000 226780 166028 229463
rect 167012 226780 167040 231911
rect 169942 230752 169998 230761
rect 169942 230687 169998 230696
rect 167918 229664 167974 229673
rect 167918 229599 167974 229608
rect 167932 226780 167960 229599
rect 168562 227080 168618 227089
rect 168562 227015 168618 227024
rect 168576 226794 168604 227015
rect 168576 226766 168958 226794
rect 169956 226780 169984 230687
rect 171874 229392 171930 229401
rect 171874 229327 171930 229336
rect 170954 228440 171010 228449
rect 170954 228375 171010 228384
rect 170968 226780 170996 228375
rect 171888 226780 171916 229327
rect 172532 226794 172560 399638
rect 175188 398268 175240 398274
rect 175188 398210 175240 398216
rect 173440 360188 173492 360194
rect 173440 360130 173492 360136
rect 173452 358562 173480 360130
rect 173440 358556 173492 358562
rect 173440 358498 173492 358504
rect 173900 262132 173952 262138
rect 173900 262074 173952 262080
rect 173912 248414 173940 262074
rect 173912 248386 174584 248414
rect 174174 233880 174230 233889
rect 174174 233815 174230 233824
rect 174188 226794 174216 233815
rect 172532 226766 172914 226794
rect 173926 226766 174216 226794
rect 174556 226794 174584 248386
rect 175200 233889 175228 398210
rect 183466 397352 183522 397361
rect 183466 397287 183522 397296
rect 183480 396982 183508 397287
rect 183468 396976 183520 396982
rect 183468 396918 183520 396924
rect 183190 396808 183246 396817
rect 183190 396743 183246 396752
rect 183204 396030 183232 396743
rect 183192 396024 183244 396030
rect 183192 395966 183244 395972
rect 179328 395956 179380 395962
rect 179328 395898 179380 395904
rect 177948 395684 178000 395690
rect 177948 395626 178000 395632
rect 177304 374672 177356 374678
rect 177304 374614 177356 374620
rect 177316 360262 177344 374614
rect 177304 360256 177356 360262
rect 177304 360198 177356 360204
rect 176568 267096 176620 267102
rect 176568 267038 176620 267044
rect 175186 233880 175242 233889
rect 175186 233815 175242 233824
rect 176580 229094 176608 267038
rect 176660 267028 176712 267034
rect 176660 266970 176712 266976
rect 176304 229066 176608 229094
rect 176304 226794 176332 229066
rect 174556 226766 174938 226794
rect 175858 226766 176332 226794
rect 176672 226794 176700 266970
rect 177960 226794 177988 395626
rect 179340 229094 179368 395898
rect 186320 387864 186372 387870
rect 186320 387806 186372 387812
rect 186332 385694 186360 387806
rect 185676 385688 185728 385694
rect 185676 385630 185728 385636
rect 186320 385688 186372 385694
rect 186320 385630 186372 385636
rect 185688 379574 185716 385630
rect 183560 379568 183612 379574
rect 183560 379510 183612 379516
rect 185676 379568 185728 379574
rect 185676 379510 185728 379516
rect 183572 374678 183600 379510
rect 183560 374672 183612 374678
rect 183560 374614 183612 374620
rect 182088 267028 182140 267034
rect 182088 266970 182140 266976
rect 181996 263492 182048 263498
rect 181996 263434 182048 263440
rect 179786 229800 179842 229809
rect 179786 229735 179842 229744
rect 179248 229066 179368 229094
rect 179248 226794 179276 229066
rect 176672 226766 176870 226794
rect 177882 226766 177988 226794
rect 178802 226766 179276 226794
rect 179800 226780 179828 229735
rect 181166 226808 181222 226817
rect 180826 226766 181166 226794
rect 158810 226743 158866 226752
rect 182008 226794 182036 263434
rect 182100 226817 182128 266970
rect 186228 261384 186280 261390
rect 186228 261326 186280 261332
rect 183742 230208 183798 230217
rect 183742 230143 183798 230152
rect 182730 229936 182786 229945
rect 182730 229871 182786 229880
rect 181838 226766 182036 226794
rect 182086 226808 182142 226817
rect 181166 226743 181222 226752
rect 182744 226780 182772 229871
rect 183756 226780 183784 230143
rect 184754 230072 184810 230081
rect 184754 230007 184810 230016
rect 184768 226780 184796 230007
rect 186240 226794 186268 261326
rect 187620 229094 187648 399638
rect 191748 399424 191800 399430
rect 191748 399366 191800 399372
rect 188988 399356 189040 399362
rect 188988 399298 189040 399304
rect 187700 396024 187752 396030
rect 187700 395966 187752 395972
rect 187712 248414 187740 395966
rect 187712 248386 188384 248414
rect 187974 233880 188030 233889
rect 187974 233815 188030 233824
rect 187160 229066 187648 229094
rect 187160 226794 187188 229066
rect 187988 226794 188016 233815
rect 185794 226766 186268 226794
rect 186714 226766 187188 226794
rect 187726 226766 188016 226794
rect 188356 226794 188384 248386
rect 189000 233889 189028 399298
rect 189080 396908 189132 396914
rect 189080 396850 189132 396856
rect 191104 396908 191156 396914
rect 191104 396850 191156 396856
rect 189092 248414 189120 396850
rect 191116 267102 191144 396850
rect 191380 390380 191432 390386
rect 191380 390322 191432 390328
rect 191392 387870 191420 390322
rect 191380 387864 191432 387870
rect 191380 387806 191432 387812
rect 191656 301504 191708 301510
rect 191656 301446 191708 301452
rect 191104 267096 191156 267102
rect 191104 267038 191156 267044
rect 189092 248386 189304 248414
rect 188986 233880 189042 233889
rect 188986 233815 189042 233824
rect 189276 226794 189304 248386
rect 190918 233880 190974 233889
rect 190918 233815 190974 233824
rect 190932 226794 190960 233815
rect 188356 226766 188738 226794
rect 189276 226766 189658 226794
rect 190670 226766 190960 226794
rect 191668 226780 191696 301446
rect 191760 233889 191788 399366
rect 193220 396840 193272 396846
rect 193220 396782 193272 396788
rect 191840 265532 191892 265538
rect 191840 265474 191892 265480
rect 191852 248414 191880 265474
rect 191852 248386 192248 248414
rect 191746 233880 191802 233889
rect 191746 233815 191802 233824
rect 192220 226794 192248 248386
rect 193232 226794 193260 396782
rect 194600 395888 194652 395894
rect 194600 395830 194652 395836
rect 193312 393304 193364 393310
rect 193312 393246 193364 393252
rect 193324 390386 193352 393246
rect 193312 390380 193364 390386
rect 193312 390322 193364 390328
rect 192220 226766 192694 226794
rect 193232 226766 193614 226794
rect 194612 226780 194640 395830
rect 195888 265464 195940 265470
rect 195888 265406 195940 265412
rect 195900 226794 195928 265406
rect 196544 236745 196572 700334
rect 196624 700324 196676 700330
rect 196624 700266 196676 700272
rect 196636 398206 196664 700266
rect 196900 566500 196952 566506
rect 196900 566442 196952 566448
rect 196714 487792 196770 487801
rect 196714 487727 196770 487736
rect 196624 398200 196676 398206
rect 196624 398142 196676 398148
rect 196624 396840 196676 396846
rect 196624 396782 196676 396788
rect 196636 263498 196664 396782
rect 196624 263492 196676 263498
rect 196624 263434 196676 263440
rect 196530 236736 196586 236745
rect 196530 236671 196586 236680
rect 196728 230217 196756 487727
rect 196806 483440 196862 483449
rect 196806 483375 196862 483384
rect 196714 230208 196770 230217
rect 196714 230143 196770 230152
rect 196820 229809 196848 483375
rect 196912 393378 196940 566442
rect 197910 486976 197966 486985
rect 197910 486911 197966 486920
rect 197358 479224 197414 479233
rect 197358 479159 197414 479168
rect 196900 393372 196952 393378
rect 196900 393314 196952 393320
rect 197268 265532 197320 265538
rect 197268 265474 197320 265480
rect 196806 229800 196862 229809
rect 196806 229735 196862 229744
rect 197280 229094 197308 265474
rect 197372 239465 197400 479159
rect 197544 264716 197596 264722
rect 197544 264658 197596 264664
rect 197452 264036 197504 264042
rect 197452 263978 197504 263984
rect 197358 239456 197414 239465
rect 197358 239391 197414 239400
rect 196912 229066 197308 229094
rect 196912 226794 196940 229066
rect 195638 226766 195928 226794
rect 196558 226766 196940 226794
rect 197464 226794 197492 263978
rect 197556 238754 197584 264658
rect 197924 239465 197952 486911
rect 198016 398138 198044 700742
rect 200764 700664 200816 700670
rect 200764 700606 200816 700612
rect 198646 486704 198702 486713
rect 198646 486639 198702 486648
rect 198278 486432 198334 486441
rect 198278 486367 198334 486376
rect 198094 485888 198150 485897
rect 198094 485823 198150 485832
rect 198004 398132 198056 398138
rect 198004 398074 198056 398080
rect 197910 239456 197966 239465
rect 197910 239391 197966 239400
rect 197556 238726 198044 238754
rect 198016 229094 198044 238726
rect 198108 229809 198136 485823
rect 198292 231169 198320 486367
rect 198462 486160 198518 486169
rect 198462 486095 198518 486104
rect 198370 485616 198426 485625
rect 198370 485551 198426 485560
rect 198278 231160 198334 231169
rect 198278 231095 198334 231104
rect 198384 230081 198412 485551
rect 198476 236881 198504 486095
rect 198554 483984 198610 483993
rect 198554 483919 198610 483928
rect 198462 236872 198518 236881
rect 198462 236807 198518 236816
rect 198370 230072 198426 230081
rect 198370 230007 198426 230016
rect 198568 229945 198596 483919
rect 198660 236745 198688 486639
rect 198830 419384 198886 419393
rect 198830 419319 198886 419328
rect 198738 417752 198794 417761
rect 198738 417687 198794 417696
rect 198646 236736 198702 236745
rect 198646 236671 198702 236680
rect 198752 236609 198780 417687
rect 198844 242185 198872 419319
rect 199014 416392 199070 416401
rect 199014 416327 199070 416336
rect 198922 413672 198978 413681
rect 198922 413607 198978 413616
rect 198936 262070 198964 413607
rect 199028 399838 199056 416327
rect 199382 414896 199438 414905
rect 199382 414831 199438 414840
rect 199016 399832 199068 399838
rect 199016 399774 199068 399780
rect 198924 262064 198976 262070
rect 198924 262006 198976 262012
rect 198830 242176 198886 242185
rect 198830 242111 198886 242120
rect 198738 236600 198794 236609
rect 198738 236535 198794 236544
rect 198554 229936 198610 229945
rect 198554 229871 198610 229880
rect 198094 229800 198150 229809
rect 198094 229735 198150 229744
rect 198016 229066 198136 229094
rect 198108 226794 198136 229066
rect 199396 228313 199424 414831
rect 200776 262478 200804 700606
rect 201408 262812 201460 262818
rect 201408 262754 201460 262760
rect 200764 262472 200816 262478
rect 200764 262414 200816 262420
rect 200028 260568 200080 260574
rect 200028 260510 200080 260516
rect 199382 228304 199438 228313
rect 199382 228239 199438 228248
rect 200040 226794 200068 260510
rect 201420 229094 201448 262754
rect 201512 260982 201540 702986
rect 218992 700874 219020 703520
rect 209136 700868 209188 700874
rect 209136 700810 209188 700816
rect 218980 700868 219032 700874
rect 218980 700810 219032 700816
rect 206284 700732 206336 700738
rect 206284 700674 206336 700680
rect 204904 700596 204956 700602
rect 204904 700538 204956 700544
rect 202878 487656 202934 487665
rect 202878 487591 202934 487600
rect 202142 486568 202198 486577
rect 202142 486503 202198 486512
rect 201684 263900 201736 263906
rect 201684 263842 201736 263848
rect 201500 260976 201552 260982
rect 201500 260918 201552 260924
rect 201696 248414 201724 263842
rect 201696 248386 202092 248414
rect 201774 233880 201830 233889
rect 201774 233815 201830 233824
rect 200960 229066 201448 229094
rect 200960 226794 200988 229066
rect 201788 226794 201816 233815
rect 202064 229094 202092 248386
rect 202156 231305 202184 486503
rect 202236 433356 202288 433362
rect 202236 433298 202288 433304
rect 202248 399362 202276 433298
rect 202236 399356 202288 399362
rect 202236 399298 202288 399304
rect 202788 262200 202840 262206
rect 202788 262142 202840 262148
rect 202800 233889 202828 262142
rect 202892 248414 202920 487591
rect 203522 486296 203578 486305
rect 203522 486231 203578 486240
rect 202892 248386 203104 248414
rect 202786 233880 202842 233889
rect 202786 233815 202842 233824
rect 202142 231296 202198 231305
rect 202142 231231 202198 231240
rect 202064 229066 202184 229094
rect 197464 226766 197570 226794
rect 198108 226766 198582 226794
rect 199594 226766 200068 226794
rect 200514 226766 200988 226794
rect 201526 226766 201816 226794
rect 202156 226794 202184 229066
rect 203076 226794 203104 248386
rect 203536 235249 203564 486231
rect 204260 266348 204312 266354
rect 204260 266290 204312 266296
rect 203522 235240 203578 235249
rect 203522 235175 203578 235184
rect 204272 226794 204300 266290
rect 204916 261118 204944 700538
rect 204996 429208 205048 429214
rect 204996 429150 205048 429156
rect 205008 267034 205036 429150
rect 204996 267028 205048 267034
rect 204996 266970 205048 266976
rect 205548 263492 205600 263498
rect 205548 263434 205600 263440
rect 204904 261112 204956 261118
rect 204904 261054 204956 261060
rect 205560 226794 205588 263434
rect 205640 262404 205692 262410
rect 205640 262346 205692 262352
rect 205652 248414 205680 262346
rect 206296 260098 206324 700674
rect 209044 700324 209096 700330
rect 209044 700266 209096 700272
rect 206376 670744 206428 670750
rect 206376 670686 206428 670692
rect 206388 260778 206416 670686
rect 206468 434784 206520 434790
rect 206468 434726 206520 434732
rect 206480 399430 206508 434726
rect 206468 399424 206520 399430
rect 206468 399366 206520 399372
rect 207020 266212 207072 266218
rect 207020 266154 207072 266160
rect 206376 260772 206428 260778
rect 206376 260714 206428 260720
rect 206284 260092 206336 260098
rect 206284 260034 206336 260040
rect 205652 248386 206048 248414
rect 205638 234832 205694 234841
rect 205638 234767 205694 234776
rect 205652 231985 205680 234767
rect 205638 231976 205694 231985
rect 205638 231911 205694 231920
rect 202156 226766 202538 226794
rect 203076 226766 203550 226794
rect 204272 226766 204470 226794
rect 205482 226766 205588 226794
rect 206020 226794 206048 248386
rect 207032 226794 207060 266154
rect 208400 264172 208452 264178
rect 208400 264114 208452 264120
rect 206020 226766 206494 226794
rect 207032 226766 207414 226794
rect 208412 226780 208440 264114
rect 209056 261254 209084 700266
rect 209148 400042 209176 700810
rect 235184 700806 235212 703520
rect 235172 700800 235224 700806
rect 235172 700742 235224 700748
rect 267660 700738 267688 703520
rect 267648 700732 267700 700738
rect 267648 700674 267700 700680
rect 283852 700670 283880 703520
rect 283840 700664 283892 700670
rect 283840 700606 283892 700612
rect 300136 700602 300164 703520
rect 300124 700596 300176 700602
rect 300124 700538 300176 700544
rect 332520 700534 332548 703520
rect 213184 700528 213236 700534
rect 213184 700470 213236 700476
rect 332508 700528 332560 700534
rect 332508 700470 332560 700476
rect 209778 485344 209834 485353
rect 209778 485279 209834 485288
rect 209136 400036 209188 400042
rect 209136 399978 209188 399984
rect 209688 264716 209740 264722
rect 209688 264658 209740 264664
rect 209044 261248 209096 261254
rect 209044 261190 209096 261196
rect 209700 226794 209728 264658
rect 209792 248414 209820 485279
rect 211804 409896 211856 409902
rect 211804 409838 211856 409844
rect 211816 398274 211844 409838
rect 213196 399974 213224 700470
rect 348804 700466 348832 703520
rect 215944 700460 215996 700466
rect 215944 700402 215996 700408
rect 348792 700460 348844 700466
rect 348792 700402 348844 700408
rect 214564 700392 214616 700398
rect 214564 700334 214616 700340
rect 213276 432404 213328 432410
rect 213276 432346 213328 432352
rect 213184 399968 213236 399974
rect 213184 399910 213236 399916
rect 211804 398268 211856 398274
rect 211804 398210 211856 398216
rect 213184 267028 213236 267034
rect 213184 266970 213236 266976
rect 211160 266280 211212 266286
rect 211160 266222 211212 266228
rect 211172 248414 211200 266222
rect 209792 248386 210096 248414
rect 211172 248386 211936 248414
rect 209438 226766 209728 226794
rect 210068 226794 210096 248386
rect 211342 230480 211398 230489
rect 211342 230415 211398 230424
rect 210068 226766 210450 226794
rect 211356 226780 211384 230415
rect 211908 226794 211936 248386
rect 213196 230489 213224 266970
rect 213288 265878 213316 432346
rect 213920 269816 213972 269822
rect 213920 269758 213972 269764
rect 213276 265872 213328 265878
rect 213276 265814 213328 265820
rect 213828 263560 213880 263566
rect 213828 263502 213880 263508
rect 213182 230480 213238 230489
rect 213182 230415 213238 230424
rect 213840 226794 213868 263502
rect 211908 226766 212382 226794
rect 213394 226766 213868 226794
rect 213932 226794 213960 269758
rect 214576 260846 214604 700334
rect 215956 399906 215984 700402
rect 364996 700398 365024 703520
rect 385684 700596 385736 700602
rect 385684 700538 385736 700544
rect 370504 700460 370556 700466
rect 370504 700402 370556 700408
rect 364984 700392 365036 700398
rect 364984 700334 365036 700340
rect 367744 616888 367796 616894
rect 367744 616830 367796 616836
rect 363604 563100 363656 563106
rect 363604 563042 363656 563048
rect 360844 510672 360896 510678
rect 360844 510614 360896 510620
rect 266082 490104 266138 490113
rect 266082 490039 266138 490048
rect 217782 489016 217838 489025
rect 217782 488951 217838 488960
rect 263598 489016 263654 489025
rect 263598 488951 263654 488960
rect 217690 487656 217746 487665
rect 217690 487591 217746 487600
rect 217322 487248 217378 487257
rect 217322 487183 217378 487192
rect 216586 485344 216642 485353
rect 216586 485279 216642 485288
rect 215944 399900 215996 399906
rect 215944 399842 215996 399848
rect 215300 264104 215352 264110
rect 215300 264046 215352 264052
rect 214564 260840 214616 260846
rect 214564 260782 214616 260788
rect 215312 248414 215340 264046
rect 215312 248386 215984 248414
rect 215574 233880 215630 233889
rect 215574 233815 215630 233824
rect 215588 226794 215616 233815
rect 213932 226766 214406 226794
rect 215326 226766 215616 226794
rect 215956 226794 215984 248386
rect 216600 233889 216628 485279
rect 217336 484537 217364 487183
rect 217414 486840 217470 486849
rect 217414 486775 217470 486784
rect 217322 484528 217378 484537
rect 217322 484463 217378 484472
rect 216678 435976 216734 435985
rect 216678 435911 216734 435920
rect 216692 434790 216720 435911
rect 216680 434784 216732 434790
rect 216680 434726 216732 434732
rect 216678 433800 216734 433809
rect 216678 433735 216734 433744
rect 216692 433362 216720 433735
rect 216680 433356 216732 433362
rect 216680 433298 216732 433304
rect 216678 432848 216734 432857
rect 216678 432783 216734 432792
rect 216692 432410 216720 432783
rect 216680 432404 216732 432410
rect 216680 432346 216732 432352
rect 216678 429992 216734 430001
rect 216678 429927 216734 429936
rect 216692 429214 216720 429927
rect 216680 429208 216732 429214
rect 216680 429150 216732 429156
rect 217230 428224 217286 428233
rect 217230 428159 217286 428168
rect 216678 410000 216734 410009
rect 216678 409935 216734 409944
rect 216692 409902 216720 409935
rect 216680 409896 216732 409902
rect 216680 409838 216732 409844
rect 217138 408096 217194 408105
rect 217138 408031 217194 408040
rect 217152 233889 217180 408031
rect 217244 399770 217272 428159
rect 217336 408377 217364 484463
rect 217322 408368 217378 408377
rect 217322 408303 217378 408312
rect 217336 400110 217364 408303
rect 217324 400104 217376 400110
rect 217324 400046 217376 400052
rect 217232 399764 217284 399770
rect 217232 399706 217284 399712
rect 216586 233880 216642 233889
rect 216586 233815 216642 233824
rect 217138 233880 217194 233889
rect 217138 233815 217194 233824
rect 217428 227089 217456 486775
rect 217598 485888 217654 485897
rect 217598 485823 217654 485832
rect 217506 431080 217562 431089
rect 217506 431015 217562 431024
rect 217520 399770 217548 431015
rect 217508 399764 217560 399770
rect 217508 399706 217560 399712
rect 217612 398206 217640 485823
rect 217704 398274 217732 487591
rect 217692 398268 217744 398274
rect 217692 398210 217744 398216
rect 217600 398200 217652 398206
rect 217600 398142 217652 398148
rect 217796 398138 217824 488951
rect 256146 487656 256202 487665
rect 256146 487591 256202 487600
rect 217874 487520 217930 487529
rect 217874 487455 217930 487464
rect 217888 398177 217916 487455
rect 218242 486976 218298 486985
rect 218242 486911 218298 486920
rect 218058 484528 218114 484537
rect 218058 484463 218114 484472
rect 217966 436928 218022 436937
rect 217966 436863 218022 436872
rect 217874 398168 217930 398177
rect 217784 398132 217836 398138
rect 217874 398103 217930 398112
rect 217784 398074 217836 398080
rect 217690 235920 217746 235929
rect 217690 235855 217746 235864
rect 217414 227080 217470 227089
rect 217414 227015 217470 227024
rect 217704 226794 217732 235855
rect 217980 229945 218008 436863
rect 218072 398041 218100 484463
rect 218150 483576 218206 483585
rect 218150 483511 218206 483520
rect 218058 398032 218114 398041
rect 218058 397967 218114 397976
rect 218164 231713 218192 483511
rect 218256 399537 218284 486911
rect 218978 486840 219034 486849
rect 218978 486775 219034 486784
rect 218610 486704 218666 486713
rect 218610 486639 218666 486648
rect 218426 486432 218482 486441
rect 218426 486367 218482 486376
rect 218334 483712 218390 483721
rect 218334 483647 218390 483656
rect 218242 399528 218298 399537
rect 218242 399463 218298 399472
rect 218150 231704 218206 231713
rect 218150 231639 218206 231648
rect 218348 231441 218376 483647
rect 218440 399838 218468 486367
rect 218518 485208 218574 485217
rect 218518 485143 218574 485152
rect 218428 399832 218480 399838
rect 218428 399774 218480 399780
rect 218426 267744 218482 267753
rect 218426 267679 218482 267688
rect 218440 258369 218468 267679
rect 218426 258360 218482 258369
rect 218426 258295 218482 258304
rect 218426 257952 218482 257961
rect 218426 257887 218482 257896
rect 218440 248441 218468 257887
rect 218426 248432 218482 248441
rect 218426 248367 218482 248376
rect 218426 248024 218482 248033
rect 218426 247959 218482 247968
rect 218440 238921 218468 247959
rect 218426 238912 218482 238921
rect 218426 238847 218482 238856
rect 218532 238754 218560 485143
rect 218624 399906 218652 486639
rect 218702 486024 218758 486033
rect 218702 485959 218758 485968
rect 218612 399900 218664 399906
rect 218612 399842 218664 399848
rect 218610 398304 218666 398313
rect 218610 398239 218666 398248
rect 218624 393417 218652 398239
rect 218610 393408 218666 393417
rect 218610 393343 218666 393352
rect 218612 260500 218664 260506
rect 218612 260442 218664 260448
rect 218440 238726 218560 238754
rect 218334 231432 218390 231441
rect 218334 231367 218390 231376
rect 218440 231033 218468 238726
rect 218518 238504 218574 238513
rect 218518 238439 218574 238448
rect 218532 235113 218560 238439
rect 218518 235104 218574 235113
rect 218518 235039 218574 235048
rect 218426 231024 218482 231033
rect 218426 230959 218482 230968
rect 217966 229936 218022 229945
rect 217966 229871 218022 229880
rect 218624 226794 218652 260442
rect 215956 226766 216338 226794
rect 217350 226766 217732 226794
rect 218270 226766 218652 226794
rect 182086 226743 182142 226752
rect 77390 226672 77446 226681
rect 77234 226630 77390 226658
rect 77390 226607 77446 226616
rect 62118 226536 62174 226545
rect 75550 226536 75606 226545
rect 62174 226494 62422 226522
rect 75210 226494 75550 226522
rect 62118 226471 62174 226480
rect 75550 226471 75606 226480
rect 68558 226400 68614 226409
rect 68310 226358 68558 226386
rect 68558 226335 68614 226344
rect 218716 226273 218744 485959
rect 218794 485072 218850 485081
rect 218794 485007 218850 485016
rect 218808 228721 218836 485007
rect 218886 483304 218942 483313
rect 218886 483239 218942 483248
rect 218900 231849 218928 483239
rect 218992 399974 219020 486775
rect 219990 486568 220046 486577
rect 219990 486503 220046 486512
rect 219806 486296 219862 486305
rect 219806 486231 219862 486240
rect 219346 486160 219402 486169
rect 219346 486095 219402 486104
rect 219254 485752 219310 485761
rect 219254 485687 219310 485696
rect 219162 483848 219218 483857
rect 219162 483783 219218 483792
rect 219070 483304 219126 483313
rect 219070 483239 219126 483248
rect 218980 399968 219032 399974
rect 218980 399910 219032 399916
rect 219084 393314 219112 483239
rect 218992 393286 219112 393314
rect 218992 374082 219020 393286
rect 219072 392964 219124 392970
rect 219072 392906 219124 392912
rect 219084 383790 219112 392906
rect 219072 383784 219124 383790
rect 219072 383726 219124 383732
rect 219070 383616 219126 383625
rect 219070 383551 219126 383560
rect 219084 374241 219112 383551
rect 219070 374232 219126 374241
rect 219070 374167 219126 374176
rect 218992 374054 219112 374082
rect 218978 373960 219034 373969
rect 218978 373895 219034 373904
rect 218992 364449 219020 373895
rect 218978 364440 219034 364449
rect 218978 364375 219034 364384
rect 218978 364304 219034 364313
rect 218978 364239 219034 364248
rect 218992 354793 219020 364239
rect 218978 354784 219034 354793
rect 218978 354719 219034 354728
rect 218978 354648 219034 354657
rect 218978 354583 219034 354592
rect 218992 345137 219020 354583
rect 218978 345128 219034 345137
rect 218978 345063 219034 345072
rect 219084 345014 219112 374054
rect 218992 344986 219112 345014
rect 218992 316146 219020 344986
rect 219070 344584 219126 344593
rect 219070 344519 219126 344528
rect 219084 335481 219112 344519
rect 219070 335472 219126 335481
rect 219070 335407 219126 335416
rect 219072 335164 219124 335170
rect 219072 335106 219124 335112
rect 219084 325854 219112 335106
rect 219072 325848 219124 325854
rect 219072 325790 219124 325796
rect 219070 325680 219126 325689
rect 219070 325615 219126 325624
rect 219084 316305 219112 325615
rect 219070 316296 219126 316305
rect 219070 316231 219126 316240
rect 218992 316118 219112 316146
rect 218978 316024 219034 316033
rect 218978 315959 219034 315968
rect 218992 306513 219020 315959
rect 218978 306504 219034 306513
rect 218978 306439 219034 306448
rect 218978 306368 219034 306377
rect 218978 306303 219034 306312
rect 218992 296857 219020 306303
rect 218978 296848 219034 296857
rect 218978 296783 219034 296792
rect 218978 296712 219034 296721
rect 218978 296647 219034 296656
rect 218992 287201 219020 296647
rect 218978 287192 219034 287201
rect 218978 287127 219034 287136
rect 218978 287056 219034 287065
rect 218978 286991 219034 287000
rect 218992 277545 219020 286991
rect 218978 277536 219034 277545
rect 218978 277471 219034 277480
rect 218978 277400 219034 277409
rect 218978 277335 219034 277344
rect 218992 267889 219020 277335
rect 218978 267880 219034 267889
rect 218978 267815 219034 267824
rect 218980 262132 219032 262138
rect 218980 262074 219032 262080
rect 218886 231840 218942 231849
rect 218886 231775 218942 231784
rect 218794 228712 218850 228721
rect 218794 228647 218850 228656
rect 218992 226794 219020 262074
rect 219084 230081 219112 316118
rect 219070 230072 219126 230081
rect 219070 230007 219126 230016
rect 219176 228585 219204 483783
rect 219268 231577 219296 485687
rect 219360 392970 219388 486095
rect 219622 486024 219678 486033
rect 219622 485959 219678 485968
rect 219636 484265 219664 485959
rect 219714 485208 219770 485217
rect 219714 485143 219770 485152
rect 219622 484256 219678 484265
rect 219622 484191 219678 484200
rect 219438 484120 219494 484129
rect 219438 484055 219494 484064
rect 219452 398478 219480 484055
rect 219530 483848 219586 483857
rect 219530 483783 219586 483792
rect 219544 398682 219572 483783
rect 219622 483712 219678 483721
rect 219622 483647 219678 483656
rect 219532 398676 219584 398682
rect 219532 398618 219584 398624
rect 219636 398614 219664 483647
rect 219728 403209 219756 485143
rect 219714 403200 219770 403209
rect 219714 403135 219770 403144
rect 219716 403096 219768 403102
rect 219716 403038 219768 403044
rect 219624 398608 219676 398614
rect 219624 398550 219676 398556
rect 219440 398472 219492 398478
rect 219440 398414 219492 398420
rect 219728 398206 219756 403038
rect 219716 398200 219768 398206
rect 219716 398142 219768 398148
rect 219348 392964 219400 392970
rect 219348 392906 219400 392912
rect 219346 392864 219402 392873
rect 219346 392799 219402 392808
rect 219360 383897 219388 392799
rect 219346 383888 219402 383897
rect 219346 383823 219402 383832
rect 219348 383716 219400 383722
rect 219348 383658 219400 383664
rect 219360 335170 219388 383658
rect 219348 335164 219400 335170
rect 219348 335106 219400 335112
rect 219346 335064 219402 335073
rect 219346 334999 219402 335008
rect 219360 325961 219388 334999
rect 219346 325952 219402 325961
rect 219346 325887 219402 325896
rect 219348 325848 219400 325854
rect 219348 325790 219400 325796
rect 219254 231568 219310 231577
rect 219254 231503 219310 231512
rect 219162 228576 219218 228585
rect 219162 228511 219218 228520
rect 219360 227225 219388 325790
rect 219440 265600 219492 265606
rect 219440 265542 219492 265548
rect 219452 229094 219480 265542
rect 219820 234025 219848 486231
rect 219898 483576 219954 483585
rect 219898 483511 219954 483520
rect 219912 403102 219940 483511
rect 219900 403096 219952 403102
rect 219900 403038 219952 403044
rect 219898 402928 219954 402937
rect 219898 402863 219954 402872
rect 219806 234016 219862 234025
rect 219806 233951 219862 233960
rect 219452 229066 219848 229094
rect 219346 227216 219402 227225
rect 219346 227151 219402 227160
rect 219820 226794 219848 229066
rect 219912 228449 219940 402863
rect 220004 229094 220032 486503
rect 256160 485897 256188 487591
rect 263612 485897 263640 488951
rect 266096 486849 266124 490039
rect 316038 489968 316094 489977
rect 316038 489903 316094 489912
rect 276202 488880 276258 488889
rect 276202 488815 276258 488824
rect 266082 486840 266138 486849
rect 266082 486775 266138 486784
rect 276216 485897 276244 488815
rect 301042 488744 301098 488753
rect 301042 488679 301098 488688
rect 256146 485888 256202 485897
rect 256146 485823 256202 485832
rect 263598 485888 263654 485897
rect 263598 485823 263654 485832
rect 276202 485888 276258 485897
rect 276202 485823 276258 485832
rect 301056 485081 301084 488679
rect 303434 488608 303490 488617
rect 303434 488543 303490 488552
rect 303448 485897 303476 488543
rect 316052 486577 316080 489903
rect 318706 487384 318762 487393
rect 318706 487319 318762 487328
rect 316038 486568 316094 486577
rect 316038 486503 316094 486512
rect 318720 486441 318748 487319
rect 340142 487248 340198 487257
rect 340142 487183 340198 487192
rect 340156 486441 340184 487183
rect 315946 486432 316002 486441
rect 315946 486367 316002 486376
rect 318706 486432 318762 486441
rect 318706 486367 318762 486376
rect 340142 486432 340198 486441
rect 340142 486367 340198 486376
rect 303434 485888 303490 485897
rect 303434 485823 303490 485832
rect 301042 485072 301098 485081
rect 301042 485007 301098 485016
rect 315960 483857 315988 486367
rect 356518 485888 356574 485897
rect 356518 485823 356574 485832
rect 315946 483848 316002 483857
rect 315946 483783 316002 483792
rect 227352 399968 227404 399974
rect 220082 399936 220138 399945
rect 227352 399910 227404 399916
rect 220082 399871 220138 399880
rect 226432 399900 226484 399906
rect 220096 398138 220124 399871
rect 226432 399842 226484 399848
rect 224960 398676 225012 398682
rect 224960 398618 225012 398624
rect 224776 398608 224828 398614
rect 224776 398550 224828 398556
rect 220084 398132 220136 398138
rect 220084 398074 220136 398080
rect 220084 396364 220136 396370
rect 220084 396306 220136 396312
rect 220096 235929 220124 396306
rect 222200 395616 222252 395622
rect 222200 395558 222252 395564
rect 224684 395616 224736 395622
rect 224684 395558 224736 395564
rect 222108 262064 222160 262070
rect 222108 262006 222160 262012
rect 220082 235920 220138 235929
rect 220082 235855 220138 235864
rect 222120 229094 222148 262006
rect 220004 229066 220584 229094
rect 219898 228440 219954 228449
rect 219898 228375 219954 228384
rect 218992 226766 219282 226794
rect 219820 226766 220294 226794
rect 220556 226273 220584 229066
rect 221752 229066 222148 229094
rect 221752 226794 221780 229066
rect 221306 226766 221780 226794
rect 222212 226780 222240 395558
rect 223580 358080 223632 358086
rect 223580 358022 223632 358028
rect 223210 230072 223266 230081
rect 223210 230007 223266 230016
rect 223224 226780 223252 230007
rect 223592 226273 223620 358022
rect 224696 238754 224724 395558
rect 224512 238726 224724 238754
rect 224512 226794 224540 238726
rect 224590 229256 224646 229265
rect 224590 229191 224646 229200
rect 224250 226766 224540 226794
rect 224604 226273 224632 229191
rect 61162 226222 61240 226250
rect 61934 226264 61990 226273
rect 61106 226199 61162 226208
rect 61934 226199 61990 226208
rect 218702 226264 218758 226273
rect 218702 226199 218758 226208
rect 220542 226264 220598 226273
rect 220542 226199 220598 226208
rect 223578 226264 223634 226273
rect 223578 226199 223634 226208
rect 224590 226264 224646 226273
rect 224590 226199 224646 226208
rect 59832 180766 59952 180794
rect 59832 175642 59860 180766
rect 59820 175636 59872 175642
rect 59820 175578 59872 175584
rect 59542 138816 59598 138825
rect 59542 138751 59598 138760
rect 59372 74506 59768 74534
rect 59266 67280 59322 67289
rect 59266 67215 59322 67224
rect 59740 60058 59768 74506
rect 224406 60344 224462 60353
rect 224462 60302 224526 60330
rect 224406 60279 224462 60288
rect 222658 60208 222714 60217
rect 222502 60166 222658 60194
rect 222658 60143 222714 60152
rect 211894 60072 211950 60081
rect 59740 60030 60122 60058
rect 60200 60030 60398 60058
rect 60476 60030 60674 60058
rect 59740 59922 59768 60030
rect 59372 59894 59768 59922
rect 59268 57996 59320 58002
rect 59268 57938 59320 57944
rect 58898 57896 58954 57905
rect 58898 57831 58954 57840
rect 59280 57322 59308 57938
rect 59268 57316 59320 57322
rect 59268 57258 59320 57264
rect 58622 57080 58678 57089
rect 58622 57015 58678 57024
rect 59268 56704 59320 56710
rect 59268 56646 59320 56652
rect 57244 56636 57296 56642
rect 57244 56578 57296 56584
rect 55772 55888 55824 55894
rect 55772 55830 55824 55836
rect 55680 20664 55732 20670
rect 55680 20606 55732 20612
rect 57256 6914 57284 56578
rect 54956 6886 55168 6914
rect 57164 6886 57284 6914
rect 53840 3052 53892 3058
rect 53840 2994 53892 3000
rect 53852 2854 53880 2994
rect 53840 2848 53892 2854
rect 53840 2790 53892 2796
rect 54956 480 54984 6886
rect 55680 3800 55732 3806
rect 55680 3742 55732 3748
rect 55772 3800 55824 3806
rect 55772 3742 55824 3748
rect 55692 3641 55720 3742
rect 55784 3670 55812 3742
rect 55772 3664 55824 3670
rect 55678 3632 55734 3641
rect 55772 3606 55824 3612
rect 55678 3567 55734 3576
rect 57164 3534 57192 6886
rect 59280 3534 59308 56646
rect 56048 3528 56100 3534
rect 56048 3470 56100 3476
rect 57152 3528 57204 3534
rect 57152 3470 57204 3476
rect 58440 3528 58492 3534
rect 58440 3470 58492 3476
rect 59268 3528 59320 3534
rect 59268 3470 59320 3476
rect 56060 480 56088 3470
rect 57244 2848 57296 2854
rect 57244 2790 57296 2796
rect 57256 480 57284 2790
rect 58452 480 58480 3470
rect 59372 3369 59400 59894
rect 60200 57610 60228 60030
rect 59556 57582 60228 57610
rect 59452 57316 59504 57322
rect 59452 57258 59504 57264
rect 59464 3602 59492 57258
rect 59452 3596 59504 3602
rect 59452 3538 59504 3544
rect 59556 3466 59584 57582
rect 60002 57488 60058 57497
rect 60002 57423 60058 57432
rect 60016 3738 60044 57423
rect 60476 57322 60504 60030
rect 60464 57316 60516 57322
rect 60464 57258 60516 57264
rect 60936 57225 60964 60044
rect 61028 60030 61226 60058
rect 61304 60030 61502 60058
rect 61580 60030 61870 60058
rect 60922 57216 60978 57225
rect 60922 57151 60978 57160
rect 60648 54664 60700 54670
rect 60648 54606 60700 54612
rect 60004 3732 60056 3738
rect 60004 3674 60056 3680
rect 59726 3632 59782 3641
rect 59726 3567 59728 3576
rect 59780 3567 59782 3576
rect 59728 3538 59780 3544
rect 60660 3534 60688 54606
rect 61028 51074 61056 60030
rect 61304 58002 61332 60030
rect 61292 57996 61344 58002
rect 61292 57938 61344 57944
rect 60844 51046 61056 51074
rect 60844 6914 60872 51046
rect 61580 45554 61608 60030
rect 62132 57769 62160 60044
rect 62118 57760 62174 57769
rect 61936 57724 61988 57730
rect 62118 57695 62174 57704
rect 61936 57666 61988 57672
rect 61842 57216 61898 57225
rect 61948 57186 61976 57666
rect 62028 57656 62080 57662
rect 62212 57656 62264 57662
rect 62080 57604 62212 57610
rect 62028 57598 62264 57604
rect 62040 57582 62252 57598
rect 62408 57361 62436 60044
rect 62684 57633 62712 60044
rect 62670 57624 62726 57633
rect 62670 57559 62726 57568
rect 62960 57497 62988 60044
rect 62946 57488 63002 57497
rect 62946 57423 63002 57432
rect 62394 57352 62450 57361
rect 62028 57316 62080 57322
rect 62394 57287 62450 57296
rect 62028 57258 62080 57264
rect 61842 57151 61844 57160
rect 61896 57151 61898 57160
rect 61936 57180 61988 57186
rect 61844 57122 61896 57128
rect 61936 57122 61988 57128
rect 60752 6886 60872 6914
rect 61028 45526 61608 45554
rect 60752 3670 60780 6886
rect 61028 3806 61056 45526
rect 61016 3800 61068 3806
rect 61016 3742 61068 3748
rect 60832 3732 60884 3738
rect 60832 3674 60884 3680
rect 60740 3664 60792 3670
rect 60740 3606 60792 3612
rect 59636 3528 59688 3534
rect 59636 3470 59688 3476
rect 60648 3528 60700 3534
rect 60648 3470 60700 3476
rect 59544 3460 59596 3466
rect 59544 3402 59596 3408
rect 59358 3360 59414 3369
rect 59358 3295 59414 3304
rect 59648 480 59676 3470
rect 60844 480 60872 3674
rect 62040 480 62068 57258
rect 63236 56817 63264 60044
rect 63604 56953 63632 60044
rect 63776 57044 63828 57050
rect 63776 56986 63828 56992
rect 63788 56953 63816 56986
rect 63590 56944 63646 56953
rect 63590 56879 63646 56888
rect 63774 56944 63830 56953
rect 63774 56879 63830 56888
rect 63408 56840 63460 56846
rect 63222 56808 63278 56817
rect 63222 56743 63278 56752
rect 63406 56808 63408 56817
rect 63460 56808 63462 56817
rect 63406 56743 63462 56752
rect 63500 55616 63552 55622
rect 63500 55558 63552 55564
rect 63512 3942 63540 55558
rect 63684 55548 63736 55554
rect 63684 55490 63736 55496
rect 63696 4010 63724 55490
rect 63684 4004 63736 4010
rect 63684 3946 63736 3952
rect 63500 3936 63552 3942
rect 63500 3878 63552 3884
rect 63880 3602 63908 60044
rect 64156 56681 64184 60044
rect 64248 60030 64446 60058
rect 64524 60030 64722 60058
rect 64142 56672 64198 56681
rect 64142 56607 64198 56616
rect 64248 55622 64276 60030
rect 64236 55616 64288 55622
rect 64236 55558 64288 55564
rect 64524 55554 64552 60030
rect 64696 57996 64748 58002
rect 64696 57938 64748 57944
rect 64708 56642 64736 57938
rect 64880 57860 64932 57866
rect 64880 57802 64932 57808
rect 64892 57526 64920 57802
rect 64880 57520 64932 57526
rect 64880 57462 64932 57468
rect 64880 57180 64932 57186
rect 64880 57122 64932 57128
rect 64788 56772 64840 56778
rect 64788 56714 64840 56720
rect 64696 56636 64748 56642
rect 64696 56578 64748 56584
rect 64800 56506 64828 56714
rect 64892 56574 64920 57122
rect 64880 56568 64932 56574
rect 64880 56510 64932 56516
rect 64788 56500 64840 56506
rect 64788 56442 64840 56448
rect 64512 55548 64564 55554
rect 64512 55490 64564 55496
rect 64984 3874 65012 60044
rect 65076 60030 65366 60058
rect 65444 60030 65642 60058
rect 65076 4078 65104 60030
rect 65248 57180 65300 57186
rect 65248 57122 65300 57128
rect 65156 56908 65208 56914
rect 65156 56850 65208 56856
rect 65168 56522 65196 56850
rect 65260 56642 65288 57122
rect 65340 56772 65392 56778
rect 65340 56714 65392 56720
rect 65248 56636 65300 56642
rect 65248 56578 65300 56584
rect 65352 56522 65380 56714
rect 65168 56494 65380 56522
rect 65444 45554 65472 60030
rect 65904 57254 65932 60044
rect 65996 60030 66194 60058
rect 65996 57458 66024 60030
rect 66168 57520 66220 57526
rect 66168 57462 66220 57468
rect 65984 57452 66036 57458
rect 65984 57394 66036 57400
rect 65892 57248 65944 57254
rect 65892 57190 65944 57196
rect 65522 56944 65578 56953
rect 65522 56879 65524 56888
rect 65576 56879 65578 56888
rect 65524 56850 65576 56856
rect 65616 56840 65668 56846
rect 65614 56808 65616 56817
rect 65668 56808 65670 56817
rect 65614 56743 65670 56752
rect 65168 45526 65472 45554
rect 65168 4146 65196 45526
rect 65156 4140 65208 4146
rect 65156 4082 65208 4088
rect 65064 4072 65116 4078
rect 65064 4014 65116 4020
rect 64972 3868 65024 3874
rect 64972 3810 65024 3816
rect 63868 3596 63920 3602
rect 63868 3538 63920 3544
rect 64328 3596 64380 3602
rect 64328 3538 64380 3544
rect 63224 3528 63276 3534
rect 63224 3470 63276 3476
rect 63236 480 63264 3470
rect 64340 480 64368 3538
rect 66180 3466 66208 57462
rect 66456 57390 66484 60044
rect 66732 57594 66760 60044
rect 66824 60030 67114 60058
rect 67192 60030 67390 60058
rect 67666 60030 67864 60058
rect 66720 57588 66772 57594
rect 66720 57530 66772 57536
rect 66444 57384 66496 57390
rect 66444 57326 66496 57332
rect 66824 51074 66852 60030
rect 66904 57588 66956 57594
rect 66904 57530 66956 57536
rect 66916 57225 66944 57530
rect 66902 57216 66958 57225
rect 66902 57151 66958 57160
rect 66364 51046 66852 51074
rect 65524 3460 65576 3466
rect 65524 3402 65576 3408
rect 66168 3460 66220 3466
rect 66168 3402 66220 3408
rect 65536 480 65564 3402
rect 66364 3398 66392 51046
rect 67192 45554 67220 60030
rect 67548 57384 67600 57390
rect 67548 57326 67600 57332
rect 66548 45526 67220 45554
rect 66352 3392 66404 3398
rect 66352 3334 66404 3340
rect 66548 3330 66576 45526
rect 67560 3466 67588 57326
rect 66720 3460 66772 3466
rect 66720 3402 66772 3408
rect 67548 3460 67600 3466
rect 67548 3402 67600 3408
rect 66536 3324 66588 3330
rect 66536 3266 66588 3272
rect 66732 480 66760 3402
rect 67836 3262 67864 60030
rect 67928 57730 67956 60044
rect 67916 57724 67968 57730
rect 67916 57666 67968 57672
rect 68204 57662 68232 60044
rect 68480 57798 68508 60044
rect 68572 60030 68862 60058
rect 69138 60030 69244 60058
rect 68468 57792 68520 57798
rect 68468 57734 68520 57740
rect 68192 57656 68244 57662
rect 68192 57598 68244 57604
rect 68572 55570 68600 60030
rect 68928 57248 68980 57254
rect 68928 57190 68980 57196
rect 68652 57180 68704 57186
rect 68652 57122 68704 57128
rect 68020 55542 68600 55570
rect 67916 3460 67968 3466
rect 67916 3402 67968 3408
rect 67824 3256 67876 3262
rect 67824 3198 67876 3204
rect 67928 480 67956 3402
rect 68020 3126 68048 55542
rect 68664 51074 68692 57122
rect 68296 51046 68692 51074
rect 68008 3120 68060 3126
rect 68008 3062 68060 3068
rect 68296 2854 68324 51046
rect 68940 3466 68968 57190
rect 69112 3596 69164 3602
rect 69112 3538 69164 3544
rect 68928 3460 68980 3466
rect 68928 3402 68980 3408
rect 68284 2848 68336 2854
rect 68284 2790 68336 2796
rect 69124 480 69152 3538
rect 69216 3194 69244 60030
rect 69400 54534 69428 60044
rect 69676 56710 69704 60044
rect 69952 57458 69980 60044
rect 70228 57594 70256 60044
rect 70216 57588 70268 57594
rect 70216 57530 70268 57536
rect 69940 57452 69992 57458
rect 69940 57394 69992 57400
rect 70216 57452 70268 57458
rect 70216 57394 70268 57400
rect 69664 56704 69716 56710
rect 69664 56646 69716 56652
rect 69388 54528 69440 54534
rect 69388 54470 69440 54476
rect 70228 16574 70256 57394
rect 70308 56704 70360 56710
rect 70308 56646 70360 56652
rect 70136 16546 70256 16574
rect 70136 3482 70164 16546
rect 70320 6914 70348 56646
rect 70228 6886 70348 6914
rect 70228 3602 70256 6886
rect 70216 3596 70268 3602
rect 70216 3538 70268 3544
rect 70136 3454 70348 3482
rect 69204 3188 69256 3194
rect 69204 3130 69256 3136
rect 70320 480 70348 3454
rect 70596 3058 70624 60044
rect 70872 57798 70900 60044
rect 70964 60030 71162 60058
rect 70860 57792 70912 57798
rect 70860 57734 70912 57740
rect 70964 45554 70992 60030
rect 71424 57050 71452 60044
rect 71516 60030 71714 60058
rect 71792 60030 71990 60058
rect 72068 60030 72358 60058
rect 72436 60030 72634 60058
rect 71412 57044 71464 57050
rect 71412 56986 71464 56992
rect 71516 56982 71544 60030
rect 71688 57588 71740 57594
rect 71688 57530 71740 57536
rect 71504 56976 71556 56982
rect 71504 56918 71556 56924
rect 70688 45526 70992 45554
rect 70584 3052 70636 3058
rect 70584 2994 70636 3000
rect 70688 2990 70716 45526
rect 71700 6914 71728 57530
rect 71792 56914 71820 60030
rect 72068 57644 72096 60030
rect 71884 57616 72096 57644
rect 71780 56908 71832 56914
rect 71780 56850 71832 56856
rect 71884 54602 71912 57616
rect 71872 54596 71924 54602
rect 71872 54538 71924 54544
rect 72436 45554 72464 60030
rect 72896 56846 72924 60044
rect 73068 57724 73120 57730
rect 73068 57666 73120 57672
rect 72884 56840 72936 56846
rect 72884 56782 72936 56788
rect 71516 6886 71728 6914
rect 72068 45526 72464 45554
rect 70676 2984 70728 2990
rect 70676 2926 70728 2932
rect 71516 480 71544 6886
rect 72068 2922 72096 45526
rect 73080 3466 73108 57666
rect 73172 56778 73200 60044
rect 73160 56772 73212 56778
rect 73160 56714 73212 56720
rect 73448 56642 73476 60044
rect 73724 57662 73752 60044
rect 73712 57656 73764 57662
rect 73712 57598 73764 57604
rect 74092 57186 74120 60044
rect 74080 57180 74132 57186
rect 74080 57122 74132 57128
rect 74368 57118 74396 60044
rect 74658 60030 74856 60058
rect 74724 57656 74776 57662
rect 74724 57598 74776 57604
rect 74356 57112 74408 57118
rect 74356 57054 74408 57060
rect 73436 56636 73488 56642
rect 73436 56578 73488 56584
rect 73804 3596 73856 3602
rect 73804 3538 73856 3544
rect 72608 3460 72660 3466
rect 72608 3402 72660 3408
rect 73068 3460 73120 3466
rect 73068 3402 73120 3408
rect 72056 2916 72108 2922
rect 72056 2858 72108 2864
rect 72620 480 72648 3402
rect 73816 480 73844 3538
rect 74736 3534 74764 57598
rect 74828 56982 74856 60030
rect 74816 56976 74868 56982
rect 74816 56918 74868 56924
rect 74816 56228 74868 56234
rect 74816 56170 74868 56176
rect 74828 3670 74856 56170
rect 74920 3738 74948 60044
rect 75196 57322 75224 60044
rect 75288 60030 75578 60058
rect 75656 60030 75854 60058
rect 75288 57662 75316 60030
rect 75276 57656 75328 57662
rect 75276 57598 75328 57604
rect 75184 57316 75236 57322
rect 75184 57258 75236 57264
rect 75000 56976 75052 56982
rect 75000 56918 75052 56924
rect 75012 54670 75040 56918
rect 75656 56234 75684 60030
rect 76116 57526 76144 60044
rect 76104 57520 76156 57526
rect 76104 57462 76156 57468
rect 76392 57390 76420 60044
rect 76484 60030 76682 60058
rect 76380 57384 76432 57390
rect 76380 57326 76432 57332
rect 76484 57254 76512 60030
rect 76656 57656 76708 57662
rect 76656 57598 76708 57604
rect 76472 57248 76524 57254
rect 76472 57190 76524 57196
rect 76564 56908 76616 56914
rect 76564 56850 76616 56856
rect 75644 56228 75696 56234
rect 75644 56170 75696 56176
rect 75000 54664 75052 54670
rect 75000 54606 75052 54612
rect 74908 3732 74960 3738
rect 74908 3674 74960 3680
rect 74816 3664 74868 3670
rect 74816 3606 74868 3612
rect 76576 3602 76604 56850
rect 76564 3596 76616 3602
rect 76564 3538 76616 3544
rect 74724 3528 74776 3534
rect 74724 3470 74776 3476
rect 76196 3528 76248 3534
rect 76196 3470 76248 3476
rect 75000 3052 75052 3058
rect 75000 2994 75052 3000
rect 75012 480 75040 2994
rect 76208 480 76236 3470
rect 76668 3058 76696 57598
rect 76944 56710 76972 60044
rect 77312 57526 77340 60044
rect 77588 57594 77616 60044
rect 77864 57730 77892 60044
rect 77852 57724 77904 57730
rect 77852 57666 77904 57672
rect 77576 57588 77628 57594
rect 77576 57530 77628 57536
rect 77300 57520 77352 57526
rect 77300 57462 77352 57468
rect 77208 57452 77260 57458
rect 77208 57394 77260 57400
rect 76932 56704 76984 56710
rect 76932 56646 76984 56652
rect 77220 3534 77248 57394
rect 78140 56914 78168 60044
rect 78416 57662 78444 60044
rect 78404 57656 78456 57662
rect 78404 57598 78456 57604
rect 78692 57458 78720 60044
rect 78784 60030 79074 60058
rect 79152 60030 79350 60058
rect 79428 60030 79626 60058
rect 78680 57452 78732 57458
rect 78680 57394 78732 57400
rect 78128 56908 78180 56914
rect 78128 56850 78180 56856
rect 78784 3602 78812 60030
rect 79152 57644 79180 60030
rect 78876 57616 79180 57644
rect 77392 3596 77444 3602
rect 77392 3538 77444 3544
rect 78772 3596 78824 3602
rect 78772 3538 78824 3544
rect 77208 3528 77260 3534
rect 77208 3470 77260 3476
rect 76656 3052 76708 3058
rect 76656 2994 76708 3000
rect 77404 480 77432 3538
rect 78876 3482 78904 57616
rect 79428 45554 79456 60030
rect 79888 57050 79916 60044
rect 80164 57594 80192 60044
rect 80440 57798 80468 60044
rect 80428 57792 80480 57798
rect 80428 57734 80480 57740
rect 80152 57588 80204 57594
rect 80152 57530 80204 57536
rect 80808 57526 80836 60044
rect 81098 60030 81204 60058
rect 81072 57656 81124 57662
rect 81072 57598 81124 57604
rect 80796 57520 80848 57526
rect 80796 57462 80848 57468
rect 79876 57044 79928 57050
rect 79876 56986 79928 56992
rect 80428 57044 80480 57050
rect 80428 56986 80480 56992
rect 79152 45526 79456 45554
rect 79152 3534 79180 45526
rect 80440 16574 80468 56986
rect 80440 16546 80928 16574
rect 78600 3454 78904 3482
rect 79140 3528 79192 3534
rect 79140 3470 79192 3476
rect 79692 3528 79744 3534
rect 79692 3470 79744 3476
rect 78600 480 78628 3454
rect 79704 480 79732 3470
rect 80900 480 80928 16546
rect 81084 2854 81112 57598
rect 81176 3738 81204 60030
rect 81360 57662 81388 60044
rect 81348 57656 81400 57662
rect 81348 57598 81400 57604
rect 81256 57588 81308 57594
rect 81256 57530 81308 57536
rect 81164 3732 81216 3738
rect 81164 3674 81216 3680
rect 81268 2922 81296 57530
rect 81348 57520 81400 57526
rect 81348 57462 81400 57468
rect 81360 3534 81388 57462
rect 81636 57458 81664 60044
rect 81912 57730 81940 60044
rect 81900 57724 81952 57730
rect 81900 57666 81952 57672
rect 81624 57452 81676 57458
rect 81624 57394 81676 57400
rect 82188 57322 82216 60044
rect 82570 60030 82676 60058
rect 82176 57316 82228 57322
rect 82176 57258 82228 57264
rect 81348 3528 81400 3534
rect 81348 3470 81400 3476
rect 82648 3466 82676 60030
rect 82832 57526 82860 60044
rect 83004 57792 83056 57798
rect 83004 57734 83056 57740
rect 82820 57520 82872 57526
rect 82820 57462 82872 57468
rect 82728 57452 82780 57458
rect 82728 57394 82780 57400
rect 82740 3602 82768 57394
rect 83016 16574 83044 57734
rect 83108 57458 83136 60044
rect 83384 57594 83412 60044
rect 83674 60030 83872 60058
rect 83740 57792 83792 57798
rect 83740 57734 83792 57740
rect 83372 57588 83424 57594
rect 83372 57530 83424 57536
rect 83096 57452 83148 57458
rect 83096 57394 83148 57400
rect 83752 57254 83780 57734
rect 83844 57644 83872 60030
rect 83936 57798 83964 60044
rect 83924 57792 83976 57798
rect 83924 57734 83976 57740
rect 83844 57616 84056 57644
rect 83924 57520 83976 57526
rect 83924 57462 83976 57468
rect 83740 57248 83792 57254
rect 83740 57190 83792 57196
rect 83016 16546 83320 16574
rect 82728 3596 82780 3602
rect 82728 3538 82780 3544
rect 82636 3460 82688 3466
rect 82636 3402 82688 3408
rect 81256 2916 81308 2922
rect 81256 2858 81308 2864
rect 82084 2916 82136 2922
rect 82084 2858 82136 2864
rect 81072 2848 81124 2854
rect 81072 2790 81124 2796
rect 82096 480 82124 2858
rect 83292 480 83320 16546
rect 83936 2922 83964 57462
rect 84028 4146 84056 57616
rect 84108 57588 84160 57594
rect 84108 57530 84160 57536
rect 84016 4140 84068 4146
rect 84016 4082 84068 4088
rect 84120 2990 84148 57530
rect 84304 57526 84332 60044
rect 84580 57934 84608 60044
rect 84568 57928 84620 57934
rect 84568 57870 84620 57876
rect 84292 57520 84344 57526
rect 84292 57462 84344 57468
rect 84856 56778 84884 60044
rect 85146 60030 85344 60058
rect 85316 57644 85344 60030
rect 85408 57866 85436 60044
rect 85396 57860 85448 57866
rect 85396 57802 85448 57808
rect 85316 57616 85528 57644
rect 85396 57520 85448 57526
rect 85396 57462 85448 57468
rect 84844 56772 84896 56778
rect 84844 56714 84896 56720
rect 85408 4078 85436 57462
rect 85396 4072 85448 4078
rect 85396 4014 85448 4020
rect 84476 3528 84528 3534
rect 84476 3470 84528 3476
rect 84108 2984 84160 2990
rect 84108 2926 84160 2932
rect 83924 2916 83976 2922
rect 83924 2858 83976 2864
rect 84488 480 84516 3470
rect 85500 3058 85528 57616
rect 85684 57526 85712 60044
rect 86052 57594 86080 60044
rect 86328 57798 86356 60044
rect 86316 57792 86368 57798
rect 86316 57734 86368 57740
rect 86604 57662 86632 60044
rect 86788 60030 86894 60058
rect 86592 57656 86644 57662
rect 86592 57598 86644 57604
rect 86040 57588 86092 57594
rect 86040 57530 86092 57536
rect 86684 57588 86736 57594
rect 86684 57530 86736 57536
rect 85672 57520 85724 57526
rect 85672 57462 85724 57468
rect 86592 57520 86644 57526
rect 86592 57462 86644 57468
rect 86224 56772 86276 56778
rect 86224 56714 86276 56720
rect 86236 9042 86264 56714
rect 86224 9036 86276 9042
rect 86224 8978 86276 8984
rect 86604 8974 86632 57462
rect 86592 8968 86644 8974
rect 86592 8910 86644 8916
rect 85672 3732 85724 3738
rect 85672 3674 85724 3680
rect 85488 3052 85540 3058
rect 85488 2994 85540 3000
rect 85684 480 85712 3674
rect 86696 3126 86724 57530
rect 86788 3262 86816 60030
rect 86868 57656 86920 57662
rect 86868 57598 86920 57604
rect 86776 3256 86828 3262
rect 86776 3198 86828 3204
rect 86880 3194 86908 57598
rect 87156 57390 87184 60044
rect 87432 57662 87460 60044
rect 87814 60030 88012 60058
rect 88090 60030 88288 60058
rect 87604 57724 87656 57730
rect 87604 57666 87656 57672
rect 87420 57656 87472 57662
rect 87420 57598 87472 57604
rect 87144 57384 87196 57390
rect 87144 57326 87196 57332
rect 87616 3534 87644 57666
rect 87984 55214 88012 60030
rect 88156 57656 88208 57662
rect 88156 57598 88208 57604
rect 87984 55186 88104 55214
rect 87972 3596 88024 3602
rect 87972 3538 88024 3544
rect 87604 3528 87656 3534
rect 87604 3470 87656 3476
rect 86868 3188 86920 3194
rect 86868 3130 86920 3136
rect 86684 3120 86736 3126
rect 86684 3062 86736 3068
rect 86868 2848 86920 2854
rect 86868 2790 86920 2796
rect 86880 480 86908 2790
rect 87984 480 88012 3538
rect 88076 3398 88104 55186
rect 88064 3392 88116 3398
rect 88064 3334 88116 3340
rect 88168 3330 88196 57598
rect 88260 4010 88288 60030
rect 88352 57594 88380 60044
rect 88628 57662 88656 60044
rect 88616 57656 88668 57662
rect 88616 57598 88668 57604
rect 88340 57588 88392 57594
rect 88340 57530 88392 57536
rect 88904 57050 88932 60044
rect 88892 57044 88944 57050
rect 88892 56986 88944 56992
rect 89180 56846 89208 60044
rect 89456 60030 89562 60058
rect 89352 57656 89404 57662
rect 89352 57598 89404 57604
rect 89168 56840 89220 56846
rect 89168 56782 89220 56788
rect 88248 4004 88300 4010
rect 88248 3946 88300 3952
rect 89364 3806 89392 57598
rect 89352 3800 89404 3806
rect 89352 3742 89404 3748
rect 89456 3738 89484 60030
rect 89628 57588 89680 57594
rect 89628 57530 89680 57536
rect 89536 56840 89588 56846
rect 89536 56782 89588 56788
rect 89548 3874 89576 56782
rect 89640 3942 89668 57530
rect 89824 57186 89852 60044
rect 89812 57180 89864 57186
rect 89812 57122 89864 57128
rect 90100 56710 90128 60044
rect 90390 60030 90588 60058
rect 90666 60030 90956 60058
rect 90560 57644 90588 60030
rect 90560 57616 90864 57644
rect 90180 57316 90232 57322
rect 90180 57258 90232 57264
rect 90088 56704 90140 56710
rect 90088 56646 90140 56652
rect 90192 16574 90220 57258
rect 90732 56840 90784 56846
rect 90732 56782 90784 56788
rect 90192 16546 90404 16574
rect 89628 3936 89680 3942
rect 89628 3878 89680 3884
rect 89536 3868 89588 3874
rect 89536 3810 89588 3816
rect 89444 3732 89496 3738
rect 89444 3674 89496 3680
rect 89168 3528 89220 3534
rect 89168 3470 89220 3476
rect 88156 3324 88208 3330
rect 88156 3266 88208 3272
rect 89180 480 89208 3470
rect 90376 480 90404 16546
rect 90744 15910 90772 56782
rect 90732 15904 90784 15910
rect 90732 15846 90784 15852
rect 90836 3602 90864 57616
rect 90824 3596 90876 3602
rect 90824 3538 90876 3544
rect 90928 3534 90956 60030
rect 91020 56846 91048 60044
rect 91296 57662 91324 60044
rect 91284 57656 91336 57662
rect 91284 57598 91336 57604
rect 91572 56846 91600 60044
rect 91848 57322 91876 60044
rect 92138 60030 92244 60058
rect 91836 57316 91888 57322
rect 91836 57258 91888 57264
rect 91008 56840 91060 56846
rect 91008 56782 91060 56788
rect 91560 56840 91612 56846
rect 91560 56782 91612 56788
rect 91008 56704 91060 56710
rect 91008 56646 91060 56652
rect 91020 3670 91048 56646
rect 92216 6186 92244 60030
rect 92296 57656 92348 57662
rect 92296 57598 92348 57604
rect 92204 6180 92256 6186
rect 92204 6122 92256 6128
rect 92308 4282 92336 57598
rect 92296 4276 92348 4282
rect 92296 4218 92348 4224
rect 91008 3664 91060 3670
rect 91008 3606 91060 3612
rect 90916 3528 90968 3534
rect 90916 3470 90968 3476
rect 92400 3466 92428 60044
rect 92768 57662 92796 60044
rect 93058 60030 93256 60058
rect 92848 57928 92900 57934
rect 92848 57870 92900 57876
rect 92756 57656 92808 57662
rect 92756 57598 92808 57604
rect 92860 57594 92888 57870
rect 92848 57588 92900 57594
rect 92848 57530 92900 57536
rect 93124 57452 93176 57458
rect 93124 57394 93176 57400
rect 93136 8362 93164 57394
rect 93228 55214 93256 60030
rect 93320 56914 93348 60044
rect 93610 60030 93808 60058
rect 93676 57656 93728 57662
rect 93676 57598 93728 57604
rect 93308 56908 93360 56914
rect 93308 56850 93360 56856
rect 93228 55186 93624 55214
rect 93124 8356 93176 8362
rect 93124 8298 93176 8304
rect 93596 8022 93624 55186
rect 93584 8016 93636 8022
rect 93584 7958 93636 7964
rect 93688 4350 93716 57598
rect 93780 4418 93808 60030
rect 93872 57526 93900 60044
rect 94148 57866 94176 60044
rect 94530 60030 94728 60058
rect 94806 60030 95004 60058
rect 94136 57860 94188 57866
rect 94136 57802 94188 57808
rect 94504 57588 94556 57594
rect 94504 57530 94556 57536
rect 93860 57520 93912 57526
rect 93860 57462 93912 57468
rect 93952 57384 94004 57390
rect 93952 57326 94004 57332
rect 93964 56982 93992 57326
rect 93952 56976 94004 56982
rect 93952 56918 94004 56924
rect 93952 8356 94004 8362
rect 93952 8298 94004 8304
rect 93768 4412 93820 4418
rect 93768 4354 93820 4360
rect 93676 4344 93728 4350
rect 93676 4286 93728 4292
rect 91560 3460 91612 3466
rect 91560 3402 91612 3408
rect 92388 3460 92440 3466
rect 92388 3402 92440 3408
rect 91572 480 91600 3402
rect 92756 2916 92808 2922
rect 92756 2858 92808 2864
rect 92768 480 92796 2858
rect 93964 480 93992 8298
rect 94516 4078 94544 57530
rect 94596 57384 94648 57390
rect 94596 57326 94648 57332
rect 94608 56846 94636 57326
rect 94700 56846 94728 60030
rect 94976 57610 95004 60030
rect 95068 57934 95096 60044
rect 95056 57928 95108 57934
rect 95056 57870 95108 57876
rect 94976 57582 95188 57610
rect 95056 57520 95108 57526
rect 95056 57462 95108 57468
rect 94596 56840 94648 56846
rect 94596 56782 94648 56788
rect 94688 56840 94740 56846
rect 94688 56782 94740 56788
rect 95068 7954 95096 57462
rect 95056 7948 95108 7954
rect 95056 7890 95108 7896
rect 95160 7886 95188 57582
rect 95344 57526 95372 60044
rect 95620 57662 95648 60044
rect 95896 57798 95924 60044
rect 96172 60030 96278 60058
rect 95884 57792 95936 57798
rect 95884 57734 95936 57740
rect 95608 57656 95660 57662
rect 95608 57598 95660 57604
rect 95332 57520 95384 57526
rect 95332 57462 95384 57468
rect 96172 57118 96200 60030
rect 96540 57746 96568 60044
rect 96816 57866 96844 60044
rect 96712 57860 96764 57866
rect 96712 57802 96764 57808
rect 96804 57860 96856 57866
rect 96804 57802 96856 57808
rect 96264 57718 96568 57746
rect 96160 57112 96212 57118
rect 96160 57054 96212 57060
rect 95148 7880 95200 7886
rect 95148 7822 95200 7828
rect 96264 7750 96292 57718
rect 96344 57656 96396 57662
rect 96344 57598 96396 57604
rect 96356 7818 96384 57598
rect 96724 57526 96752 57802
rect 97092 57662 97120 60044
rect 97382 60030 97580 60058
rect 97080 57656 97132 57662
rect 97080 57598 97132 57604
rect 97264 57588 97316 57594
rect 97264 57530 97316 57536
rect 96436 57520 96488 57526
rect 96436 57462 96488 57468
rect 96712 57520 96764 57526
rect 96712 57462 96764 57468
rect 96344 7812 96396 7818
rect 96344 7754 96396 7760
rect 96252 7744 96304 7750
rect 96252 7686 96304 7692
rect 96448 4486 96476 57462
rect 96712 57248 96764 57254
rect 96712 57190 96764 57196
rect 96528 57112 96580 57118
rect 96528 57054 96580 57060
rect 96540 4622 96568 57054
rect 96724 16574 96752 57190
rect 96724 16546 97212 16574
rect 96528 4616 96580 4622
rect 96528 4558 96580 4564
rect 96436 4480 96488 4486
rect 96436 4422 96488 4428
rect 96252 4140 96304 4146
rect 96252 4082 96304 4088
rect 94412 4072 94464 4078
rect 94412 4014 94464 4020
rect 94504 4072 94556 4078
rect 94504 4014 94556 4020
rect 94424 2922 94452 4014
rect 95148 2984 95200 2990
rect 95148 2926 95200 2932
rect 94412 2916 94464 2922
rect 94412 2858 94464 2864
rect 95160 480 95188 2926
rect 96264 480 96292 4082
rect 97184 3482 97212 16546
rect 97276 4146 97304 57530
rect 97552 55214 97580 60030
rect 97644 56642 97672 60044
rect 98012 56710 98040 60044
rect 98288 57118 98316 60044
rect 98564 57662 98592 60044
rect 98552 57656 98604 57662
rect 98552 57598 98604 57604
rect 98276 57112 98328 57118
rect 98276 57054 98328 57060
rect 98840 56778 98868 60044
rect 98932 60030 99130 60058
rect 98828 56772 98880 56778
rect 98828 56714 98880 56720
rect 98000 56704 98052 56710
rect 98000 56646 98052 56652
rect 97632 56636 97684 56642
rect 97632 56578 97684 56584
rect 97552 55186 97948 55214
rect 97920 7682 97948 55186
rect 98932 9382 98960 60030
rect 99288 57656 99340 57662
rect 99288 57598 99340 57604
rect 99012 57112 99064 57118
rect 99012 57054 99064 57060
rect 99104 57112 99156 57118
rect 99104 57054 99156 57060
rect 98920 9376 98972 9382
rect 98920 9318 98972 9324
rect 97908 7676 97960 7682
rect 97908 7618 97960 7624
rect 99024 7614 99052 57054
rect 99116 56846 99144 57054
rect 99104 56840 99156 56846
rect 99104 56782 99156 56788
rect 99196 56772 99248 56778
rect 99196 56714 99248 56720
rect 99104 56704 99156 56710
rect 99104 56646 99156 56652
rect 99012 7608 99064 7614
rect 99012 7550 99064 7556
rect 99116 4554 99144 56646
rect 99208 4690 99236 56714
rect 99196 4684 99248 4690
rect 99196 4626 99248 4632
rect 99104 4548 99156 4554
rect 99104 4490 99156 4496
rect 99300 4214 99328 57598
rect 99392 56778 99420 60044
rect 99760 56846 99788 60044
rect 100036 57662 100064 60044
rect 100326 60030 100524 60058
rect 100024 57656 100076 57662
rect 100024 57598 100076 57604
rect 99748 56840 99800 56846
rect 99748 56782 99800 56788
rect 99380 56772 99432 56778
rect 99380 56714 99432 56720
rect 100496 9314 100524 60030
rect 100588 57934 100616 60044
rect 100576 57928 100628 57934
rect 100576 57870 100628 57876
rect 100576 57656 100628 57662
rect 100576 57598 100628 57604
rect 100484 9308 100536 9314
rect 100484 9250 100536 9256
rect 100588 4758 100616 57598
rect 100864 57526 100892 60044
rect 101140 57662 101168 60044
rect 101508 57798 101536 60044
rect 101798 60030 101996 60058
rect 101496 57792 101548 57798
rect 101496 57734 101548 57740
rect 101588 57724 101640 57730
rect 101588 57666 101640 57672
rect 101772 57724 101824 57730
rect 101772 57666 101824 57672
rect 101128 57656 101180 57662
rect 101128 57598 101180 57604
rect 100760 57520 100812 57526
rect 100760 57462 100812 57468
rect 100852 57520 100904 57526
rect 100852 57462 100904 57468
rect 100772 56778 100800 57462
rect 101600 57458 101628 57666
rect 101404 57452 101456 57458
rect 101404 57394 101456 57400
rect 101588 57452 101640 57458
rect 101588 57394 101640 57400
rect 100668 56772 100720 56778
rect 100668 56714 100720 56720
rect 100760 56772 100812 56778
rect 100760 56714 100812 56720
rect 100576 4752 100628 4758
rect 100576 4694 100628 4700
rect 99288 4208 99340 4214
rect 99288 4150 99340 4156
rect 97264 4140 97316 4146
rect 97264 4082 97316 4088
rect 100680 4078 100708 56714
rect 101036 9036 101088 9042
rect 101036 8978 101088 8984
rect 99840 4072 99892 4078
rect 99840 4014 99892 4020
rect 100668 4072 100720 4078
rect 100668 4014 100720 4020
rect 97184 3454 97488 3482
rect 97460 480 97488 3454
rect 98644 2916 98696 2922
rect 98644 2858 98696 2864
rect 98656 480 98684 2858
rect 99852 480 99880 4014
rect 101048 480 101076 8978
rect 101416 2854 101444 57394
rect 101784 9178 101812 57666
rect 101864 57656 101916 57662
rect 101864 57598 101916 57604
rect 101968 57610 101996 60030
rect 102060 57730 102088 60044
rect 102140 57996 102192 58002
rect 102140 57938 102192 57944
rect 102048 57724 102100 57730
rect 102048 57666 102100 57672
rect 101876 9246 101904 57598
rect 101968 57582 102088 57610
rect 101956 57520 102008 57526
rect 101956 57462 102008 57468
rect 101864 9240 101916 9246
rect 101864 9182 101916 9188
rect 101772 9172 101824 9178
rect 101772 9114 101824 9120
rect 101968 5506 101996 57462
rect 101956 5500 102008 5506
rect 101956 5442 102008 5448
rect 102060 5438 102088 57582
rect 102152 57526 102180 57938
rect 102336 57730 102364 60044
rect 102324 57724 102376 57730
rect 102324 57666 102376 57672
rect 102140 57520 102192 57526
rect 102140 57462 102192 57468
rect 102612 56710 102640 60044
rect 102902 60030 103192 60058
rect 103060 57588 103112 57594
rect 103060 57530 103112 57536
rect 103072 57497 103100 57530
rect 103058 57488 103114 57497
rect 103058 57423 103114 57432
rect 102876 57044 102928 57050
rect 102876 56986 102928 56992
rect 103060 57044 103112 57050
rect 103060 56986 103112 56992
rect 102784 56976 102836 56982
rect 102784 56918 102836 56924
rect 102600 56704 102652 56710
rect 102600 56646 102652 56652
rect 102048 5432 102100 5438
rect 102048 5374 102100 5380
rect 102232 3052 102284 3058
rect 102232 2994 102284 3000
rect 101404 2848 101456 2854
rect 101404 2790 101456 2796
rect 102244 480 102272 2994
rect 102796 2922 102824 56918
rect 102888 2990 102916 56986
rect 103072 56778 103100 56986
rect 103060 56772 103112 56778
rect 103060 56714 103112 56720
rect 103164 55214 103192 60030
rect 103256 57662 103284 60044
rect 103546 60030 103744 60058
rect 103244 57656 103296 57662
rect 103244 57598 103296 57604
rect 103518 57488 103574 57497
rect 103518 57423 103574 57432
rect 103532 57186 103560 57423
rect 103612 57384 103664 57390
rect 103612 57326 103664 57332
rect 103520 57180 103572 57186
rect 103520 57122 103572 57128
rect 103624 56778 103652 57326
rect 103716 57118 103744 60030
rect 103808 57390 103836 60044
rect 103796 57384 103848 57390
rect 103796 57326 103848 57332
rect 103704 57112 103756 57118
rect 103704 57054 103756 57060
rect 103612 56772 103664 56778
rect 103612 56714 103664 56720
rect 104084 56710 104112 60044
rect 104360 57594 104388 60044
rect 104348 57588 104400 57594
rect 104348 57530 104400 57536
rect 104532 57384 104584 57390
rect 104532 57326 104584 57332
rect 104164 57248 104216 57254
rect 104164 57190 104216 57196
rect 103336 56704 103388 56710
rect 104072 56704 104124 56710
rect 103388 56664 103468 56692
rect 103336 56646 103388 56652
rect 103164 55186 103376 55214
rect 103348 9110 103376 55186
rect 103336 9104 103388 9110
rect 103336 9046 103388 9052
rect 103440 5370 103468 56664
rect 104072 56646 104124 56652
rect 103428 5364 103480 5370
rect 103428 5306 103480 5312
rect 103336 4140 103388 4146
rect 103336 4082 103388 4088
rect 102876 2984 102928 2990
rect 102876 2926 102928 2932
rect 102784 2916 102836 2922
rect 102784 2858 102836 2864
rect 103348 480 103376 4082
rect 104176 3058 104204 57190
rect 104544 16574 104572 57326
rect 104452 16546 104572 16574
rect 104452 9042 104480 16546
rect 104440 9036 104492 9042
rect 104440 8978 104492 8984
rect 104636 8974 104664 60044
rect 104716 57588 104768 57594
rect 104716 57530 104768 57536
rect 104532 8968 104584 8974
rect 104532 8910 104584 8916
rect 104624 8968 104676 8974
rect 104624 8910 104676 8916
rect 104164 3052 104216 3058
rect 104164 2994 104216 3000
rect 104544 480 104572 8910
rect 104728 5234 104756 57530
rect 105004 57254 105032 60044
rect 104992 57248 105044 57254
rect 104992 57190 105044 57196
rect 104808 57112 104860 57118
rect 104808 57054 104860 57060
rect 105176 57112 105228 57118
rect 105176 57054 105228 57060
rect 104820 5302 104848 57054
rect 105188 56846 105216 57054
rect 105280 56846 105308 60044
rect 105570 60030 105768 60058
rect 105176 56840 105228 56846
rect 105176 56782 105228 56788
rect 105268 56840 105320 56846
rect 105268 56782 105320 56788
rect 105544 56772 105596 56778
rect 105544 56714 105596 56720
rect 105556 6254 105584 56714
rect 105740 55214 105768 60030
rect 105832 57390 105860 60044
rect 105820 57384 105872 57390
rect 105820 57326 105872 57332
rect 105740 55186 106044 55214
rect 106016 10946 106044 55186
rect 106004 10940 106056 10946
rect 106004 10882 106056 10888
rect 105544 6248 105596 6254
rect 105544 6190 105596 6196
rect 104808 5296 104860 5302
rect 104808 5238 104860 5244
rect 104716 5228 104768 5234
rect 104716 5170 104768 5176
rect 106108 5098 106136 60044
rect 106292 60030 106490 60058
rect 106188 56840 106240 56846
rect 106188 56782 106240 56788
rect 106200 5166 106228 56782
rect 106292 45554 106320 60030
rect 106752 57594 106780 60044
rect 107042 60030 107240 60058
rect 107318 60030 107424 60058
rect 106740 57588 106792 57594
rect 106740 57530 106792 57536
rect 106372 56772 106424 56778
rect 106372 56714 106424 56720
rect 106384 50386 106412 56714
rect 107212 55214 107240 60030
rect 107212 55186 107332 55214
rect 106372 50380 106424 50386
rect 106372 50322 106424 50328
rect 106292 45526 107240 45554
rect 107212 10878 107240 45526
rect 107200 10872 107252 10878
rect 107200 10814 107252 10820
rect 107304 10810 107332 55186
rect 107292 10804 107344 10810
rect 107292 10746 107344 10752
rect 107396 10742 107424 60030
rect 107476 57588 107528 57594
rect 107476 57530 107528 57536
rect 107384 10736 107436 10742
rect 107384 10678 107436 10684
rect 106188 5160 106240 5166
rect 106188 5102 106240 5108
rect 106096 5092 106148 5098
rect 106096 5034 106148 5040
rect 107488 5030 107516 57530
rect 107580 56778 107608 60044
rect 107856 56846 107884 60044
rect 108238 60030 108436 60058
rect 108212 57588 108264 57594
rect 108212 57530 108264 57536
rect 108224 57254 108252 57530
rect 108212 57248 108264 57254
rect 108212 57190 108264 57196
rect 108304 57248 108356 57254
rect 108304 57190 108356 57196
rect 107844 56840 107896 56846
rect 107844 56782 107896 56788
rect 107568 56772 107620 56778
rect 107568 56714 107620 56720
rect 107660 56772 107712 56778
rect 107660 56714 107712 56720
rect 107672 50386 107700 56714
rect 108316 56642 108344 57190
rect 108304 56636 108356 56642
rect 108304 56578 108356 56584
rect 108408 55214 108436 60030
rect 108500 56778 108528 60044
rect 108790 60030 108896 60058
rect 108764 56840 108816 56846
rect 108764 56782 108816 56788
rect 108488 56772 108540 56778
rect 108488 56714 108540 56720
rect 108408 55186 108712 55214
rect 107568 50380 107620 50386
rect 107568 50322 107620 50328
rect 107660 50380 107712 50386
rect 107660 50322 107712 50328
rect 107476 5024 107528 5030
rect 107476 4966 107528 4972
rect 107580 4962 107608 50322
rect 108684 10606 108712 55186
rect 108776 10674 108804 56782
rect 108764 10668 108816 10674
rect 108764 10610 108816 10616
rect 108672 10600 108724 10606
rect 108672 10542 108724 10548
rect 108868 10538 108896 60030
rect 109052 50386 109080 60044
rect 109328 56642 109356 60044
rect 109618 60030 109908 60058
rect 109986 60030 110184 60058
rect 109316 56636 109368 56642
rect 109316 56578 109368 56584
rect 109880 51074 109908 60030
rect 110156 51074 110184 60030
rect 110248 56846 110276 60044
rect 110236 56840 110288 56846
rect 110236 56782 110288 56788
rect 110524 56642 110552 60044
rect 110800 56710 110828 60044
rect 110788 56704 110840 56710
rect 110788 56646 110840 56652
rect 110328 56636 110380 56642
rect 110328 56578 110380 56584
rect 110512 56636 110564 56642
rect 110512 56578 110564 56584
rect 109880 51046 110092 51074
rect 110156 51046 110276 51074
rect 108948 50380 109000 50386
rect 108948 50322 109000 50328
rect 109040 50380 109092 50386
rect 109040 50322 109092 50328
rect 108856 10532 108908 10538
rect 108856 10474 108908 10480
rect 107568 4956 107620 4962
rect 107568 4898 107620 4904
rect 108960 4894 108988 50322
rect 110064 10334 110092 51046
rect 110144 50380 110196 50386
rect 110144 50322 110196 50328
rect 110156 10470 110184 50322
rect 110144 10464 110196 10470
rect 110144 10406 110196 10412
rect 110248 10402 110276 51046
rect 110236 10396 110288 10402
rect 110236 10338 110288 10344
rect 110052 10328 110104 10334
rect 110052 10270 110104 10276
rect 108948 4888 109000 4894
rect 108948 4830 109000 4836
rect 110340 4826 110368 56578
rect 111076 55486 111104 60044
rect 111366 60030 111472 60058
rect 111064 55480 111116 55486
rect 111064 55422 111116 55428
rect 111444 9858 111472 60030
rect 111536 60030 111734 60058
rect 111536 15366 111564 60030
rect 111616 56636 111668 56642
rect 111616 56578 111668 56584
rect 111524 15360 111576 15366
rect 111524 15302 111576 15308
rect 111432 9852 111484 9858
rect 111432 9794 111484 9800
rect 111628 9790 111656 56578
rect 111996 55418 112024 60044
rect 112272 56642 112300 60044
rect 112562 60030 112760 60058
rect 112260 56636 112312 56642
rect 112260 56578 112312 56584
rect 111984 55412 112036 55418
rect 111984 55354 112036 55360
rect 112732 55350 112760 60030
rect 112824 55826 112852 60044
rect 112916 60030 113114 60058
rect 112812 55820 112864 55826
rect 112812 55762 112864 55768
rect 112916 55706 112944 60030
rect 113468 56710 113496 60044
rect 113758 60030 113956 60058
rect 114034 60030 114232 60058
rect 113928 57746 113956 60030
rect 113928 57718 114140 57746
rect 113732 57588 113784 57594
rect 113732 57530 113784 57536
rect 113824 57588 113876 57594
rect 113824 57530 113876 57536
rect 113744 56846 113772 57530
rect 113836 57458 113864 57530
rect 113824 57452 113876 57458
rect 113824 57394 113876 57400
rect 113916 57452 113968 57458
rect 113916 57394 113968 57400
rect 113640 56840 113692 56846
rect 113640 56782 113692 56788
rect 113732 56840 113784 56846
rect 113732 56782 113784 56788
rect 113456 56704 113508 56710
rect 113456 56646 113508 56652
rect 112996 56636 113048 56642
rect 112996 56578 113048 56584
rect 112824 55678 112944 55706
rect 112720 55344 112772 55350
rect 112720 55286 112772 55292
rect 112824 9994 112852 55678
rect 112904 55344 112956 55350
rect 112904 55286 112956 55292
rect 112916 15434 112944 55286
rect 112904 15428 112956 15434
rect 112904 15370 112956 15376
rect 112812 9988 112864 9994
rect 112812 9930 112864 9936
rect 113008 9926 113036 56578
rect 113652 56506 113680 56782
rect 113928 56778 113956 57394
rect 114112 56778 114140 57718
rect 113916 56772 113968 56778
rect 113916 56714 113968 56720
rect 114100 56772 114152 56778
rect 114100 56714 114152 56720
rect 114204 56642 114232 60030
rect 114192 56636 114244 56642
rect 114192 56578 114244 56584
rect 113640 56500 113692 56506
rect 113640 56442 113692 56448
rect 114296 15570 114324 60044
rect 114376 56704 114428 56710
rect 114376 56646 114428 56652
rect 114284 15564 114336 15570
rect 114284 15506 114336 15512
rect 114388 15502 114416 56646
rect 114468 56636 114520 56642
rect 114468 56578 114520 56584
rect 114376 15496 114428 15502
rect 114376 15438 114428 15444
rect 114480 10062 114508 56578
rect 114572 55622 114600 60044
rect 114848 56642 114876 60044
rect 115216 56710 115244 60044
rect 115506 60030 115704 60058
rect 115782 60030 115888 60058
rect 115204 56704 115256 56710
rect 115204 56646 115256 56652
rect 114836 56636 114888 56642
rect 114836 56578 114888 56584
rect 115572 56636 115624 56642
rect 115572 56578 115624 56584
rect 114560 55616 114612 55622
rect 114560 55558 114612 55564
rect 115584 10130 115612 56578
rect 115676 18902 115704 60030
rect 115756 56704 115808 56710
rect 115756 56646 115808 56652
rect 115664 18896 115716 18902
rect 115664 18838 115716 18844
rect 115768 15638 115796 56646
rect 115860 52902 115888 60030
rect 116044 56710 116072 60044
rect 116032 56704 116084 56710
rect 116032 56646 116084 56652
rect 116320 55690 116348 60044
rect 116308 55684 116360 55690
rect 116308 55626 116360 55632
rect 116596 52970 116624 60044
rect 116978 60030 117084 60058
rect 116858 57080 116914 57089
rect 116858 57015 116914 57024
rect 116872 56642 116900 57015
rect 116860 56636 116912 56642
rect 116860 56578 116912 56584
rect 116952 56636 117004 56642
rect 116952 56578 117004 56584
rect 116584 52964 116636 52970
rect 116584 52906 116636 52912
rect 115848 52896 115900 52902
rect 115848 52838 115900 52844
rect 115756 15632 115808 15638
rect 115756 15574 115808 15580
rect 115572 10124 115624 10130
rect 115572 10066 115624 10072
rect 114468 10056 114520 10062
rect 114468 9998 114520 10004
rect 112996 9920 113048 9926
rect 112996 9862 113048 9868
rect 111616 9784 111668 9790
rect 111616 9726 111668 9732
rect 116964 5574 116992 56578
rect 117056 15774 117084 60030
rect 117136 56704 117188 56710
rect 117136 56646 117188 56652
rect 117044 15768 117096 15774
rect 117044 15710 117096 15716
rect 117148 15706 117176 56646
rect 117240 56642 117268 60044
rect 117320 57384 117372 57390
rect 117320 57326 117372 57332
rect 117228 56636 117280 56642
rect 117228 56578 117280 56584
rect 117332 56438 117360 57326
rect 117516 56681 117544 60044
rect 117608 60030 117806 60058
rect 118082 60030 118280 60058
rect 117502 56672 117558 56681
rect 117502 56607 117558 56616
rect 117320 56432 117372 56438
rect 117320 56374 117372 56380
rect 117608 45554 117636 60030
rect 118252 51074 118280 60030
rect 118344 57225 118372 60044
rect 118608 57452 118660 57458
rect 118608 57394 118660 57400
rect 118516 57316 118568 57322
rect 118516 57258 118568 57264
rect 118330 57216 118386 57225
rect 118330 57151 118386 57160
rect 118528 56574 118556 57258
rect 118620 56953 118648 57394
rect 118606 56944 118662 56953
rect 118606 56879 118662 56888
rect 118606 56808 118662 56817
rect 118712 56778 118740 60044
rect 118896 60030 119002 60058
rect 118792 57452 118844 57458
rect 118792 57394 118844 57400
rect 118804 56817 118832 57394
rect 118790 56808 118846 56817
rect 118606 56743 118608 56752
rect 118660 56743 118662 56752
rect 118700 56772 118752 56778
rect 118608 56714 118660 56720
rect 118790 56743 118846 56752
rect 118700 56714 118752 56720
rect 118516 56568 118568 56574
rect 118516 56510 118568 56516
rect 118252 51046 118648 51074
rect 117608 45526 118556 45554
rect 118528 15842 118556 45526
rect 118516 15836 118568 15842
rect 118516 15778 118568 15784
rect 117136 15700 117188 15706
rect 117136 15642 117188 15648
rect 118620 5642 118648 51046
rect 118896 46238 118924 60030
rect 118976 57384 119028 57390
rect 118976 57326 119028 57332
rect 118988 57089 119016 57326
rect 118974 57080 119030 57089
rect 118974 57015 119030 57024
rect 119264 53038 119292 60044
rect 119356 60030 119554 60058
rect 119632 60030 119830 60058
rect 120198 60030 120396 60058
rect 119252 53032 119304 53038
rect 119252 52974 119304 52980
rect 118884 46232 118936 46238
rect 118884 46174 118936 46180
rect 119356 45422 119384 60030
rect 119632 46288 119660 60030
rect 120368 58002 120396 60030
rect 120356 57996 120408 58002
rect 120356 57938 120408 57944
rect 120460 57322 120488 60044
rect 120448 57316 120500 57322
rect 120448 57258 120500 57264
rect 120736 56778 120764 60044
rect 121012 57361 121040 60044
rect 120998 57352 121054 57361
rect 120998 57287 121054 57296
rect 121184 57316 121236 57322
rect 121184 57258 121236 57264
rect 119804 56772 119856 56778
rect 119804 56714 119856 56720
rect 120080 56772 120132 56778
rect 120080 56714 120132 56720
rect 120724 56772 120776 56778
rect 120724 56714 120776 56720
rect 119540 46260 119660 46288
rect 119344 45416 119396 45422
rect 119344 45358 119396 45364
rect 119540 38654 119568 46260
rect 119712 45416 119764 45422
rect 119712 45358 119764 45364
rect 119540 38626 119660 38654
rect 119632 5778 119660 38626
rect 119724 16522 119752 45358
rect 119816 16590 119844 56714
rect 120092 46238 120120 56714
rect 120724 56568 120776 56574
rect 120724 56510 120776 56516
rect 119896 46232 119948 46238
rect 119896 46174 119948 46180
rect 120080 46232 120132 46238
rect 120080 46174 120132 46180
rect 119804 16584 119856 16590
rect 119804 16526 119856 16532
rect 119712 16516 119764 16522
rect 119712 16458 119764 16464
rect 119620 5772 119672 5778
rect 119620 5714 119672 5720
rect 119908 5710 119936 46174
rect 119896 5704 119948 5710
rect 119896 5646 119948 5652
rect 118608 5636 118660 5642
rect 118608 5578 118660 5584
rect 116952 5568 117004 5574
rect 116952 5510 117004 5516
rect 110328 4820 110380 4826
rect 110328 4762 110380 4768
rect 114008 4004 114060 4010
rect 114008 3946 114060 3952
rect 112812 3392 112864 3398
rect 112812 3334 112864 3340
rect 111616 3324 111668 3330
rect 111616 3266 111668 3272
rect 109316 3256 109368 3262
rect 109316 3198 109368 3204
rect 108120 3188 108172 3194
rect 108120 3130 108172 3136
rect 105728 3120 105780 3126
rect 105728 3062 105780 3068
rect 105740 480 105768 3062
rect 106924 2848 106976 2854
rect 106924 2790 106976 2796
rect 106936 480 106964 2790
rect 108132 480 108160 3130
rect 109328 480 109356 3198
rect 110512 2916 110564 2922
rect 110512 2858 110564 2864
rect 110524 480 110552 2858
rect 111628 480 111656 3266
rect 112824 480 112852 3334
rect 114020 480 114048 3946
rect 115204 3936 115256 3942
rect 115204 3878 115256 3884
rect 115216 480 115244 3878
rect 118792 3868 118844 3874
rect 118792 3810 118844 3816
rect 116400 3800 116452 3806
rect 116400 3742 116452 3748
rect 116412 480 116440 3742
rect 117596 2984 117648 2990
rect 117596 2926 117648 2932
rect 117608 480 117636 2926
rect 118804 480 118832 3810
rect 120736 3738 120764 56510
rect 121196 16454 121224 57258
rect 121184 16448 121236 16454
rect 121184 16390 121236 16396
rect 121288 16386 121316 60044
rect 121578 60030 121684 60058
rect 121368 46232 121420 46238
rect 121368 46174 121420 46180
rect 121276 16380 121328 16386
rect 121276 16322 121328 16328
rect 121380 5846 121408 46174
rect 121656 41414 121684 60030
rect 121932 52426 121960 60044
rect 122024 60030 122222 60058
rect 122498 60030 122696 60058
rect 121920 52420 121972 52426
rect 121920 52362 121972 52368
rect 122024 51074 122052 60030
rect 122024 51046 122604 51074
rect 121656 41386 122420 41414
rect 122392 5914 122420 41386
rect 122576 16318 122604 51046
rect 122564 16312 122616 16318
rect 122564 16254 122616 16260
rect 122668 5982 122696 60030
rect 122760 52358 122788 60044
rect 122944 60030 123050 60058
rect 122840 57316 122892 57322
rect 122840 57258 122892 57264
rect 122748 52352 122800 52358
rect 122748 52294 122800 52300
rect 122852 46238 122880 57258
rect 122840 46232 122892 46238
rect 122840 46174 122892 46180
rect 122944 41414 122972 60030
rect 123312 57322 123340 60044
rect 123694 60030 123892 60058
rect 123300 57316 123352 57322
rect 123300 57258 123352 57264
rect 123300 56772 123352 56778
rect 123300 56714 123352 56720
rect 123312 46186 123340 56714
rect 123482 56672 123538 56681
rect 123482 56607 123538 56616
rect 123496 52834 123524 56607
rect 123484 52828 123536 52834
rect 123484 52770 123536 52776
rect 123864 51074 123892 60030
rect 123956 56778 123984 60044
rect 124246 60030 124352 60058
rect 123944 56772 123996 56778
rect 123944 56714 123996 56720
rect 123864 51046 124076 51074
rect 123312 46158 123984 46186
rect 122944 41386 123892 41414
rect 123864 16250 123892 41386
rect 123852 16244 123904 16250
rect 123852 16186 123904 16192
rect 123956 16182 123984 46158
rect 123944 16176 123996 16182
rect 123944 16118 123996 16124
rect 123576 15904 123628 15910
rect 123576 15846 123628 15852
rect 122656 5976 122708 5982
rect 122656 5918 122708 5924
rect 122380 5908 122432 5914
rect 122380 5850 122432 5856
rect 121368 5840 121420 5846
rect 121368 5782 121420 5788
rect 119896 3732 119948 3738
rect 119896 3674 119948 3680
rect 120724 3732 120776 3738
rect 120724 3674 120776 3680
rect 119908 480 119936 3674
rect 122288 3664 122340 3670
rect 122288 3606 122340 3612
rect 121092 3052 121144 3058
rect 121092 2994 121144 3000
rect 121104 480 121132 2994
rect 122300 480 122328 3606
rect 123484 3596 123536 3602
rect 123484 3538 123536 3544
rect 123496 480 123524 3538
rect 123588 3194 123616 15846
rect 124048 11218 124076 51046
rect 124128 46232 124180 46238
rect 124128 46174 124180 46180
rect 124036 11212 124088 11218
rect 124036 11154 124088 11160
rect 124140 6050 124168 46174
rect 124324 46170 124352 60030
rect 124404 57316 124456 57322
rect 124404 57258 124456 57264
rect 124416 46374 124444 57258
rect 124404 46368 124456 46374
rect 124404 46310 124456 46316
rect 124508 46238 124536 60044
rect 124798 60030 124996 60058
rect 124588 56772 124640 56778
rect 124588 56714 124640 56720
rect 124600 46306 124628 56714
rect 124968 51074 124996 60030
rect 125060 57322 125088 60044
rect 125048 57316 125100 57322
rect 125048 57258 125100 57264
rect 125428 56778 125456 60044
rect 125704 57322 125732 60044
rect 125796 60030 125994 60058
rect 125692 57316 125744 57322
rect 125692 57258 125744 57264
rect 125416 56772 125468 56778
rect 125416 56714 125468 56720
rect 125600 56772 125652 56778
rect 125600 56714 125652 56720
rect 124968 51046 125180 51074
rect 124588 46300 124640 46306
rect 124588 46242 124640 46248
rect 124496 46232 124548 46238
rect 124496 46174 124548 46180
rect 124312 46164 124364 46170
rect 124312 46106 124364 46112
rect 125152 17134 125180 51046
rect 125508 46368 125560 46374
rect 125508 46310 125560 46316
rect 125324 46300 125376 46306
rect 125324 46242 125376 46248
rect 125232 46232 125284 46238
rect 125232 46174 125284 46180
rect 125140 17128 125192 17134
rect 125140 17070 125192 17076
rect 125244 11286 125272 46174
rect 125336 11354 125364 46242
rect 125416 46164 125468 46170
rect 125416 46106 125468 46112
rect 125324 11348 125376 11354
rect 125324 11290 125376 11296
rect 125232 11280 125284 11286
rect 125232 11222 125284 11228
rect 125428 6118 125456 46106
rect 125520 6866 125548 46310
rect 125612 46238 125640 56714
rect 125796 46306 125824 60030
rect 126256 56778 126284 60044
rect 126334 56944 126390 56953
rect 126334 56879 126390 56888
rect 126348 56778 126376 56879
rect 126244 56772 126296 56778
rect 126244 56714 126296 56720
rect 126336 56772 126388 56778
rect 126336 56714 126388 56720
rect 125784 46300 125836 46306
rect 125784 46242 125836 46248
rect 125600 46232 125652 46238
rect 125600 46174 125652 46180
rect 126532 17950 126560 60044
rect 126612 57316 126664 57322
rect 126612 57258 126664 57264
rect 126520 17944 126572 17950
rect 126520 17886 126572 17892
rect 126624 17202 126652 57258
rect 126704 46232 126756 46238
rect 126704 46174 126756 46180
rect 126612 17196 126664 17202
rect 126612 17138 126664 17144
rect 126716 11422 126744 46174
rect 126704 11416 126756 11422
rect 126704 11358 126756 11364
rect 125508 6860 125560 6866
rect 125508 6802 125560 6808
rect 126808 6730 126836 60044
rect 126992 60030 127190 60058
rect 127466 60030 127664 60058
rect 127742 60030 127940 60058
rect 126992 46306 127020 60030
rect 127072 57316 127124 57322
rect 127072 57258 127124 57264
rect 126888 46300 126940 46306
rect 126888 46242 126940 46248
rect 126980 46300 127032 46306
rect 126980 46242 127032 46248
rect 126900 6798 126928 46242
rect 127084 46238 127112 57258
rect 127636 51074 127664 60030
rect 127912 55758 127940 60030
rect 128004 57322 128032 60044
rect 128096 60030 128294 60058
rect 127992 57316 128044 57322
rect 127992 57258 128044 57264
rect 127900 55752 127952 55758
rect 127900 55694 127952 55700
rect 128096 51074 128124 60030
rect 128176 57996 128228 58002
rect 128176 57938 128228 57944
rect 128188 57322 128216 57938
rect 128556 57458 128584 60044
rect 128938 60030 129136 60058
rect 128268 57452 128320 57458
rect 128268 57394 128320 57400
rect 128544 57452 128596 57458
rect 128544 57394 128596 57400
rect 128176 57316 128228 57322
rect 128176 57258 128228 57264
rect 128280 56574 128308 57394
rect 128268 56568 128320 56574
rect 128268 56510 128320 56516
rect 128176 55752 128228 55758
rect 128176 55694 128228 55700
rect 127636 51046 127940 51074
rect 127072 46232 127124 46238
rect 127072 46174 127124 46180
rect 127912 17882 127940 51046
rect 128004 51046 128124 51074
rect 127900 17876 127952 17882
rect 127900 17818 127952 17824
rect 128004 17814 128032 51046
rect 128084 46232 128136 46238
rect 128084 46174 128136 46180
rect 127992 17808 128044 17814
rect 127992 17750 128044 17756
rect 128096 11490 128124 46174
rect 128084 11484 128136 11490
rect 128084 11426 128136 11432
rect 126888 6792 126940 6798
rect 126888 6734 126940 6740
rect 126796 6724 126848 6730
rect 126796 6666 126848 6672
rect 128188 6662 128216 55694
rect 129108 55214 129136 60030
rect 129200 57089 129228 60044
rect 129490 60030 129596 60058
rect 129766 60030 129964 60058
rect 129186 57080 129242 57089
rect 129186 57015 129242 57024
rect 129108 55186 129504 55214
rect 128268 46300 128320 46306
rect 128268 46242 128320 46248
rect 128176 6656 128228 6662
rect 128176 6598 128228 6604
rect 128176 6248 128228 6254
rect 128176 6190 128228 6196
rect 125416 6112 125468 6118
rect 125416 6054 125468 6060
rect 124128 6044 124180 6050
rect 124128 5986 124180 5992
rect 126980 4276 127032 4282
rect 126980 4218 127032 4224
rect 124680 3528 124732 3534
rect 124680 3470 124732 3476
rect 123576 3188 123628 3194
rect 123576 3130 123628 3136
rect 124692 480 124720 3470
rect 125876 3188 125928 3194
rect 125876 3130 125928 3136
rect 125888 480 125916 3130
rect 126992 480 127020 4218
rect 128188 480 128216 6190
rect 128280 3126 128308 46242
rect 129476 11558 129504 55186
rect 129464 11552 129516 11558
rect 129464 11494 129516 11500
rect 129568 6526 129596 60030
rect 129648 57452 129700 57458
rect 129648 57394 129700 57400
rect 129660 6594 129688 57394
rect 129832 57316 129884 57322
rect 129832 57258 129884 57264
rect 129844 56778 129872 57258
rect 129936 56953 129964 60030
rect 130028 57322 130056 60044
rect 130120 60030 130318 60058
rect 130686 60030 130884 60058
rect 130016 57316 130068 57322
rect 130016 57258 130068 57264
rect 129922 56944 129978 56953
rect 129922 56879 129978 56888
rect 129740 56772 129792 56778
rect 129740 56714 129792 56720
rect 129832 56772 129884 56778
rect 129832 56714 129884 56720
rect 129752 55962 129780 56714
rect 129832 56568 129884 56574
rect 129832 56510 129884 56516
rect 129740 55956 129792 55962
rect 129740 55898 129792 55904
rect 129844 55842 129872 56510
rect 129752 55814 129872 55842
rect 129752 54262 129780 55814
rect 129740 54256 129792 54262
rect 129740 54198 129792 54204
rect 130120 50386 130148 60030
rect 130752 57452 130804 57458
rect 130752 57394 130804 57400
rect 130384 56772 130436 56778
rect 130384 56714 130436 56720
rect 130108 50380 130160 50386
rect 130108 50322 130160 50328
rect 130396 24138 130424 56714
rect 130384 24132 130436 24138
rect 130384 24074 130436 24080
rect 130764 17746 130792 57394
rect 130752 17740 130804 17746
rect 130752 17682 130804 17688
rect 130856 11626 130884 60030
rect 130948 57458 130976 60044
rect 130936 57452 130988 57458
rect 130936 57394 130988 57400
rect 131120 57452 131172 57458
rect 131120 57394 131172 57400
rect 131028 57316 131080 57322
rect 131028 57258 131080 57264
rect 130936 50380 130988 50386
rect 130936 50322 130988 50328
rect 130844 11620 130896 11626
rect 130844 11562 130896 11568
rect 129648 6588 129700 6594
rect 129648 6530 129700 6536
rect 129556 6520 129608 6526
rect 129556 6462 129608 6468
rect 130948 6458 130976 50322
rect 130936 6452 130988 6458
rect 130936 6394 130988 6400
rect 130568 6180 130620 6186
rect 130568 6122 130620 6128
rect 129372 3732 129424 3738
rect 129372 3674 129424 3680
rect 128268 3120 128320 3126
rect 128268 3062 128320 3068
rect 129384 480 129412 3674
rect 130580 480 130608 6122
rect 131040 3194 131068 57258
rect 131132 54330 131160 57394
rect 131224 56778 131252 60044
rect 131500 57322 131528 60044
rect 131790 60030 131988 60058
rect 131960 57497 131988 60030
rect 131946 57488 132002 57497
rect 132052 57458 132080 60044
rect 132236 60030 132434 60058
rect 132710 60030 132908 60058
rect 132986 60030 133184 60058
rect 131946 57423 132002 57432
rect 132040 57452 132092 57458
rect 132040 57394 132092 57400
rect 131488 57316 131540 57322
rect 131488 57258 131540 57264
rect 132132 57316 132184 57322
rect 132132 57258 132184 57264
rect 131212 56772 131264 56778
rect 131212 56714 131264 56720
rect 131120 54324 131172 54330
rect 131120 54266 131172 54272
rect 132144 11694 132172 57258
rect 132236 12442 132264 60030
rect 132880 58002 132908 60030
rect 132868 57996 132920 58002
rect 132868 57938 132920 57944
rect 133052 57520 133104 57526
rect 132866 57488 132922 57497
rect 132776 57452 132828 57458
rect 133052 57462 133104 57468
rect 132866 57423 132922 57432
rect 132776 57394 132828 57400
rect 132500 57316 132552 57322
rect 132500 57258 132552 57264
rect 132512 56953 132540 57258
rect 132684 57044 132736 57050
rect 132684 56986 132736 56992
rect 132696 56953 132724 56986
rect 132498 56944 132554 56953
rect 132498 56879 132554 56888
rect 132682 56944 132738 56953
rect 132682 56879 132738 56888
rect 132500 56840 132552 56846
rect 132684 56840 132736 56846
rect 132552 56788 132684 56794
rect 132500 56782 132736 56788
rect 132408 56772 132460 56778
rect 132512 56766 132724 56782
rect 132408 56714 132460 56720
rect 132316 54324 132368 54330
rect 132316 54266 132368 54272
rect 132224 12436 132276 12442
rect 132224 12378 132276 12384
rect 132132 11688 132184 11694
rect 132132 11630 132184 11636
rect 132328 6322 132356 54266
rect 132420 6390 132448 56714
rect 132788 54330 132816 57394
rect 132880 57050 132908 57423
rect 133064 57089 133092 57462
rect 133050 57080 133106 57089
rect 132868 57044 132920 57050
rect 133050 57015 133106 57024
rect 132868 56986 132920 56992
rect 133156 55214 133184 60030
rect 133248 57526 133276 60044
rect 133538 60030 133644 60058
rect 133236 57520 133288 57526
rect 133236 57462 133288 57468
rect 133156 55186 133552 55214
rect 132776 54324 132828 54330
rect 132776 54266 132828 54272
rect 132408 6384 132460 6390
rect 132408 6326 132460 6332
rect 132316 6316 132368 6322
rect 132316 6258 132368 6264
rect 133524 6254 133552 55186
rect 133616 17610 133644 60030
rect 133696 57520 133748 57526
rect 133696 57462 133748 57468
rect 133604 17604 133656 17610
rect 133604 17546 133656 17552
rect 133708 12374 133736 57462
rect 133800 57458 133828 60044
rect 134168 57526 134196 60044
rect 134156 57520 134208 57526
rect 134156 57462 134208 57468
rect 134444 57458 134472 60044
rect 133788 57452 133840 57458
rect 133788 57394 133840 57400
rect 134432 57452 134484 57458
rect 134432 57394 134484 57400
rect 133788 56976 133840 56982
rect 133788 56918 133840 56924
rect 133800 56778 133828 56918
rect 134720 56914 134748 60044
rect 135010 60030 135116 60058
rect 134892 57520 134944 57526
rect 134892 57462 134944 57468
rect 134798 57080 134854 57089
rect 134798 57015 134854 57024
rect 134812 56914 134840 57015
rect 133972 56908 134024 56914
rect 133972 56850 134024 56856
rect 134708 56908 134760 56914
rect 134708 56850 134760 56856
rect 134800 56908 134852 56914
rect 134800 56850 134852 56856
rect 133788 56772 133840 56778
rect 133788 56714 133840 56720
rect 133984 54398 134012 56850
rect 133972 54392 134024 54398
rect 133972 54334 134024 54340
rect 133696 12368 133748 12374
rect 133696 12310 133748 12316
rect 134904 12306 134932 57462
rect 134984 57452 135036 57458
rect 134984 57394 135036 57400
rect 134996 17542 135024 57394
rect 134984 17536 135036 17542
rect 134984 17478 135036 17484
rect 134892 12300 134944 12306
rect 134892 12242 134944 12248
rect 135088 12238 135116 60030
rect 135272 50386 135300 60044
rect 135640 57458 135668 60044
rect 135916 57526 135944 60044
rect 136206 60030 136312 60058
rect 135904 57520 135956 57526
rect 135904 57462 135956 57468
rect 135628 57452 135680 57458
rect 135628 57394 135680 57400
rect 135444 56976 135496 56982
rect 135444 56918 135496 56924
rect 135260 50380 135312 50386
rect 135260 50322 135312 50328
rect 135456 45554 135484 56918
rect 135272 45526 135484 45554
rect 135076 12232 135128 12238
rect 135076 12174 135128 12180
rect 134156 8016 134208 8022
rect 134156 7958 134208 7964
rect 133512 6248 133564 6254
rect 133512 6190 133564 6196
rect 132960 4344 133012 4350
rect 132960 4286 133012 4292
rect 131764 3460 131816 3466
rect 131764 3402 131816 3408
rect 131028 3188 131080 3194
rect 131028 3130 131080 3136
rect 131776 480 131804 3402
rect 132972 480 133000 4286
rect 134168 480 134196 7958
rect 135272 480 135300 45526
rect 136284 17474 136312 60030
rect 136468 57526 136496 60044
rect 136364 57520 136416 57526
rect 136364 57462 136416 57468
rect 136456 57520 136508 57526
rect 136456 57462 136508 57468
rect 136272 17468 136324 17474
rect 136272 17410 136324 17416
rect 136376 12170 136404 57462
rect 136744 57458 136772 60044
rect 136548 57452 136600 57458
rect 136548 57394 136600 57400
rect 136732 57452 136784 57458
rect 136732 57394 136784 57400
rect 136456 50380 136508 50386
rect 136456 50322 136508 50328
rect 136364 12164 136416 12170
rect 136364 12106 136416 12112
rect 136468 6914 136496 50322
rect 136376 6886 136496 6914
rect 136376 3330 136404 6886
rect 136456 4412 136508 4418
rect 136456 4354 136508 4360
rect 136364 3324 136416 3330
rect 136364 3266 136416 3272
rect 136468 480 136496 4354
rect 136560 3398 136588 57394
rect 137020 56982 137048 60044
rect 137112 60030 137402 60058
rect 137008 56976 137060 56982
rect 137008 56918 137060 56924
rect 136822 56808 136878 56817
rect 136732 56772 136784 56778
rect 136822 56743 136824 56752
rect 136732 56714 136784 56720
rect 136876 56743 136878 56752
rect 136824 56714 136876 56720
rect 136744 45554 136772 56714
rect 137112 55214 137140 60030
rect 137192 57520 137244 57526
rect 137192 57462 137244 57468
rect 137100 55208 137152 55214
rect 137100 55150 137152 55156
rect 137204 54466 137232 57462
rect 137192 54460 137244 54466
rect 137192 54402 137244 54408
rect 136744 45526 137324 45554
rect 137296 3534 137324 45526
rect 137664 12034 137692 60044
rect 137756 60030 137954 60058
rect 138230 60030 138336 60058
rect 137756 17406 137784 60030
rect 138112 57520 138164 57526
rect 138112 57462 138164 57468
rect 137836 57452 137888 57458
rect 137836 57394 137888 57400
rect 137744 17400 137796 17406
rect 137744 17342 137796 17348
rect 137848 12102 137876 57394
rect 137926 56944 137982 56953
rect 137926 56879 137982 56888
rect 137940 50250 137968 56879
rect 138020 56772 138072 56778
rect 138020 56714 138072 56720
rect 137928 50244 137980 50250
rect 137928 50186 137980 50192
rect 138032 16574 138060 56714
rect 138124 55078 138152 57462
rect 138308 55146 138336 60030
rect 138492 56778 138520 60044
rect 138768 56914 138796 60044
rect 139136 57526 139164 60044
rect 139124 57520 139176 57526
rect 139124 57462 139176 57468
rect 139412 57458 139440 60044
rect 139702 60030 139900 60058
rect 139400 57452 139452 57458
rect 139400 57394 139452 57400
rect 138664 56908 138716 56914
rect 138664 56850 138716 56856
rect 138756 56908 138808 56914
rect 138756 56850 138808 56856
rect 138860 56868 139256 56896
rect 138676 56794 138704 56850
rect 138860 56794 138888 56868
rect 138480 56772 138532 56778
rect 138676 56766 138888 56794
rect 139228 56778 139256 56868
rect 139124 56772 139176 56778
rect 138480 56714 138532 56720
rect 139124 56714 139176 56720
rect 139216 56772 139268 56778
rect 139216 56714 139268 56720
rect 138296 55140 138348 55146
rect 138296 55082 138348 55088
rect 138112 55072 138164 55078
rect 138112 55014 138164 55020
rect 138032 16546 138888 16574
rect 137836 12096 137888 12102
rect 137836 12038 137888 12044
rect 137652 12028 137704 12034
rect 137652 11970 137704 11976
rect 137652 7948 137704 7954
rect 137652 7890 137704 7896
rect 137284 3528 137336 3534
rect 137284 3470 137336 3476
rect 136548 3392 136600 3398
rect 136548 3334 136600 3340
rect 137664 480 137692 7890
rect 138860 480 138888 16546
rect 139136 11966 139164 56714
rect 139872 56506 139900 60030
rect 139964 57526 139992 60044
rect 140240 58546 140268 60044
rect 140424 60030 140530 60058
rect 140228 58540 140280 58546
rect 140228 58482 140280 58488
rect 139952 57520 140004 57526
rect 140424 57497 140452 60030
rect 140688 58540 140740 58546
rect 140688 58482 140740 58488
rect 139952 57462 140004 57468
rect 140410 57488 140466 57497
rect 140410 57423 140466 57432
rect 140596 57452 140648 57458
rect 140596 57394 140648 57400
rect 139860 56500 139912 56506
rect 139860 56442 139912 56448
rect 139124 11960 139176 11966
rect 139124 11902 139176 11908
rect 140608 11898 140636 57394
rect 140596 11892 140648 11898
rect 140596 11834 140648 11840
rect 140700 11830 140728 58482
rect 140780 57520 140832 57526
rect 140780 57462 140832 57468
rect 140792 55010 140820 57462
rect 140780 55004 140832 55010
rect 140780 54946 140832 54952
rect 140884 54942 140912 60044
rect 140964 57996 141016 58002
rect 140964 57938 141016 57944
rect 140976 57458 141004 57938
rect 141160 57526 141188 60044
rect 141148 57520 141200 57526
rect 141148 57462 141200 57468
rect 140964 57452 141016 57458
rect 140964 57394 141016 57400
rect 141436 56982 141464 60044
rect 141726 60030 141832 60058
rect 141332 56976 141384 56982
rect 141332 56918 141384 56924
rect 141424 56976 141476 56982
rect 141424 56918 141476 56924
rect 140872 54936 140924 54942
rect 140872 54878 140924 54884
rect 141344 49162 141372 56918
rect 141332 49156 141384 49162
rect 141332 49098 141384 49104
rect 140688 11824 140740 11830
rect 140688 11766 140740 11772
rect 141240 7880 141292 7886
rect 141240 7822 141292 7828
rect 140044 3528 140096 3534
rect 140044 3470 140096 3476
rect 140056 480 140084 3470
rect 141252 480 141280 7822
rect 141804 7070 141832 60030
rect 141896 60030 142002 60058
rect 141896 17270 141924 60030
rect 142264 57526 142292 60044
rect 142632 57594 142660 60044
rect 142816 60030 142922 60058
rect 143198 60030 143304 60058
rect 142528 57588 142580 57594
rect 142528 57530 142580 57536
rect 142620 57588 142672 57594
rect 142620 57530 142672 57536
rect 141976 57520 142028 57526
rect 141976 57462 142028 57468
rect 142252 57520 142304 57526
rect 142252 57462 142304 57468
rect 141884 17264 141936 17270
rect 141884 17206 141936 17212
rect 141988 11762 142016 57462
rect 142066 57216 142122 57225
rect 142066 57151 142122 57160
rect 142250 57216 142306 57225
rect 142250 57151 142306 57160
rect 142080 56914 142108 57151
rect 142264 57050 142292 57151
rect 142160 57044 142212 57050
rect 142160 56986 142212 56992
rect 142252 57044 142304 57050
rect 142252 56986 142304 56992
rect 142172 56930 142200 56986
rect 142068 56908 142120 56914
rect 142172 56902 142292 56930
rect 142540 56914 142568 57530
rect 142068 56850 142120 56856
rect 142068 56772 142120 56778
rect 142068 56714 142120 56720
rect 142080 56438 142108 56714
rect 142264 56710 142292 56902
rect 142528 56908 142580 56914
rect 142528 56850 142580 56856
rect 142252 56704 142304 56710
rect 142252 56646 142304 56652
rect 142160 56636 142212 56642
rect 142160 56578 142212 56584
rect 142172 56522 142200 56578
rect 142172 56494 142752 56522
rect 142068 56432 142120 56438
rect 142068 56374 142120 56380
rect 142620 56432 142672 56438
rect 142620 56374 142672 56380
rect 141976 11756 142028 11762
rect 141976 11698 142028 11704
rect 141792 7064 141844 7070
rect 141792 7006 141844 7012
rect 142632 6914 142660 56374
rect 142724 45554 142752 56494
rect 142816 52290 142844 60030
rect 143172 58064 143224 58070
rect 143172 58006 143224 58012
rect 143184 57866 143212 58006
rect 143276 58002 143304 60030
rect 143368 60030 143474 60058
rect 143264 57996 143316 58002
rect 143264 57938 143316 57944
rect 143172 57860 143224 57866
rect 143172 57802 143224 57808
rect 143264 57860 143316 57866
rect 143264 57802 143316 57808
rect 143276 57186 143304 57802
rect 143264 57180 143316 57186
rect 143264 57122 143316 57128
rect 142894 57080 142950 57089
rect 142894 57015 142950 57024
rect 142908 52766 142936 57015
rect 142896 52760 142948 52766
rect 142896 52702 142948 52708
rect 142804 52284 142856 52290
rect 142804 52226 142856 52232
rect 142724 45526 142844 45554
rect 142448 6886 142660 6914
rect 142448 480 142476 6886
rect 142816 4418 142844 45526
rect 143368 7206 143396 60030
rect 143448 57996 143500 58002
rect 143448 57938 143500 57944
rect 143460 57746 143488 57938
rect 143460 57718 143580 57746
rect 143552 57594 143580 57718
rect 143448 57588 143500 57594
rect 143448 57530 143500 57536
rect 143540 57588 143592 57594
rect 143540 57530 143592 57536
rect 143356 7200 143408 7206
rect 143356 7142 143408 7148
rect 143460 7138 143488 57530
rect 143540 57180 143592 57186
rect 143540 57122 143592 57128
rect 143552 52154 143580 57122
rect 143736 52222 143764 60044
rect 144026 60030 144316 60058
rect 144394 60030 144592 60058
rect 143906 57624 143962 57633
rect 143906 57559 143962 57568
rect 143724 52216 143776 52222
rect 143724 52158 143776 52164
rect 143540 52148 143592 52154
rect 143540 52090 143592 52096
rect 143920 51678 143948 57559
rect 144288 57526 144316 60030
rect 144184 57520 144236 57526
rect 144184 57462 144236 57468
rect 144276 57520 144328 57526
rect 144276 57462 144328 57468
rect 143908 51672 143960 51678
rect 143908 51614 143960 51620
rect 144196 17338 144224 57462
rect 144564 55214 144592 60030
rect 144656 57186 144684 60044
rect 144946 60030 145144 60058
rect 144828 57520 144880 57526
rect 144828 57462 144880 57468
rect 144840 57186 144868 57462
rect 144644 57180 144696 57186
rect 144644 57122 144696 57128
rect 144828 57180 144880 57186
rect 144828 57122 144880 57128
rect 145116 56914 145144 60030
rect 145208 57526 145236 60044
rect 145196 57520 145248 57526
rect 145196 57462 145248 57468
rect 144920 56908 144972 56914
rect 144920 56850 144972 56856
rect 145104 56908 145156 56914
rect 145104 56850 145156 56856
rect 144564 55186 144868 55214
rect 144184 17332 144236 17338
rect 144184 17274 144236 17280
rect 144736 7812 144788 7818
rect 144736 7754 144788 7760
rect 143448 7132 143500 7138
rect 143448 7074 143500 7080
rect 143540 4480 143592 4486
rect 143540 4422 143592 4428
rect 142804 4412 142856 4418
rect 142804 4354 142856 4360
rect 143552 480 143580 4422
rect 144748 480 144776 7754
rect 144840 7274 144868 55186
rect 144932 16574 144960 56850
rect 145484 52086 145512 60044
rect 145774 60030 146064 60058
rect 146142 60030 146248 60058
rect 146036 57610 146064 60030
rect 146220 57746 146248 60030
rect 146220 57718 146340 57746
rect 146036 57582 146248 57610
rect 146116 57520 146168 57526
rect 146116 57462 146168 57468
rect 145472 52080 145524 52086
rect 145472 52022 145524 52028
rect 144932 16546 145972 16574
rect 144828 7268 144880 7274
rect 144828 7210 144880 7216
rect 145944 480 145972 16546
rect 146128 7342 146156 57462
rect 146116 7336 146168 7342
rect 146116 7278 146168 7284
rect 146220 4010 146248 57582
rect 146312 57361 146340 57718
rect 146298 57352 146354 57361
rect 146298 57287 146354 57296
rect 146404 57186 146432 60044
rect 146680 57594 146708 60044
rect 146970 60030 147168 60058
rect 147246 60030 147444 60058
rect 147522 60030 147628 60058
rect 146668 57588 146720 57594
rect 146668 57530 146720 57536
rect 146300 57180 146352 57186
rect 146300 57122 146352 57128
rect 146392 57180 146444 57186
rect 146392 57122 146444 57128
rect 146312 57066 146340 57122
rect 146312 57038 146708 57066
rect 146680 56846 146708 57038
rect 146944 56976 146996 56982
rect 146944 56918 146996 56924
rect 146576 56840 146628 56846
rect 146576 56782 146628 56788
rect 146668 56840 146720 56846
rect 146668 56782 146720 56788
rect 146588 45554 146616 56782
rect 146956 56778 146984 56918
rect 146852 56772 146904 56778
rect 146852 56714 146904 56720
rect 146944 56772 146996 56778
rect 146944 56714 146996 56720
rect 146864 55214 146892 56714
rect 147140 55214 147168 60030
rect 147312 57520 147364 57526
rect 147312 57462 147364 57468
rect 147324 56982 147352 57462
rect 147312 56976 147364 56982
rect 147312 56918 147364 56924
rect 146864 55186 147076 55214
rect 147140 55186 147352 55214
rect 146588 45526 146984 45554
rect 146956 4486 146984 45526
rect 147048 16574 147076 55186
rect 147048 16546 147260 16574
rect 147232 4622 147260 16546
rect 147324 7410 147352 55186
rect 147312 7404 147364 7410
rect 147312 7346 147364 7352
rect 147128 4616 147180 4622
rect 147128 4558 147180 4564
rect 147220 4616 147272 4622
rect 147220 4558 147272 4564
rect 146944 4480 146996 4486
rect 146944 4422 146996 4428
rect 146208 4004 146260 4010
rect 146208 3946 146260 3952
rect 147140 480 147168 4558
rect 147416 3874 147444 60030
rect 147496 57588 147548 57594
rect 147496 57530 147548 57536
rect 147508 3942 147536 57530
rect 147496 3936 147548 3942
rect 147496 3878 147548 3884
rect 147404 3868 147456 3874
rect 147404 3810 147456 3816
rect 147600 3806 147628 60030
rect 147680 57588 147732 57594
rect 147680 57530 147732 57536
rect 147692 57254 147720 57530
rect 147680 57248 147732 57254
rect 147680 57190 147732 57196
rect 147876 56710 147904 60044
rect 148048 57520 148100 57526
rect 148048 57462 148100 57468
rect 147956 57248 148008 57254
rect 147956 57190 148008 57196
rect 147772 56704 147824 56710
rect 147772 56646 147824 56652
rect 147864 56704 147916 56710
rect 147864 56646 147916 56652
rect 147784 56522 147812 56646
rect 147968 56522 147996 57190
rect 147784 56494 147996 56522
rect 148060 51074 148088 57462
rect 148152 52018 148180 60044
rect 148442 60030 148640 60058
rect 148718 60030 148916 60058
rect 148324 57860 148376 57866
rect 148324 57802 148376 57808
rect 148140 52012 148192 52018
rect 148140 51954 148192 51960
rect 147692 51046 148088 51074
rect 147692 50318 147720 51046
rect 147680 50312 147732 50318
rect 147680 50254 147732 50260
rect 148232 7744 148284 7750
rect 148232 7686 148284 7692
rect 147588 3800 147640 3806
rect 147588 3742 147640 3748
rect 148244 1578 148272 7686
rect 148336 3466 148364 57802
rect 148612 3738 148640 60030
rect 148784 56704 148836 56710
rect 148784 56646 148836 56652
rect 148796 7478 148824 56646
rect 148888 7546 148916 60030
rect 148980 57526 149008 60044
rect 149256 57866 149284 60044
rect 149428 58064 149480 58070
rect 149428 58006 149480 58012
rect 149244 57860 149296 57866
rect 149244 57802 149296 57808
rect 148968 57520 149020 57526
rect 148968 57462 149020 57468
rect 149440 16574 149468 58006
rect 149624 56710 149652 60044
rect 149612 56704 149664 56710
rect 149612 56646 149664 56652
rect 149900 51950 149928 60044
rect 150190 60030 150388 60058
rect 150256 57520 150308 57526
rect 150256 57462 150308 57468
rect 150268 56982 150296 57462
rect 150256 56976 150308 56982
rect 150256 56918 150308 56924
rect 150256 56704 150308 56710
rect 150256 56646 150308 56652
rect 149888 51944 149940 51950
rect 149888 51886 149940 51892
rect 149440 16546 149560 16574
rect 148876 7540 148928 7546
rect 148876 7482 148928 7488
rect 148784 7472 148836 7478
rect 148784 7414 148836 7420
rect 148600 3732 148652 3738
rect 148600 3674 148652 3680
rect 148324 3460 148376 3466
rect 148324 3402 148376 3408
rect 148244 1550 148364 1578
rect 148336 480 148364 1550
rect 149532 480 149560 16546
rect 150268 8294 150296 56646
rect 150256 8288 150308 8294
rect 150256 8230 150308 8236
rect 150360 3670 150388 60030
rect 150452 56982 150480 60044
rect 150742 60030 151032 60058
rect 150440 56976 150492 56982
rect 150440 56918 150492 56924
rect 151004 51074 151032 60030
rect 151096 56710 151124 60044
rect 151386 60030 151492 60058
rect 151662 60030 151768 60058
rect 151084 56704 151136 56710
rect 151084 56646 151136 56652
rect 151004 51046 151400 51074
rect 151372 12646 151400 51046
rect 151360 12640 151412 12646
rect 151360 12582 151412 12588
rect 151464 8158 151492 60030
rect 151544 56976 151596 56982
rect 151544 56918 151596 56924
rect 151556 8226 151584 56918
rect 151636 56704 151688 56710
rect 151636 56646 151688 56652
rect 151544 8220 151596 8226
rect 151544 8162 151596 8168
rect 151452 8152 151504 8158
rect 151452 8094 151504 8100
rect 151648 6186 151676 56646
rect 151636 6180 151688 6186
rect 151636 6122 151688 6128
rect 151740 5817 151768 60030
rect 151820 57248 151872 57254
rect 151820 57190 151872 57196
rect 151832 49366 151860 57190
rect 151924 56982 151952 60044
rect 152214 60030 152412 60058
rect 152490 60030 152780 60058
rect 152188 57588 152240 57594
rect 152188 57530 152240 57536
rect 151912 56976 151964 56982
rect 151912 56918 151964 56924
rect 151820 49360 151872 49366
rect 151820 49302 151872 49308
rect 151820 7676 151872 7682
rect 151820 7618 151872 7624
rect 151726 5808 151782 5817
rect 151726 5743 151782 5752
rect 150348 3664 150400 3670
rect 150348 3606 150400 3612
rect 150624 3460 150676 3466
rect 150624 3402 150676 3408
rect 150636 480 150664 3402
rect 151832 480 151860 7618
rect 152200 6914 152228 57530
rect 152384 55758 152412 60030
rect 152464 57588 152516 57594
rect 152464 57530 152516 57536
rect 152476 57186 152504 57530
rect 152464 57180 152516 57186
rect 152464 57122 152516 57128
rect 152372 55752 152424 55758
rect 152372 55694 152424 55700
rect 152752 12714 152780 60030
rect 152844 56710 152872 60044
rect 152936 60030 153134 60058
rect 152832 56704 152884 56710
rect 152832 56646 152884 56652
rect 152832 55752 152884 55758
rect 152832 55694 152884 55700
rect 152740 12708 152792 12714
rect 152740 12650 152792 12656
rect 152844 8090 152872 55694
rect 152832 8084 152884 8090
rect 152832 8026 152884 8032
rect 152936 8022 152964 60030
rect 153396 56982 153424 60044
rect 153672 57118 153700 60044
rect 153660 57112 153712 57118
rect 153660 57054 153712 57060
rect 153108 56976 153160 56982
rect 153108 56918 153160 56924
rect 153384 56976 153436 56982
rect 153384 56918 153436 56924
rect 153016 56704 153068 56710
rect 153016 56646 153068 56652
rect 152924 8016 152976 8022
rect 152924 7958 152976 7964
rect 152200 6886 152964 6914
rect 152936 3482 152964 6886
rect 153028 3602 153056 56646
rect 153120 3602 153148 56918
rect 153948 56710 153976 60044
rect 154238 60030 154344 60058
rect 154212 56976 154264 56982
rect 154212 56918 154264 56924
rect 153936 56704 153988 56710
rect 153936 56646 153988 56652
rect 154224 12782 154252 56918
rect 154316 12850 154344 60030
rect 154488 57112 154540 57118
rect 154488 57054 154540 57060
rect 154396 56704 154448 56710
rect 154396 56646 154448 56652
rect 154304 12844 154356 12850
rect 154304 12786 154356 12792
rect 154212 12776 154264 12782
rect 154212 12718 154264 12724
rect 154408 7954 154436 56646
rect 154396 7948 154448 7954
rect 154396 7890 154448 7896
rect 154212 4548 154264 4554
rect 154212 4490 154264 4496
rect 153016 3596 153068 3602
rect 153016 3538 153068 3544
rect 153108 3596 153160 3602
rect 153108 3538 153160 3544
rect 152936 3454 153056 3482
rect 153028 480 153056 3454
rect 154224 480 154252 4490
rect 154500 3466 154528 57054
rect 154592 56982 154620 60044
rect 154580 56976 154632 56982
rect 154580 56918 154632 56924
rect 154868 56710 154896 60044
rect 155158 60030 155356 60058
rect 154856 56704 154908 56710
rect 154856 56646 154908 56652
rect 155328 51074 155356 60030
rect 155420 57254 155448 60044
rect 155408 57248 155460 57254
rect 155408 57190 155460 57196
rect 155328 51046 155632 51074
rect 155604 12918 155632 51046
rect 155592 12912 155644 12918
rect 155592 12854 155644 12860
rect 155696 7818 155724 60044
rect 155972 56982 156000 60044
rect 156144 57180 156196 57186
rect 156144 57122 156196 57128
rect 155868 56976 155920 56982
rect 155868 56918 155920 56924
rect 155960 56976 156012 56982
rect 155960 56918 156012 56924
rect 155776 56704 155828 56710
rect 155776 56646 155828 56652
rect 155788 7886 155816 56646
rect 155776 7880 155828 7886
rect 155776 7822 155828 7828
rect 155684 7812 155736 7818
rect 155684 7754 155736 7760
rect 155408 7608 155460 7614
rect 155408 7550 155460 7556
rect 154488 3460 154540 3466
rect 154488 3402 154540 3408
rect 155420 480 155448 7550
rect 155880 5953 155908 56918
rect 156052 56840 156104 56846
rect 156052 56782 156104 56788
rect 156064 49094 156092 56782
rect 156156 52698 156184 57122
rect 156340 57118 156368 60044
rect 156630 60030 156828 60058
rect 156906 60030 157012 60058
rect 157182 60030 157288 60058
rect 157458 60030 157656 60058
rect 157734 60030 158024 60058
rect 156800 58018 156828 60030
rect 156800 57990 156920 58018
rect 156892 57866 156920 57990
rect 156788 57860 156840 57866
rect 156788 57802 156840 57808
rect 156880 57860 156932 57866
rect 156880 57802 156932 57808
rect 156328 57112 156380 57118
rect 156328 57054 156380 57060
rect 156800 56710 156828 57802
rect 156788 56704 156840 56710
rect 156788 56646 156840 56652
rect 156696 56636 156748 56642
rect 156696 56578 156748 56584
rect 156144 52692 156196 52698
rect 156144 52634 156196 52640
rect 156708 49230 156736 56578
rect 156696 49224 156748 49230
rect 156696 49166 156748 49172
rect 156052 49088 156104 49094
rect 156052 49030 156104 49036
rect 156984 13054 157012 60030
rect 157156 57860 157208 57866
rect 157156 57802 157208 57808
rect 157064 56976 157116 56982
rect 157064 56918 157116 56924
rect 156972 13048 157024 13054
rect 156972 12990 157024 12996
rect 157076 12986 157104 56918
rect 157064 12980 157116 12986
rect 157064 12922 157116 12928
rect 157168 7750 157196 57802
rect 157156 7744 157208 7750
rect 157156 7686 157208 7692
rect 157260 6089 157288 60030
rect 157628 54874 157656 60030
rect 157996 55570 158024 60030
rect 158088 56642 158116 60044
rect 158378 60030 158484 60058
rect 158076 56636 158128 56642
rect 158076 56578 158128 56584
rect 157996 55542 158392 55570
rect 158260 55344 158312 55350
rect 158260 55286 158312 55292
rect 157616 54868 157668 54874
rect 157616 54810 157668 54816
rect 158272 13734 158300 55286
rect 158364 13802 158392 55542
rect 158352 13796 158404 13802
rect 158352 13738 158404 13744
rect 158260 13728 158312 13734
rect 158260 13670 158312 13676
rect 158456 7614 158484 60030
rect 158548 60030 158654 60058
rect 158548 55350 158576 60030
rect 158916 56642 158944 60044
rect 159192 57866 159220 60044
rect 159482 60030 159772 60058
rect 159180 57860 159232 57866
rect 159180 57802 159232 57808
rect 158628 56636 158680 56642
rect 158628 56578 158680 56584
rect 158904 56636 158956 56642
rect 158904 56578 158956 56584
rect 158536 55344 158588 55350
rect 158536 55286 158588 55292
rect 158536 54868 158588 54874
rect 158536 54810 158588 54816
rect 158548 7682 158576 54810
rect 158536 7676 158588 7682
rect 158536 7618 158588 7624
rect 158444 7608 158496 7614
rect 158444 7550 158496 7556
rect 158640 6905 158668 56578
rect 159744 51074 159772 60030
rect 159836 57934 159864 60044
rect 159824 57928 159876 57934
rect 159824 57870 159876 57876
rect 160008 56636 160060 56642
rect 160008 56578 160060 56584
rect 159744 51046 159956 51074
rect 159928 13666 159956 51046
rect 159916 13660 159968 13666
rect 159916 13602 159968 13608
rect 158904 9376 158956 9382
rect 158904 9318 158956 9324
rect 158626 6896 158682 6905
rect 158626 6831 158682 6840
rect 157246 6080 157302 6089
rect 157246 6015 157302 6024
rect 155866 5944 155922 5953
rect 155866 5879 155922 5888
rect 157800 4684 157852 4690
rect 157800 4626 157852 4632
rect 156604 4140 156656 4146
rect 156604 4082 156656 4088
rect 156616 480 156644 4082
rect 157812 480 157840 4626
rect 158916 480 158944 9318
rect 160020 2174 160048 56578
rect 160112 54874 160140 60044
rect 160402 60030 160600 60058
rect 160678 60030 160876 60058
rect 160466 57488 160522 57497
rect 160466 57423 160522 57432
rect 160100 54868 160152 54874
rect 160100 54810 160152 54816
rect 160192 52692 160244 52698
rect 160192 52634 160244 52640
rect 160204 6914 160232 52634
rect 160480 51074 160508 57423
rect 160572 55434 160600 60030
rect 160848 55570 160876 60030
rect 160940 56642 160968 60044
rect 160928 56636 160980 56642
rect 160928 56578 160980 56584
rect 160848 55542 161152 55570
rect 160572 55406 161060 55434
rect 160480 51046 160784 51074
rect 160756 18766 160784 51046
rect 160744 18760 160796 18766
rect 160744 18702 160796 18708
rect 161032 13598 161060 55406
rect 161020 13592 161072 13598
rect 161020 13534 161072 13540
rect 160204 6886 161060 6914
rect 160100 4072 160152 4078
rect 160100 4014 160152 4020
rect 160008 2168 160060 2174
rect 160008 2110 160060 2116
rect 160112 480 160140 4014
rect 161032 3482 161060 6886
rect 161124 3913 161152 55542
rect 161216 13530 161244 60044
rect 161584 57050 161612 60044
rect 161572 57044 161624 57050
rect 161572 56986 161624 56992
rect 161388 56636 161440 56642
rect 161388 56578 161440 56584
rect 161400 53786 161428 56578
rect 161860 54806 161888 60044
rect 162032 57792 162084 57798
rect 162032 57734 162084 57740
rect 162044 57118 162072 57734
rect 162032 57112 162084 57118
rect 162032 57054 162084 57060
rect 162136 56642 162164 60044
rect 162426 60030 162532 60058
rect 162216 58132 162268 58138
rect 162216 58074 162268 58080
rect 162228 57798 162256 58074
rect 162216 57792 162268 57798
rect 162216 57734 162268 57740
rect 162124 56636 162176 56642
rect 162124 56578 162176 56584
rect 161848 54800 161900 54806
rect 161848 54742 161900 54748
rect 161388 53780 161440 53786
rect 161388 53722 161440 53728
rect 162504 16574 162532 60030
rect 162596 60030 162702 60058
rect 162596 53718 162624 60030
rect 162768 56976 162820 56982
rect 162768 56918 162820 56924
rect 162780 56642 162808 56918
rect 162964 56778 162992 60044
rect 163332 56982 163360 60044
rect 163320 56976 163372 56982
rect 163320 56918 163372 56924
rect 162952 56772 163004 56778
rect 162952 56714 163004 56720
rect 162676 56636 162728 56642
rect 162676 56578 162728 56584
rect 162768 56636 162820 56642
rect 162768 56578 162820 56584
rect 162584 53712 162636 53718
rect 162584 53654 162636 53660
rect 162504 16546 162624 16574
rect 161204 13524 161256 13530
rect 161204 13466 161256 13472
rect 162492 4752 162544 4758
rect 162492 4694 162544 4700
rect 161110 3904 161166 3913
rect 161110 3839 161166 3848
rect 161032 3454 161336 3482
rect 161308 480 161336 3454
rect 162504 480 162532 4694
rect 162596 3777 162624 16546
rect 162688 13462 162716 56578
rect 163608 55758 163636 60044
rect 163898 60030 164004 60058
rect 163872 56636 163924 56642
rect 163872 56578 163924 56584
rect 163596 55752 163648 55758
rect 163596 55694 163648 55700
rect 162676 13456 162728 13462
rect 162676 13398 162728 13404
rect 163688 9308 163740 9314
rect 163688 9250 163740 9256
rect 162582 3768 162638 3777
rect 162582 3703 162638 3712
rect 163700 480 163728 9250
rect 163884 3641 163912 56578
rect 163976 13326 164004 60030
rect 164056 56772 164108 56778
rect 164056 56714 164108 56720
rect 164068 13394 164096 56714
rect 164160 56642 164188 60044
rect 164148 56636 164200 56642
rect 164148 56578 164200 56584
rect 164436 53650 164464 60044
rect 164516 57792 164568 57798
rect 164516 57734 164568 57740
rect 164424 53644 164476 53650
rect 164424 53586 164476 53592
rect 164528 51074 164556 57734
rect 164712 56642 164740 60044
rect 165094 60030 165292 60058
rect 164608 56636 164660 56642
rect 164608 56578 164660 56584
rect 164700 56636 164752 56642
rect 164700 56578 164752 56584
rect 164620 56522 164648 56578
rect 164620 56494 164740 56522
rect 164712 51074 164740 56494
rect 164528 51046 164648 51074
rect 164712 51046 164924 51074
rect 164620 16574 164648 51046
rect 164896 18834 164924 51046
rect 164884 18828 164936 18834
rect 164884 18770 164936 18776
rect 164620 16546 164924 16574
rect 164056 13388 164108 13394
rect 164056 13330 164108 13336
rect 163964 13320 164016 13326
rect 163964 13262 164016 13268
rect 163870 3632 163926 3641
rect 163870 3567 163926 3576
rect 164896 480 164924 16546
rect 165264 6769 165292 60030
rect 165356 53514 165384 60044
rect 165632 56778 165660 60044
rect 165908 57934 165936 60044
rect 165804 57928 165856 57934
rect 165804 57870 165856 57876
rect 165896 57928 165948 57934
rect 165896 57870 165948 57876
rect 165816 57780 165844 57870
rect 165896 57792 165948 57798
rect 165816 57752 165896 57780
rect 165896 57734 165948 57740
rect 165620 56772 165672 56778
rect 165620 56714 165672 56720
rect 165436 56636 165488 56642
rect 165436 56578 165488 56584
rect 165344 53508 165396 53514
rect 165344 53450 165396 53456
rect 165448 13258 165476 56578
rect 166184 54738 166212 60044
rect 166448 57248 166500 57254
rect 166448 57190 166500 57196
rect 166354 57080 166410 57089
rect 166354 57015 166356 57024
rect 166408 57015 166410 57024
rect 166356 56986 166408 56992
rect 166460 56574 166488 57190
rect 166552 56642 166580 60044
rect 166644 60030 166842 60058
rect 166540 56636 166592 56642
rect 166540 56578 166592 56584
rect 166448 56568 166500 56574
rect 166448 56510 166500 56516
rect 166172 54732 166224 54738
rect 166172 54674 166224 54680
rect 165436 13252 165488 13258
rect 165436 13194 165488 13200
rect 165250 6760 165306 6769
rect 165250 6695 165306 6704
rect 166644 6497 166672 60030
rect 166816 57860 166868 57866
rect 166816 57802 166868 57808
rect 167000 57860 167052 57866
rect 167000 57802 167052 57808
rect 166828 57254 166856 57802
rect 166908 57792 166960 57798
rect 166908 57734 166960 57740
rect 166816 57248 166868 57254
rect 166816 57190 166868 57196
rect 166920 57050 166948 57734
rect 166908 57044 166960 57050
rect 166908 56986 166960 56992
rect 166816 56976 166868 56982
rect 166816 56918 166868 56924
rect 166828 56778 166856 56918
rect 166724 56772 166776 56778
rect 166724 56714 166776 56720
rect 166816 56772 166868 56778
rect 166816 56714 166868 56720
rect 166736 13190 166764 56714
rect 166816 56636 166868 56642
rect 166816 56578 166868 56584
rect 166724 13184 166776 13190
rect 166724 13126 166776 13132
rect 166828 13122 166856 56578
rect 167012 54670 167040 57802
rect 167104 57798 167132 60044
rect 167092 57792 167144 57798
rect 167092 57734 167144 57740
rect 167184 56976 167236 56982
rect 167184 56918 167236 56924
rect 167196 56778 167224 56918
rect 167184 56772 167236 56778
rect 167184 56714 167236 56720
rect 167380 55826 167408 60044
rect 167670 60030 167868 60058
rect 167946 60030 168236 60058
rect 167368 55820 167420 55826
rect 167368 55762 167420 55768
rect 167840 55214 167868 60030
rect 168104 57792 168156 57798
rect 168104 57734 168156 57740
rect 167840 55186 168052 55214
rect 167000 54664 167052 54670
rect 167000 54606 167052 54612
rect 166816 13116 166868 13122
rect 166816 13058 166868 13064
rect 167184 9240 167236 9246
rect 167184 9182 167236 9188
rect 166630 6488 166686 6497
rect 166630 6423 166686 6432
rect 166080 5500 166132 5506
rect 166080 5442 166132 5448
rect 166092 480 166120 5442
rect 167196 480 167224 9182
rect 168024 6361 168052 55186
rect 168116 8362 168144 57734
rect 168208 8430 168236 60030
rect 168300 57866 168328 60044
rect 168576 57934 168604 60044
rect 168564 57928 168616 57934
rect 168564 57870 168616 57876
rect 168852 57866 168880 60044
rect 168288 57860 168340 57866
rect 168288 57802 168340 57808
rect 168840 57860 168892 57866
rect 168840 57802 168892 57808
rect 168564 57112 168616 57118
rect 168656 57112 168708 57118
rect 168564 57054 168616 57060
rect 168654 57080 168656 57089
rect 168708 57080 168710 57089
rect 168380 56772 168432 56778
rect 168380 56714 168432 56720
rect 168392 51882 168420 56714
rect 168576 55214 168604 57054
rect 168654 57015 168710 57024
rect 169128 56778 169156 60044
rect 169404 57798 169432 60044
rect 169496 60030 169694 60058
rect 169772 60030 170062 60058
rect 169392 57792 169444 57798
rect 169392 57734 169444 57740
rect 169116 56772 169168 56778
rect 169116 56714 169168 56720
rect 168576 55186 168880 55214
rect 168380 51876 168432 51882
rect 168380 51818 168432 51824
rect 168196 8424 168248 8430
rect 168196 8366 168248 8372
rect 168104 8356 168156 8362
rect 168104 8298 168156 8304
rect 168852 6914 168880 55186
rect 169496 8566 169524 60030
rect 169576 57860 169628 57866
rect 169576 57802 169628 57808
rect 169484 8560 169536 8566
rect 169484 8502 169536 8508
rect 169588 8498 169616 57802
rect 169668 57792 169720 57798
rect 169668 57734 169720 57740
rect 169576 8492 169628 8498
rect 169576 8434 169628 8440
rect 168392 6886 168880 6914
rect 168010 6352 168066 6361
rect 168010 6287 168066 6296
rect 168392 480 168420 6886
rect 169576 5432 169628 5438
rect 169576 5374 169628 5380
rect 169588 480 169616 5374
rect 169680 3505 169708 57734
rect 169772 50998 169800 60030
rect 169852 57792 169904 57798
rect 169852 57734 169904 57740
rect 169760 50992 169812 50998
rect 169760 50934 169812 50940
rect 169864 50930 169892 57734
rect 170324 56778 170352 60044
rect 170614 60030 170812 60058
rect 170312 56772 170364 56778
rect 170312 56714 170364 56720
rect 170404 56704 170456 56710
rect 170404 56646 170456 56652
rect 169852 50924 169904 50930
rect 169852 50866 169904 50872
rect 170416 18698 170444 56646
rect 170784 55214 170812 60030
rect 170876 57798 170904 60044
rect 170864 57792 170916 57798
rect 170864 57734 170916 57740
rect 171152 57730 171180 60044
rect 171048 57724 171100 57730
rect 171048 57666 171100 57672
rect 171140 57724 171192 57730
rect 171140 57666 171192 57672
rect 171060 57633 171088 57666
rect 171046 57624 171102 57633
rect 171046 57559 171102 57568
rect 171428 56778 171456 60044
rect 171520 60030 171810 60058
rect 172086 60030 172192 60058
rect 171048 56772 171100 56778
rect 171048 56714 171100 56720
rect 171416 56772 171468 56778
rect 171416 56714 171468 56720
rect 170784 55186 170996 55214
rect 170404 18692 170456 18698
rect 170404 18634 170456 18640
rect 170772 9172 170824 9178
rect 170772 9114 170824 9120
rect 169666 3496 169722 3505
rect 169666 3431 169722 3440
rect 170784 480 170812 9114
rect 170968 8634 170996 55186
rect 170956 8628 171008 8634
rect 170956 8570 171008 8576
rect 171060 4214 171088 56714
rect 171520 53446 171548 60030
rect 172164 58138 172192 60030
rect 172256 60030 172362 60058
rect 172152 58132 172204 58138
rect 172152 58074 172204 58080
rect 172152 57724 172204 57730
rect 172152 57666 172204 57672
rect 171598 57624 171654 57633
rect 171598 57559 171654 57568
rect 171508 53440 171560 53446
rect 171508 53382 171560 53388
rect 171612 16574 171640 57559
rect 171612 16546 172008 16574
rect 171048 4208 171100 4214
rect 171048 4150 171100 4156
rect 171980 480 172008 16546
rect 172164 4282 172192 57666
rect 172256 8770 172284 60030
rect 172336 56772 172388 56778
rect 172336 56714 172388 56720
rect 172244 8764 172296 8770
rect 172244 8706 172296 8712
rect 172348 8702 172376 56714
rect 172624 50862 172652 60044
rect 172900 57730 172928 60044
rect 173190 60030 173480 60058
rect 172888 57724 172940 57730
rect 172888 57666 172940 57672
rect 172704 57656 172756 57662
rect 172704 57598 172756 57604
rect 172796 57656 172848 57662
rect 172796 57598 172848 57604
rect 172716 56846 172744 57598
rect 172704 56840 172756 56846
rect 172704 56782 172756 56788
rect 172808 51066 172836 57598
rect 173452 55214 173480 60030
rect 173544 57662 173572 60044
rect 173716 57860 173768 57866
rect 173716 57802 173768 57808
rect 173624 57724 173676 57730
rect 173624 57666 173676 57672
rect 173532 57656 173584 57662
rect 173532 57598 173584 57604
rect 173636 56556 173664 57666
rect 173728 56710 173756 57802
rect 173820 57610 173848 60044
rect 174096 57730 174124 60044
rect 174280 60030 174386 60058
rect 174176 57792 174228 57798
rect 174176 57734 174228 57740
rect 174084 57724 174136 57730
rect 174084 57666 174136 57672
rect 174188 57610 174216 57734
rect 173820 57582 174216 57610
rect 173716 56704 173768 56710
rect 173716 56646 173768 56652
rect 173636 56528 173848 56556
rect 173452 55186 173756 55214
rect 172796 51060 172848 51066
rect 172796 51002 172848 51008
rect 172612 50856 172664 50862
rect 172612 50798 172664 50804
rect 173728 8838 173756 55186
rect 173716 8832 173768 8838
rect 173716 8774 173768 8780
rect 172336 8696 172388 8702
rect 172336 8638 172388 8644
rect 173164 5364 173216 5370
rect 173164 5306 173216 5312
rect 172152 4276 172204 4282
rect 172152 4218 172204 4224
rect 173176 480 173204 5306
rect 173820 4350 173848 56528
rect 174280 50794 174308 60030
rect 174648 57662 174676 60044
rect 174938 60030 175136 60058
rect 175004 57724 175056 57730
rect 175004 57666 175056 57672
rect 174636 57656 174688 57662
rect 174636 57598 174688 57604
rect 174912 56840 174964 56846
rect 174912 56782 174964 56788
rect 174924 56574 174952 56782
rect 174912 56568 174964 56574
rect 174912 56510 174964 56516
rect 174268 50788 174320 50794
rect 174268 50730 174320 50736
rect 174268 9104 174320 9110
rect 174268 9046 174320 9052
rect 173808 4344 173860 4350
rect 173808 4286 173860 4292
rect 174280 480 174308 9046
rect 175016 8906 175044 57666
rect 175108 9654 175136 60030
rect 175188 57656 175240 57662
rect 175188 57598 175240 57604
rect 175096 9648 175148 9654
rect 175096 9590 175148 9596
rect 175004 8900 175056 8906
rect 175004 8842 175056 8848
rect 175200 3369 175228 57598
rect 175292 56846 175320 60044
rect 175568 57866 175596 60044
rect 175556 57860 175608 57866
rect 175556 57802 175608 57808
rect 175280 56840 175332 56846
rect 175280 56782 175332 56788
rect 175844 56778 175872 60044
rect 176134 60030 176332 60058
rect 176410 60030 176608 60058
rect 176304 57644 176332 60030
rect 176304 57616 176516 57644
rect 176384 56840 176436 56846
rect 176384 56782 176436 56788
rect 175740 56772 175792 56778
rect 175740 56714 175792 56720
rect 175832 56772 175884 56778
rect 175832 56714 175884 56720
rect 175280 56568 175332 56574
rect 175280 56510 175332 56516
rect 175292 55214 175320 56510
rect 175752 56438 175780 56714
rect 175740 56432 175792 56438
rect 175740 56374 175792 56380
rect 175292 55186 175596 55214
rect 175568 6914 175596 55186
rect 176396 13938 176424 56782
rect 176488 14006 176516 57616
rect 176580 56930 176608 60030
rect 176672 57730 176700 60044
rect 176660 57724 176712 57730
rect 176660 57666 176712 57672
rect 177040 57662 177068 60044
rect 177132 60030 177330 60058
rect 177028 57656 177080 57662
rect 177028 57598 177080 57604
rect 176580 56902 176792 56930
rect 176764 56778 176792 56902
rect 176568 56772 176620 56778
rect 176568 56714 176620 56720
rect 176752 56772 176804 56778
rect 176752 56714 176804 56720
rect 176476 14000 176528 14006
rect 176476 13942 176528 13948
rect 176384 13932 176436 13938
rect 176384 13874 176436 13880
rect 176580 9586 176608 56714
rect 177132 51406 177160 60030
rect 177592 57882 177620 60044
rect 177882 60030 177988 60058
rect 177592 57854 177896 57882
rect 177500 57730 177804 57746
rect 177488 57724 177804 57730
rect 177540 57718 177804 57724
rect 177488 57666 177540 57672
rect 177580 57656 177632 57662
rect 177580 57598 177632 57604
rect 177672 57656 177724 57662
rect 177672 57598 177724 57604
rect 177120 51400 177172 51406
rect 177120 51342 177172 51348
rect 177592 14074 177620 57598
rect 177684 14142 177712 57598
rect 177672 14136 177724 14142
rect 177672 14078 177724 14084
rect 177580 14068 177632 14074
rect 177580 14010 177632 14016
rect 176568 9580 176620 9586
rect 176568 9522 176620 9528
rect 177776 9518 177804 57718
rect 177764 9512 177816 9518
rect 177764 9454 177816 9460
rect 177868 9382 177896 57854
rect 177960 57662 177988 60030
rect 178144 57730 178172 60044
rect 178132 57724 178184 57730
rect 178132 57666 178184 57672
rect 177948 57656 178000 57662
rect 177948 57598 178000 57604
rect 178132 56432 178184 56438
rect 178132 56374 178184 56380
rect 178040 55956 178092 55962
rect 178040 55898 178092 55904
rect 177948 51400 178000 51406
rect 177948 51342 178000 51348
rect 177960 9450 177988 51342
rect 178052 16574 178080 55898
rect 178144 49298 178172 56374
rect 178420 56302 178448 60044
rect 178788 57662 178816 60044
rect 179078 60030 179184 60058
rect 179052 57724 179104 57730
rect 179052 57666 179104 57672
rect 178776 57656 178828 57662
rect 178776 57598 178828 57604
rect 178408 56296 178460 56302
rect 178408 56238 178460 56244
rect 178132 49292 178184 49298
rect 178132 49234 178184 49240
rect 178052 16546 179000 16574
rect 177948 9444 178000 9450
rect 177948 9386 178000 9392
rect 177856 9376 177908 9382
rect 177856 9318 177908 9324
rect 177856 9036 177908 9042
rect 177856 8978 177908 8984
rect 175476 6886 175596 6914
rect 175186 3360 175242 3369
rect 175186 3295 175242 3304
rect 175476 480 175504 6886
rect 176660 5296 176712 5302
rect 176660 5238 176712 5244
rect 176672 480 176700 5238
rect 177868 480 177896 8978
rect 178972 1986 179000 16546
rect 179064 2106 179092 57666
rect 179156 14210 179184 60030
rect 179236 58132 179288 58138
rect 179236 58074 179288 58080
rect 179248 57798 179276 58074
rect 179236 57792 179288 57798
rect 179236 57734 179288 57740
rect 179236 57656 179288 57662
rect 179236 57598 179288 57604
rect 179144 14204 179196 14210
rect 179144 14146 179196 14152
rect 179248 9314 179276 57598
rect 179340 56166 179368 60044
rect 179616 57662 179644 60044
rect 179604 57656 179656 57662
rect 179604 57598 179656 57604
rect 179892 56710 179920 60044
rect 179880 56704 179932 56710
rect 179880 56646 179932 56652
rect 180260 56506 180288 60044
rect 180550 60030 180656 60058
rect 180826 60030 181024 60058
rect 180432 57656 180484 57662
rect 180432 57598 180484 57604
rect 180248 56500 180300 56506
rect 180248 56442 180300 56448
rect 179328 56160 179380 56166
rect 179328 56102 179380 56108
rect 179236 9308 179288 9314
rect 179236 9250 179288 9256
rect 180444 9246 180472 57598
rect 180524 56704 180576 56710
rect 180524 56646 180576 56652
rect 180536 14278 180564 56646
rect 180524 14272 180576 14278
rect 180524 14214 180576 14220
rect 180432 9240 180484 9246
rect 180432 9182 180484 9188
rect 180628 9178 180656 60030
rect 180996 56914 181024 60030
rect 180892 56908 180944 56914
rect 180892 56850 180944 56856
rect 180984 56908 181036 56914
rect 180984 56850 181036 56856
rect 180706 56808 180762 56817
rect 180904 56778 180932 56850
rect 180706 56743 180708 56752
rect 180760 56743 180762 56752
rect 180892 56772 180944 56778
rect 180708 56714 180760 56720
rect 180892 56714 180944 56720
rect 180800 56704 180852 56710
rect 180798 56672 180800 56681
rect 180852 56672 180854 56681
rect 180798 56607 180854 56616
rect 181088 56234 181116 60044
rect 181378 60030 181576 60058
rect 181654 60030 181944 60058
rect 182022 60030 182128 60058
rect 181076 56228 181128 56234
rect 181076 56170 181128 56176
rect 181548 55214 181576 60030
rect 181916 57644 181944 60030
rect 181916 57616 182036 57644
rect 181904 56908 181956 56914
rect 181904 56850 181956 56856
rect 181548 55186 181852 55214
rect 180616 9172 180668 9178
rect 180616 9114 180668 9120
rect 181824 9110 181852 55186
rect 181916 14346 181944 56850
rect 182008 14414 182036 57616
rect 182100 56438 182128 60030
rect 182284 57662 182312 60044
rect 182272 57656 182324 57662
rect 182272 57598 182324 57604
rect 182560 56914 182588 60044
rect 182548 56908 182600 56914
rect 182548 56850 182600 56856
rect 182088 56432 182140 56438
rect 182088 56374 182140 56380
rect 182836 56370 182864 60044
rect 183112 57866 183140 60044
rect 183204 60030 183402 60058
rect 183008 57860 183060 57866
rect 183008 57802 183060 57808
rect 183100 57860 183152 57866
rect 183100 57802 183152 57808
rect 183020 56778 183048 57802
rect 183100 57656 183152 57662
rect 183100 57598 183152 57604
rect 182916 56772 182968 56778
rect 182916 56714 182968 56720
rect 183008 56772 183060 56778
rect 183008 56714 183060 56720
rect 182928 56574 182956 56714
rect 182916 56568 182968 56574
rect 182916 56510 182968 56516
rect 182824 56364 182876 56370
rect 182824 56306 182876 56312
rect 181996 14408 182048 14414
rect 181996 14350 182048 14356
rect 181904 14340 181956 14346
rect 181904 14282 181956 14288
rect 181812 9104 181864 9110
rect 181812 9046 181864 9052
rect 183112 9042 183140 57598
rect 183204 15094 183232 60030
rect 183376 57860 183428 57866
rect 183376 57802 183428 57808
rect 183284 56908 183336 56914
rect 183284 56850 183336 56856
rect 183296 15162 183324 56850
rect 183284 15156 183336 15162
rect 183284 15098 183336 15104
rect 183192 15088 183244 15094
rect 183192 15030 183244 15036
rect 183100 9036 183152 9042
rect 183100 8978 183152 8984
rect 183388 8974 183416 57802
rect 183756 56098 183784 60044
rect 183848 60030 184046 60058
rect 184322 60030 184520 60058
rect 183744 56092 183796 56098
rect 183744 56034 183796 56040
rect 183848 53310 183876 60030
rect 183928 57656 183980 57662
rect 183928 57598 183980 57604
rect 183940 53378 183968 57598
rect 184204 56568 184256 56574
rect 184204 56510 184256 56516
rect 184388 56568 184440 56574
rect 184388 56510 184440 56516
rect 183928 53372 183980 53378
rect 183928 53314 183980 53320
rect 183836 53304 183888 53310
rect 183836 53246 183888 53252
rect 184216 17678 184244 56510
rect 184400 56234 184428 56510
rect 184388 56228 184440 56234
rect 184388 56170 184440 56176
rect 184492 55214 184520 60030
rect 184584 56234 184612 60044
rect 184860 57662 184888 60044
rect 185136 57866 185164 60044
rect 185124 57860 185176 57866
rect 185124 57802 185176 57808
rect 184848 57656 184900 57662
rect 184848 57598 184900 57604
rect 185032 57656 185084 57662
rect 185032 57598 185084 57604
rect 184572 56228 184624 56234
rect 184572 56170 184624 56176
rect 184492 55186 184612 55214
rect 184204 17672 184256 17678
rect 184204 17614 184256 17620
rect 184584 15026 184612 55186
rect 185044 54602 185072 57598
rect 185504 56030 185532 60044
rect 185780 57662 185808 60044
rect 186070 60030 186176 60058
rect 186044 57860 186096 57866
rect 186044 57802 186096 57808
rect 185768 57656 185820 57662
rect 185768 57598 185820 57604
rect 185492 56024 185544 56030
rect 185492 55966 185544 55972
rect 185032 54596 185084 54602
rect 185032 54538 185084 54544
rect 184572 15020 184624 15026
rect 184572 14962 184624 14968
rect 186056 14958 186084 57802
rect 186044 14952 186096 14958
rect 186044 14894 186096 14900
rect 186148 14890 186176 60030
rect 186332 56914 186360 60044
rect 186320 56908 186372 56914
rect 186320 56850 186372 56856
rect 186608 53242 186636 60044
rect 186898 60030 187188 60058
rect 187266 60030 187464 60058
rect 186780 57860 186832 57866
rect 186780 57802 186832 57808
rect 186792 53582 186820 57802
rect 187160 57644 187188 60030
rect 187436 57746 187464 60030
rect 187528 57866 187556 60044
rect 187712 60030 187818 60058
rect 187516 57860 187568 57866
rect 187516 57802 187568 57808
rect 187436 57718 187556 57746
rect 187160 57616 187464 57644
rect 187240 56908 187292 56914
rect 187240 56850 187292 56856
rect 186780 53576 186832 53582
rect 186780 53518 186832 53524
rect 186596 53236 186648 53242
rect 186596 53178 186648 53184
rect 186136 14884 186188 14890
rect 186136 14826 186188 14832
rect 184940 10940 184992 10946
rect 184940 10882 184992 10888
rect 181444 8968 181496 8974
rect 181444 8910 181496 8916
rect 183376 8968 183428 8974
rect 183376 8910 183428 8916
rect 180248 5228 180300 5234
rect 180248 5170 180300 5176
rect 179052 2100 179104 2106
rect 179052 2042 179104 2048
rect 178972 1958 179092 1986
rect 179064 480 179092 1958
rect 180260 480 180288 5170
rect 181456 480 181484 8910
rect 183744 5160 183796 5166
rect 183744 5102 183796 5108
rect 182548 4480 182600 4486
rect 182548 4422 182600 4428
rect 182560 480 182588 4422
rect 183756 480 183784 5102
rect 184952 480 184980 10882
rect 187252 5166 187280 56850
rect 187436 14822 187464 57616
rect 187424 14816 187476 14822
rect 187424 14758 187476 14764
rect 187240 5160 187292 5166
rect 187240 5102 187292 5108
rect 187332 5092 187384 5098
rect 187332 5034 187384 5040
rect 186136 4412 186188 4418
rect 186136 4354 186188 4360
rect 186148 480 186176 4354
rect 187344 480 187372 5034
rect 187528 4418 187556 57718
rect 187712 50386 187740 60030
rect 188080 57866 188108 60044
rect 188172 60030 188370 60058
rect 188646 60030 188752 60058
rect 188068 57860 188120 57866
rect 188068 57802 188120 57808
rect 188172 53174 188200 60030
rect 188620 57656 188672 57662
rect 188620 57598 188672 57604
rect 188160 53168 188212 53174
rect 188160 53110 188212 53116
rect 187700 50380 187752 50386
rect 187700 50322 187752 50328
rect 188528 10872 188580 10878
rect 188528 10814 188580 10820
rect 187516 4412 187568 4418
rect 187516 4354 187568 4360
rect 188540 480 188568 10814
rect 188632 4486 188660 57598
rect 188724 14686 188752 60030
rect 188896 57860 188948 57866
rect 188896 57802 188948 57808
rect 188804 50380 188856 50386
rect 188804 50322 188856 50328
rect 188816 14754 188844 50322
rect 188804 14748 188856 14754
rect 188804 14690 188856 14696
rect 188712 14680 188764 14686
rect 188712 14622 188764 14628
rect 188908 4554 188936 57802
rect 189000 57662 189028 60044
rect 188988 57656 189040 57662
rect 188988 57598 189040 57604
rect 189276 55962 189304 60044
rect 189552 57866 189580 60044
rect 189842 60030 190040 60058
rect 189540 57860 189592 57866
rect 189540 57802 189592 57808
rect 189356 57656 189408 57662
rect 189356 57598 189408 57604
rect 189264 55956 189316 55962
rect 189264 55898 189316 55904
rect 189368 54534 189396 57598
rect 190012 55214 190040 60030
rect 190104 57662 190132 60044
rect 190196 60030 190394 60058
rect 190092 57656 190144 57662
rect 190092 57598 190144 57604
rect 190012 55186 190132 55214
rect 189356 54528 189408 54534
rect 189356 54470 189408 54476
rect 189724 5024 189776 5030
rect 189724 4966 189776 4972
rect 188896 4548 188948 4554
rect 188896 4490 188948 4496
rect 188620 4480 188672 4486
rect 188620 4422 188672 4428
rect 189736 480 189764 4966
rect 190104 4690 190132 55186
rect 190196 14550 190224 60030
rect 190276 57860 190328 57866
rect 190276 57802 190328 57808
rect 190288 14618 190316 57802
rect 190368 57656 190420 57662
rect 190368 57598 190420 57604
rect 190380 56778 190408 57598
rect 190748 56914 190776 60044
rect 190840 60030 191038 60058
rect 190736 56908 190788 56914
rect 190736 56850 190788 56856
rect 190368 56772 190420 56778
rect 190368 56714 190420 56720
rect 190840 53106 190868 60030
rect 191300 57866 191328 60044
rect 191484 60030 191590 60058
rect 191288 57860 191340 57866
rect 191288 57802 191340 57808
rect 190828 53100 190880 53106
rect 190828 53042 190880 53048
rect 190276 14612 190328 14618
rect 190276 14554 190328 14560
rect 190184 14544 190236 14550
rect 190184 14486 190236 14492
rect 190828 10804 190880 10810
rect 190828 10746 190880 10752
rect 190092 4684 190144 4690
rect 190092 4626 190144 4632
rect 190840 480 190868 10746
rect 191484 5506 191512 60030
rect 191564 57860 191616 57866
rect 191564 57802 191616 57808
rect 191576 14482 191604 57802
rect 191852 56914 191880 60044
rect 191656 56908 191708 56914
rect 191656 56850 191708 56856
rect 191840 56908 191892 56914
rect 191840 56850 191892 56856
rect 191564 14476 191616 14482
rect 191564 14418 191616 14424
rect 191472 5500 191524 5506
rect 191472 5442 191524 5448
rect 191668 4758 191696 56850
rect 192128 51814 192156 60044
rect 192510 60030 192708 60058
rect 192786 60030 192984 60058
rect 192208 57860 192260 57866
rect 192208 57802 192260 57808
rect 192116 51808 192168 51814
rect 192116 51750 192168 51756
rect 192220 50182 192248 57802
rect 192680 55214 192708 60030
rect 192680 55186 192800 55214
rect 192208 50176 192260 50182
rect 192208 50118 192260 50124
rect 192024 10736 192076 10742
rect 192024 10678 192076 10684
rect 191656 4752 191708 4758
rect 191656 4694 191708 4700
rect 192036 480 192064 10678
rect 192772 5438 192800 55186
rect 192956 10266 192984 60030
rect 193048 57866 193076 60044
rect 193036 57860 193088 57866
rect 193036 57802 193088 57808
rect 193220 57860 193272 57866
rect 193220 57802 193272 57808
rect 193036 56908 193088 56914
rect 193036 56850 193088 56856
rect 192944 10260 192996 10266
rect 192944 10202 192996 10208
rect 193048 10198 193076 56850
rect 193232 51746 193260 57802
rect 193324 56778 193352 60044
rect 193600 56914 193628 60044
rect 193876 57866 193904 60044
rect 194152 60030 194258 60058
rect 194336 60030 194534 60058
rect 194704 60030 194810 60058
rect 193864 57860 193916 57866
rect 193864 57802 193916 57808
rect 193588 56908 193640 56914
rect 193588 56850 193640 56856
rect 193312 56772 193364 56778
rect 193312 56714 193364 56720
rect 193220 51740 193272 51746
rect 193220 51682 193272 51688
rect 193220 10668 193272 10674
rect 193220 10610 193272 10616
rect 193036 10192 193088 10198
rect 193036 10134 193088 10140
rect 192760 5432 192812 5438
rect 192760 5374 192812 5380
rect 193232 3262 193260 10610
rect 194152 4962 194180 60030
rect 194232 56908 194284 56914
rect 194232 56850 194284 56856
rect 194244 11014 194272 56850
rect 194232 11008 194284 11014
rect 194232 10950 194284 10956
rect 194336 10946 194364 60030
rect 194600 56908 194652 56914
rect 194600 56850 194652 56856
rect 194416 56772 194468 56778
rect 194416 56714 194468 56720
rect 194324 10940 194376 10946
rect 194324 10882 194376 10888
rect 194428 5370 194456 56714
rect 194612 50658 194640 56850
rect 194600 50652 194652 50658
rect 194600 50594 194652 50600
rect 194704 50522 194732 60030
rect 195072 57866 195100 60044
rect 195362 60030 195652 60058
rect 195060 57860 195112 57866
rect 195060 57802 195112 57808
rect 195624 55214 195652 60030
rect 195716 56914 195744 60044
rect 196006 60030 196112 60058
rect 195888 57860 195940 57866
rect 195888 57802 195940 57808
rect 195704 56908 195756 56914
rect 195704 56850 195756 56856
rect 195624 55186 195836 55214
rect 194692 50516 194744 50522
rect 194692 50458 194744 50464
rect 195808 10878 195836 55186
rect 195796 10872 195848 10878
rect 195796 10814 195848 10820
rect 195612 10600 195664 10606
rect 195612 10542 195664 10548
rect 194416 5364 194468 5370
rect 194416 5306 194468 5312
rect 195336 5160 195388 5166
rect 195336 5102 195388 5108
rect 193312 4956 193364 4962
rect 193312 4898 193364 4904
rect 194140 4956 194192 4962
rect 194140 4898 194192 4904
rect 193220 3256 193272 3262
rect 193220 3198 193272 3204
rect 193324 2530 193352 4898
rect 193864 4888 193916 4894
rect 194048 4888 194100 4894
rect 193916 4848 194048 4876
rect 193864 4830 193916 4836
rect 194048 4830 194100 4836
rect 195060 4820 195112 4826
rect 195060 4762 195112 4768
rect 195072 4622 195100 4762
rect 195060 4616 195112 4622
rect 195060 4558 195112 4564
rect 195152 4616 195204 4622
rect 195152 4558 195204 4564
rect 195164 4486 195192 4558
rect 195152 4480 195204 4486
rect 195152 4422 195204 4428
rect 195348 4418 195376 5102
rect 195336 4412 195388 4418
rect 195336 4354 195388 4360
rect 194416 3256 194468 3262
rect 194416 3198 194468 3204
rect 193232 2502 193352 2530
rect 193232 480 193260 2502
rect 194428 480 194456 3198
rect 195624 480 195652 10542
rect 195900 5234 195928 57802
rect 196084 50386 196112 60030
rect 196268 57866 196296 60044
rect 196452 60030 196558 60058
rect 196834 60030 196940 60058
rect 196256 57860 196308 57866
rect 196256 57802 196308 57808
rect 196452 50726 196480 60030
rect 196440 50720 196492 50726
rect 196440 50662 196492 50668
rect 196072 50380 196124 50386
rect 196072 50322 196124 50328
rect 196912 5302 196940 60030
rect 196992 57860 197044 57866
rect 196992 57802 197044 57808
rect 197004 10810 197032 57802
rect 196992 10804 197044 10810
rect 196992 10746 197044 10752
rect 197096 10742 197124 60044
rect 197478 60030 197584 60058
rect 197360 57860 197412 57866
rect 197360 57802 197412 57808
rect 197176 50380 197228 50386
rect 197176 50322 197228 50328
rect 197084 10736 197136 10742
rect 197084 10678 197136 10684
rect 196900 5296 196952 5302
rect 196900 5238 196952 5244
rect 195888 5228 195940 5234
rect 195888 5170 195940 5176
rect 197188 5166 197216 50322
rect 197372 49026 197400 57802
rect 197556 50590 197584 60030
rect 197740 56778 197768 60044
rect 198030 60030 198228 60058
rect 198200 57610 198228 60030
rect 198292 57866 198320 60044
rect 198280 57860 198332 57866
rect 198280 57802 198332 57808
rect 198200 57582 198504 57610
rect 198280 56908 198332 56914
rect 198280 56850 198332 56856
rect 197728 56772 197780 56778
rect 197728 56714 197780 56720
rect 197544 50584 197596 50590
rect 197544 50526 197596 50532
rect 197360 49020 197412 49026
rect 197360 48962 197412 48968
rect 197912 10532 197964 10538
rect 197912 10474 197964 10480
rect 197176 5160 197228 5166
rect 197176 5102 197228 5108
rect 196808 4888 196860 4894
rect 196808 4830 196860 4836
rect 196820 480 196848 4830
rect 197924 480 197952 10474
rect 198292 4962 198320 56850
rect 198476 10674 198504 57582
rect 198568 56914 198596 60044
rect 198844 57866 198872 60044
rect 198832 57860 198884 57866
rect 198832 57802 198884 57808
rect 198556 56908 198608 56914
rect 198556 56850 198608 56856
rect 198740 56908 198792 56914
rect 198740 56850 198792 56856
rect 198556 56772 198608 56778
rect 198556 56714 198608 56720
rect 198464 10668 198516 10674
rect 198464 10610 198516 10616
rect 198568 5030 198596 56714
rect 198752 50386 198780 56850
rect 199212 50454 199240 60044
rect 199502 60030 199700 60058
rect 199778 60030 199976 60058
rect 199200 50448 199252 50454
rect 199200 50390 199252 50396
rect 198740 50380 198792 50386
rect 198740 50322 198792 50328
rect 199108 10464 199160 10470
rect 199108 10406 199160 10412
rect 198556 5024 198608 5030
rect 198556 4966 198608 4972
rect 198280 4956 198332 4962
rect 198280 4898 198332 4904
rect 199120 480 199148 10406
rect 199672 5137 199700 60030
rect 199844 57860 199896 57866
rect 199844 57802 199896 57808
rect 199752 50380 199804 50386
rect 199752 50322 199804 50328
rect 199764 16114 199792 50322
rect 199752 16108 199804 16114
rect 199752 16050 199804 16056
rect 199856 10606 199884 57802
rect 199844 10600 199896 10606
rect 199844 10542 199896 10548
rect 199948 10538 199976 60030
rect 200040 56914 200068 60044
rect 200132 60030 200330 60058
rect 200028 56908 200080 56914
rect 200028 56850 200080 56856
rect 200028 50516 200080 50522
rect 200028 50458 200080 50464
rect 200040 50182 200068 50458
rect 200132 50182 200160 60030
rect 200592 57798 200620 60044
rect 200974 60030 201172 60058
rect 201250 60030 201448 60058
rect 201526 60030 201632 60058
rect 200488 57792 200540 57798
rect 200488 57734 200540 57740
rect 200580 57792 200632 57798
rect 200580 57734 200632 57740
rect 200500 56778 200528 57734
rect 200488 56772 200540 56778
rect 200488 56714 200540 56720
rect 200028 50176 200080 50182
rect 200028 50118 200080 50124
rect 200120 50176 200172 50182
rect 200120 50118 200172 50124
rect 201144 16046 201172 60030
rect 201224 57792 201276 57798
rect 201224 57734 201276 57740
rect 201132 16040 201184 16046
rect 201132 15982 201184 15988
rect 199936 10532 199988 10538
rect 199936 10474 199988 10480
rect 201236 10470 201264 57734
rect 201316 50176 201368 50182
rect 201316 50118 201368 50124
rect 201224 10464 201276 10470
rect 201224 10406 201276 10412
rect 199658 5128 199714 5137
rect 201328 5098 201356 50118
rect 199658 5063 199714 5072
rect 200304 5092 200356 5098
rect 200304 5034 200356 5040
rect 201316 5092 201368 5098
rect 201316 5034 201368 5040
rect 200316 480 200344 5034
rect 201420 5001 201448 60030
rect 201604 50114 201632 60030
rect 201788 57866 201816 60044
rect 201776 57860 201828 57866
rect 201776 57802 201828 57808
rect 201684 57792 201736 57798
rect 201684 57734 201736 57740
rect 201696 50182 201724 57734
rect 202064 57390 202092 60044
rect 202340 57798 202368 60044
rect 202432 60030 202722 60058
rect 202328 57792 202380 57798
rect 202328 57734 202380 57740
rect 201776 57384 201828 57390
rect 201776 57326 201828 57332
rect 202052 57384 202104 57390
rect 202052 57326 202104 57332
rect 201788 56914 201816 57326
rect 201776 56908 201828 56914
rect 201776 56850 201828 56856
rect 201684 50176 201736 50182
rect 201684 50118 201736 50124
rect 201592 50108 201644 50114
rect 201592 50050 201644 50056
rect 202432 15910 202460 60030
rect 202984 57866 203012 60044
rect 202512 57860 202564 57866
rect 202512 57802 202564 57808
rect 202972 57860 203024 57866
rect 202972 57802 203024 57808
rect 202524 15978 202552 57802
rect 203260 57798 203288 60044
rect 203248 57792 203300 57798
rect 203248 57734 203300 57740
rect 202788 57384 202840 57390
rect 202788 57326 202840 57332
rect 202604 50176 202656 50182
rect 202604 50118 202656 50124
rect 202512 15972 202564 15978
rect 202512 15914 202564 15920
rect 202420 15904 202472 15910
rect 202420 15846 202472 15852
rect 202616 14906 202644 50118
rect 202696 50108 202748 50114
rect 202696 50050 202748 50056
rect 202524 14878 202644 14906
rect 202524 10334 202552 14878
rect 202708 10588 202736 50050
rect 202800 10690 202828 57326
rect 203536 57225 203564 60044
rect 203812 59294 203840 60044
rect 203996 60030 204102 60058
rect 203800 59288 203852 59294
rect 203800 59230 203852 59236
rect 203996 57390 204024 60030
rect 204168 57860 204220 57866
rect 204168 57802 204220 57808
rect 204076 57792 204128 57798
rect 204076 57734 204128 57740
rect 203984 57384 204036 57390
rect 203984 57326 204036 57332
rect 203522 57216 203578 57225
rect 203522 57151 203578 57160
rect 203524 56908 203576 56914
rect 203524 56850 203576 56856
rect 202800 10662 203012 10690
rect 202708 10560 202920 10588
rect 202892 10402 202920 10560
rect 202696 10396 202748 10402
rect 202696 10338 202748 10344
rect 202880 10396 202932 10402
rect 202880 10338 202932 10344
rect 201592 10328 201644 10334
rect 201592 10270 201644 10276
rect 202512 10328 202564 10334
rect 202512 10270 202564 10276
rect 201406 4992 201462 5001
rect 201406 4927 201462 4936
rect 201604 3482 201632 10270
rect 201512 3454 201632 3482
rect 201512 480 201540 3454
rect 202708 480 202736 10338
rect 202984 10282 203012 10662
rect 202800 10254 203012 10282
rect 202800 4865 202828 10254
rect 202786 4856 202842 4865
rect 202786 4791 202842 4800
rect 203536 3262 203564 56850
rect 204088 6225 204116 57734
rect 204074 6216 204130 6225
rect 204074 6151 204130 6160
rect 204180 4826 204208 57802
rect 204456 56817 204484 60044
rect 204732 59809 204760 60044
rect 204718 59800 204774 59809
rect 204718 59735 204774 59744
rect 205008 58138 205036 60044
rect 204996 58132 205048 58138
rect 204996 58074 205048 58080
rect 205284 56914 205312 60044
rect 205560 59430 205588 60044
rect 205548 59424 205600 59430
rect 205548 59366 205600 59372
rect 205836 58274 205864 60044
rect 206204 58721 206232 60044
rect 206190 58712 206246 58721
rect 206190 58647 206246 58656
rect 205824 58268 205876 58274
rect 205824 58210 205876 58216
rect 204720 56908 204772 56914
rect 204720 56850 204772 56856
rect 205272 56908 205324 56914
rect 205272 56850 205324 56856
rect 204442 56808 204498 56817
rect 204442 56743 204498 56752
rect 204732 56710 204760 56850
rect 204812 56840 204864 56846
rect 204864 56800 204944 56828
rect 204812 56782 204864 56788
rect 204720 56704 204772 56710
rect 204720 56646 204772 56652
rect 204916 20126 204944 56800
rect 206480 56778 206508 60044
rect 206756 57633 206784 60044
rect 207032 57769 207060 60044
rect 207308 59498 207336 60044
rect 207296 59492 207348 59498
rect 207296 59434 207348 59440
rect 207584 59022 207612 60044
rect 207966 60030 208164 60058
rect 208136 59906 208164 60030
rect 208124 59900 208176 59906
rect 208124 59842 208176 59848
rect 207572 59016 207624 59022
rect 207572 58958 207624 58964
rect 208228 58954 208256 60044
rect 208216 58948 208268 58954
rect 208216 58890 208268 58896
rect 208504 57866 208532 60044
rect 208492 57860 208544 57866
rect 208492 57802 208544 57808
rect 207018 57760 207074 57769
rect 207018 57695 207074 57704
rect 206742 57624 206798 57633
rect 206742 57559 206798 57568
rect 208492 57384 208544 57390
rect 208492 57326 208544 57332
rect 206468 56772 206520 56778
rect 206468 56714 206520 56720
rect 208504 56710 208532 57326
rect 208780 56953 208808 60044
rect 209056 59673 209084 60044
rect 209042 59664 209098 59673
rect 209042 59599 209098 59608
rect 209332 58886 209360 60044
rect 209320 58880 209372 58886
rect 209320 58822 209372 58828
rect 209700 57497 209728 60044
rect 209976 57769 210004 60044
rect 209962 57760 210018 57769
rect 209962 57695 210018 57704
rect 209686 57488 209742 57497
rect 209686 57423 209742 57432
rect 210252 57390 210280 60044
rect 210528 57905 210556 60044
rect 210804 58478 210832 60044
rect 210792 58472 210844 58478
rect 210792 58414 210844 58420
rect 210514 57896 210570 57905
rect 210514 57831 210570 57840
rect 210884 57792 210936 57798
rect 210884 57734 210936 57740
rect 210240 57384 210292 57390
rect 210240 57326 210292 57332
rect 210896 57186 210924 57734
rect 210884 57180 210936 57186
rect 210884 57122 210936 57128
rect 208766 56944 208822 56953
rect 208766 56879 208822 56888
rect 209872 56840 209924 56846
rect 209872 56782 209924 56788
rect 208400 56704 208452 56710
rect 208400 56646 208452 56652
rect 208492 56704 208544 56710
rect 208492 56646 208544 56652
rect 207020 55480 207072 55486
rect 207020 55422 207072 55428
rect 204904 20120 204956 20126
rect 204904 20062 204956 20068
rect 207032 16574 207060 55422
rect 208412 55214 208440 56646
rect 209780 55412 209832 55418
rect 209780 55354 209832 55360
rect 208412 55186 209084 55214
rect 209056 20058 209084 55186
rect 209044 20052 209096 20058
rect 209044 19994 209096 20000
rect 207032 16546 207428 16574
rect 205088 9784 205140 9790
rect 205088 9726 205140 9732
rect 204732 5358 205036 5386
rect 204732 4894 204760 5358
rect 205008 5302 205036 5358
rect 204904 5296 204956 5302
rect 204904 5238 204956 5244
rect 204996 5296 205048 5302
rect 204996 5238 205048 5244
rect 204916 5098 204944 5238
rect 204812 5092 204864 5098
rect 204812 5034 204864 5040
rect 204904 5092 204956 5098
rect 204904 5034 204956 5040
rect 204720 4888 204772 4894
rect 204720 4830 204772 4836
rect 204824 4842 204852 5034
rect 204996 4888 205048 4894
rect 204824 4836 204996 4842
rect 204824 4830 205048 4836
rect 203892 4820 203944 4826
rect 203892 4762 203944 4768
rect 204168 4820 204220 4826
rect 204824 4814 205036 4830
rect 204168 4762 204220 4768
rect 203524 3256 203576 3262
rect 203524 3198 203576 3204
rect 203904 480 203932 4762
rect 205100 480 205128 9726
rect 206192 3256 206244 3262
rect 206192 3198 206244 3204
rect 206204 480 206232 3198
rect 207400 480 207428 16546
rect 209792 11150 209820 55354
rect 209884 55214 209912 56782
rect 211172 56681 211200 60044
rect 211448 57905 211476 60044
rect 211738 60030 211894 60058
rect 223578 60072 223634 60081
rect 211894 60007 211950 60016
rect 212000 58682 212028 60044
rect 211988 58676 212040 58682
rect 211988 58618 212040 58624
rect 211434 57896 211490 57905
rect 211434 57831 211490 57840
rect 212276 57186 212304 60044
rect 212448 59696 212500 59702
rect 212448 59638 212500 59644
rect 212460 59430 212488 59638
rect 212448 59424 212500 59430
rect 212448 59366 212500 59372
rect 212552 58342 212580 60044
rect 212920 59362 212948 60044
rect 213210 60030 213408 60058
rect 212908 59356 212960 59362
rect 212908 59298 212960 59304
rect 212540 58336 212592 58342
rect 212540 58278 212592 58284
rect 213184 57928 213236 57934
rect 213184 57870 213236 57876
rect 212264 57180 212316 57186
rect 212264 57122 212316 57128
rect 211158 56672 211214 56681
rect 211158 56607 211214 56616
rect 209884 55186 210464 55214
rect 209872 15360 209924 15366
rect 209872 15302 209924 15308
rect 209780 11144 209832 11150
rect 209780 11086 209832 11092
rect 208584 9852 208636 9858
rect 208584 9794 208636 9800
rect 208596 480 208624 9794
rect 209884 3482 209912 15302
rect 210436 6633 210464 55186
rect 213092 15428 213144 15434
rect 213092 15370 213144 15376
rect 210976 11144 211028 11150
rect 210976 11086 211028 11092
rect 210422 6624 210478 6633
rect 210422 6559 210478 6568
rect 209792 3454 209912 3482
rect 209792 480 209820 3454
rect 210988 480 211016 11086
rect 212172 9920 212224 9926
rect 212172 9862 212224 9868
rect 212184 480 212212 9862
rect 213104 3482 213132 15370
rect 213196 4049 213224 57870
rect 213380 57730 213408 60030
rect 213276 57724 213328 57730
rect 213276 57666 213328 57672
rect 213368 57724 213420 57730
rect 213368 57666 213420 57672
rect 213288 18630 213316 57666
rect 213368 57112 213420 57118
rect 213368 57054 213420 57060
rect 213276 18624 213328 18630
rect 213276 18566 213328 18572
rect 213380 16574 213408 57054
rect 213472 56846 213500 60044
rect 213748 57186 213776 60044
rect 213828 59628 213880 59634
rect 213828 59570 213880 59576
rect 213736 57180 213788 57186
rect 213736 57122 213788 57128
rect 213552 56976 213604 56982
rect 213552 56918 213604 56924
rect 213460 56840 213512 56846
rect 213460 56782 213512 56788
rect 213380 16546 213500 16574
rect 213182 4040 213238 4049
rect 213182 3975 213238 3984
rect 213104 3454 213408 3482
rect 213380 480 213408 3454
rect 213472 3097 213500 16546
rect 213564 3233 213592 56918
rect 213840 56914 213868 59570
rect 214024 58206 214052 60044
rect 214314 60030 214604 60058
rect 214576 59838 214604 60030
rect 214564 59832 214616 59838
rect 214564 59774 214616 59780
rect 214668 58585 214696 60044
rect 214944 58614 214972 60044
rect 214932 58608 214984 58614
rect 214654 58576 214710 58585
rect 214932 58550 214984 58556
rect 214654 58511 214710 58520
rect 214012 58200 214064 58206
rect 214012 58142 214064 58148
rect 215220 57730 215248 60044
rect 215116 57724 215168 57730
rect 215116 57666 215168 57672
rect 215208 57724 215260 57730
rect 215208 57666 215260 57672
rect 215128 57526 215156 57666
rect 214564 57520 214616 57526
rect 214564 57462 214616 57468
rect 215116 57520 215168 57526
rect 215116 57462 215168 57468
rect 214380 57384 214432 57390
rect 214380 57326 214432 57332
rect 214472 57384 214524 57390
rect 214472 57326 214524 57332
rect 213828 56908 213880 56914
rect 213828 56850 213880 56856
rect 214392 56658 214420 57326
rect 214484 56778 214512 57326
rect 214576 57050 214604 57462
rect 215496 57118 215524 60044
rect 215772 59294 215800 60044
rect 215760 59288 215812 59294
rect 215760 59230 215812 59236
rect 216048 57934 216076 60044
rect 216416 58818 216444 60044
rect 216404 58812 216456 58818
rect 216404 58754 216456 58760
rect 216692 58750 216720 60044
rect 216968 59362 216996 60044
rect 216956 59356 217008 59362
rect 216956 59298 217008 59304
rect 216680 58744 216732 58750
rect 216680 58686 216732 58692
rect 216036 57928 216088 57934
rect 216036 57870 216088 57876
rect 217244 57662 217272 60044
rect 217520 58410 217548 60044
rect 217796 58546 217824 60044
rect 218060 59764 218112 59770
rect 218060 59706 218112 59712
rect 217784 58540 217836 58546
rect 217784 58482 217836 58488
rect 217508 58404 217560 58410
rect 217508 58346 217560 58352
rect 218072 57866 218100 59706
rect 218164 59265 218192 60044
rect 218150 59256 218206 59265
rect 218440 59226 218468 60044
rect 218150 59191 218206 59200
rect 218428 59220 218480 59226
rect 218428 59162 218480 59168
rect 218716 58993 218744 60044
rect 218702 58984 218758 58993
rect 218702 58919 218758 58928
rect 218060 57860 218112 57866
rect 218060 57802 218112 57808
rect 216036 57656 216088 57662
rect 216036 57598 216088 57604
rect 217232 57656 217284 57662
rect 217232 57598 217284 57604
rect 215392 57112 215444 57118
rect 215392 57054 215444 57060
rect 215484 57112 215536 57118
rect 215484 57054 215536 57060
rect 214564 57044 214616 57050
rect 214564 56986 214616 56992
rect 214748 56908 214800 56914
rect 214748 56850 214800 56856
rect 214472 56772 214524 56778
rect 214472 56714 214524 56720
rect 214656 56772 214708 56778
rect 214656 56714 214708 56720
rect 214668 56658 214696 56714
rect 214760 56710 214788 56850
rect 215404 56710 215432 57054
rect 215944 56976 215996 56982
rect 215944 56918 215996 56924
rect 214392 56630 214696 56658
rect 214748 56704 214800 56710
rect 214748 56646 214800 56652
rect 215392 56704 215444 56710
rect 215392 56646 215444 56652
rect 213920 55548 213972 55554
rect 213920 55490 213972 55496
rect 213932 16574 213960 55490
rect 213932 16546 214512 16574
rect 213550 3224 213606 3233
rect 213550 3159 213606 3168
rect 213458 3088 213514 3097
rect 213458 3023 213514 3032
rect 214484 480 214512 16546
rect 215668 9988 215720 9994
rect 215668 9930 215720 9936
rect 215680 480 215708 9930
rect 215956 4078 215984 56918
rect 216048 19990 216076 57598
rect 216772 57520 216824 57526
rect 216772 57462 216824 57468
rect 216784 57186 216812 57462
rect 216772 57180 216824 57186
rect 216772 57122 216824 57128
rect 216588 57112 216640 57118
rect 218992 57089 219020 60044
rect 219268 59129 219296 60044
rect 219558 60030 219848 60058
rect 219254 59120 219310 59129
rect 219254 59055 219310 59064
rect 219622 58984 219678 58993
rect 219622 58919 219678 58928
rect 219636 58585 219664 58919
rect 219622 58576 219678 58585
rect 219440 58540 219492 58546
rect 219622 58511 219678 58520
rect 219440 58482 219492 58488
rect 219452 58426 219480 58482
rect 219452 58398 219572 58426
rect 219544 58138 219572 58398
rect 219532 58132 219584 58138
rect 219532 58074 219584 58080
rect 219820 58070 219848 60030
rect 219808 58064 219860 58070
rect 219808 58006 219860 58012
rect 219254 57760 219310 57769
rect 219254 57695 219310 57704
rect 219268 57610 219296 57695
rect 219268 57582 219480 57610
rect 219452 57526 219480 57582
rect 219440 57520 219492 57526
rect 219440 57462 219492 57468
rect 216588 57054 216640 57060
rect 218978 57080 219034 57089
rect 216600 56982 216628 57054
rect 218978 57015 219034 57024
rect 216588 56976 216640 56982
rect 216588 56918 216640 56924
rect 216496 56840 216548 56846
rect 216324 56788 216496 56794
rect 216324 56782 216548 56788
rect 216324 56778 216536 56782
rect 216312 56772 216536 56778
rect 216364 56766 216536 56772
rect 216312 56714 216364 56720
rect 219912 56642 219940 60044
rect 220188 59265 220216 60044
rect 220174 59256 220230 59265
rect 220174 59191 220230 59200
rect 220464 57905 220492 60044
rect 220450 57896 220506 57905
rect 220450 57831 220506 57840
rect 220176 57792 220228 57798
rect 220176 57734 220228 57740
rect 219624 56636 219676 56642
rect 219624 56578 219676 56584
rect 219900 56636 219952 56642
rect 219900 56578 219952 56584
rect 219636 55214 219664 56578
rect 219636 55186 220124 55214
rect 218060 54256 218112 54262
rect 218060 54198 218112 54204
rect 216036 19984 216088 19990
rect 216036 19926 216088 19932
rect 216864 15496 216916 15502
rect 216864 15438 216916 15444
rect 215944 4072 215996 4078
rect 215944 4014 215996 4020
rect 216876 480 216904 15438
rect 218072 480 218100 54198
rect 219992 15564 220044 15570
rect 219992 15506 220044 15512
rect 219256 10056 219308 10062
rect 219256 9998 219308 10004
rect 219268 480 219296 9998
rect 220004 2802 220032 15506
rect 220096 3262 220124 55186
rect 220188 4146 220216 57734
rect 220740 57050 220768 60044
rect 221016 59294 221044 60044
rect 221004 59288 221056 59294
rect 221004 59230 221056 59236
rect 221292 57934 221320 60044
rect 221660 59401 221688 60044
rect 221646 59392 221702 59401
rect 221646 59327 221702 59336
rect 221830 58304 221886 58313
rect 221830 58239 221886 58248
rect 221844 58206 221872 58239
rect 221936 58206 221964 60044
rect 221832 58200 221884 58206
rect 221832 58142 221884 58148
rect 221924 58200 221976 58206
rect 221924 58142 221976 58148
rect 221280 57928 221332 57934
rect 221280 57870 221332 57876
rect 221832 57860 221884 57866
rect 221832 57802 221884 57808
rect 220268 57044 220320 57050
rect 220268 56986 220320 56992
rect 220728 57044 220780 57050
rect 220728 56986 220780 56992
rect 220176 4140 220228 4146
rect 220176 4082 220228 4088
rect 220084 3256 220136 3262
rect 220084 3198 220136 3204
rect 220280 2990 220308 56986
rect 221844 56710 221872 57802
rect 222212 57186 222240 60044
rect 222764 59537 222792 60044
rect 222750 59528 222806 59537
rect 222750 59463 222806 59472
rect 222476 58880 222528 58886
rect 222476 58822 222528 58828
rect 222292 58608 222344 58614
rect 222292 58550 222344 58556
rect 222304 58342 222332 58550
rect 222488 58478 222516 58822
rect 222384 58472 222436 58478
rect 222384 58414 222436 58420
rect 222476 58472 222528 58478
rect 222476 58414 222528 58420
rect 222396 58342 222424 58414
rect 222292 58336 222344 58342
rect 222292 58278 222344 58284
rect 222384 58336 222436 58342
rect 222384 58278 222436 58284
rect 223040 57866 223068 60044
rect 223422 60030 223578 60058
rect 223698 60030 223896 60058
rect 223578 60007 223634 60016
rect 223868 59906 223896 60030
rect 223856 59900 223908 59906
rect 223856 59842 223908 59848
rect 223960 59430 223988 60044
rect 224250 60030 224448 60058
rect 224420 59809 224448 60030
rect 224406 59800 224462 59809
rect 224406 59735 224462 59744
rect 224132 59560 224184 59566
rect 224132 59502 224184 59508
rect 223948 59424 224000 59430
rect 223948 59366 224000 59372
rect 223578 59120 223634 59129
rect 223396 59084 223448 59090
rect 223578 59055 223634 59064
rect 223946 59120 224002 59129
rect 223946 59055 224002 59064
rect 223396 59026 223448 59032
rect 222936 57860 222988 57866
rect 222936 57802 222988 57808
rect 223028 57860 223080 57866
rect 223028 57802 223080 57808
rect 222948 57746 222976 57802
rect 222948 57718 223068 57746
rect 223408 57730 223436 59026
rect 223486 57760 223542 57769
rect 223040 57594 223068 57718
rect 223396 57724 223448 57730
rect 223592 57746 223620 59055
rect 223764 58880 223816 58886
rect 223764 58822 223816 58828
rect 223776 58274 223804 58822
rect 223764 58268 223816 58274
rect 223764 58210 223816 58216
rect 223542 57718 223620 57746
rect 223486 57695 223542 57704
rect 223396 57666 223448 57672
rect 223960 57662 223988 59055
rect 223948 57656 224000 57662
rect 223948 57598 224000 57604
rect 222936 57588 222988 57594
rect 222936 57530 222988 57536
rect 223028 57588 223080 57594
rect 223028 57530 223080 57536
rect 222384 57452 222436 57458
rect 222384 57394 222436 57400
rect 222200 57180 222252 57186
rect 222200 57122 222252 57128
rect 222016 57112 222068 57118
rect 222016 57054 222068 57060
rect 222028 56846 222056 57054
rect 221924 56840 221976 56846
rect 221924 56782 221976 56788
rect 222016 56840 222068 56846
rect 222016 56782 222068 56788
rect 221936 56710 221964 56782
rect 221832 56704 221884 56710
rect 221832 56646 221884 56652
rect 221924 56704 221976 56710
rect 221924 56646 221976 56652
rect 220820 55616 220872 55622
rect 220820 55558 220872 55564
rect 220832 16574 220860 55558
rect 222396 55214 222424 57394
rect 222396 55186 222884 55214
rect 220832 16546 221596 16574
rect 220268 2984 220320 2990
rect 220268 2926 220320 2932
rect 220004 2774 220492 2802
rect 220464 480 220492 2774
rect 221568 480 221596 16546
rect 222752 10124 222804 10130
rect 222752 10066 222804 10072
rect 222764 480 222792 10066
rect 222856 2922 222884 55186
rect 222948 3058 222976 57530
rect 223028 57316 223080 57322
rect 223028 57258 223080 57264
rect 222936 3052 222988 3058
rect 222936 2994 222988 3000
rect 222844 2916 222896 2922
rect 222844 2858 222896 2864
rect 223040 2854 223068 57258
rect 224144 57118 224172 59502
rect 224788 59362 224816 398550
rect 224868 398472 224920 398478
rect 224868 398414 224920 398420
rect 224776 59356 224828 59362
rect 224776 59298 224828 59304
rect 224314 59120 224370 59129
rect 224314 59055 224370 59064
rect 224224 58744 224276 58750
rect 224224 58686 224276 58692
rect 224236 58274 224264 58686
rect 224224 58268 224276 58274
rect 224224 58210 224276 58216
rect 224328 57798 224356 59055
rect 224408 58744 224460 58750
rect 224408 58686 224460 58692
rect 224420 58313 224448 58686
rect 224880 58546 224908 398414
rect 224972 59226 225000 398618
rect 225052 397248 225104 397254
rect 225052 397190 225104 397196
rect 224960 59220 225012 59226
rect 224960 59162 225012 59168
rect 224868 58540 224920 58546
rect 224868 58482 224920 58488
rect 224406 58304 224462 58313
rect 224406 58239 224462 58248
rect 225064 58002 225092 397190
rect 225144 266144 225196 266150
rect 225144 266086 225196 266092
rect 225052 57996 225104 58002
rect 225052 57938 225104 57944
rect 224316 57792 224368 57798
rect 224316 57734 224368 57740
rect 225156 57497 225184 266086
rect 226064 261316 226116 261322
rect 226064 261258 226116 261264
rect 225236 260432 225288 260438
rect 225236 260374 225288 260380
rect 225248 64161 225276 260374
rect 225326 244896 225382 244905
rect 225326 244831 225382 244840
rect 225234 64152 225290 64161
rect 225234 64087 225290 64096
rect 225340 60489 225368 244831
rect 225418 240816 225474 240825
rect 225418 240751 225474 240760
rect 225326 60480 225382 60489
rect 225326 60415 225382 60424
rect 225326 60344 225382 60353
rect 225326 60279 225382 60288
rect 225234 60208 225290 60217
rect 225234 60143 225290 60152
rect 225248 59090 225276 60143
rect 225236 59084 225288 59090
rect 225236 59026 225288 59032
rect 225142 57488 225198 57497
rect 225142 57423 225198 57432
rect 225340 57390 225368 60279
rect 225432 59906 225460 240751
rect 225510 238096 225566 238105
rect 225510 238031 225566 238040
rect 225420 59900 225472 59906
rect 225420 59842 225472 59848
rect 225524 59786 225552 238031
rect 225786 232792 225842 232801
rect 225786 232727 225842 232736
rect 225694 232656 225750 232665
rect 225694 232591 225750 232600
rect 225602 232520 225658 232529
rect 225602 232455 225658 232464
rect 225432 59758 225552 59786
rect 225328 57384 225380 57390
rect 225328 57326 225380 57332
rect 224132 57112 224184 57118
rect 224132 57054 224184 57060
rect 225432 56681 225460 59758
rect 225616 57633 225644 232455
rect 225708 62801 225736 232591
rect 225800 65657 225828 232727
rect 225878 231432 225934 231441
rect 225878 231367 225934 231376
rect 225786 65648 225842 65657
rect 225786 65583 225842 65592
rect 225892 65521 225920 231367
rect 225970 228304 226026 228313
rect 225970 228239 226026 228248
rect 225984 65657 226012 228239
rect 226076 132433 226104 261258
rect 226156 260704 226208 260710
rect 226156 260646 226208 260652
rect 226168 143585 226196 260646
rect 226246 250472 226302 250481
rect 226246 250407 226302 250416
rect 226260 148889 226288 250407
rect 226338 231568 226394 231577
rect 226338 231503 226394 231512
rect 226352 222737 226380 231503
rect 226338 222728 226394 222737
rect 226338 222663 226394 222672
rect 226338 204232 226394 204241
rect 226338 204167 226394 204176
rect 226352 203561 226380 204167
rect 226338 203552 226394 203561
rect 226338 203487 226394 203496
rect 226246 148880 226302 148889
rect 226246 148815 226302 148824
rect 226246 147792 226302 147801
rect 226246 147727 226302 147736
rect 226154 143576 226210 143585
rect 226154 143511 226210 143520
rect 226154 143440 226210 143449
rect 226154 143375 226210 143384
rect 226062 132424 226118 132433
rect 226062 132359 226118 132368
rect 225970 65648 226026 65657
rect 225970 65583 226026 65592
rect 225878 65512 225934 65521
rect 225878 65447 225934 65456
rect 226062 65512 226118 65521
rect 226062 65447 226118 65456
rect 225970 65376 226026 65385
rect 225970 65311 226026 65320
rect 225786 65240 225842 65249
rect 225786 65175 225842 65184
rect 225694 62792 225750 62801
rect 225694 62727 225750 62736
rect 225694 60480 225750 60489
rect 225694 60415 225750 60424
rect 225602 57624 225658 57633
rect 225602 57559 225658 57568
rect 225708 56778 225736 60415
rect 225800 57934 225828 65175
rect 225878 62792 225934 62801
rect 225878 62727 225934 62736
rect 225788 57928 225840 57934
rect 225788 57870 225840 57876
rect 225892 57594 225920 62727
rect 225880 57588 225932 57594
rect 225880 57530 225932 57536
rect 225696 56772 225748 56778
rect 225696 56714 225748 56720
rect 225984 56710 226012 65311
rect 226076 60081 226104 65447
rect 226062 60072 226118 60081
rect 226062 60007 226118 60016
rect 226064 59900 226116 59906
rect 226064 59842 226116 59848
rect 226076 59566 226104 59842
rect 226064 59560 226116 59566
rect 226064 59502 226116 59508
rect 226168 57526 226196 143375
rect 226156 57520 226208 57526
rect 226156 57462 226208 57468
rect 226260 56846 226288 147727
rect 226444 146169 226472 399842
rect 226524 399832 226576 399838
rect 226524 399774 226576 399780
rect 226536 181801 226564 399774
rect 226984 396432 227036 396438
rect 226984 396374 227036 396380
rect 226996 261390 227024 396374
rect 226984 261384 227036 261390
rect 226984 261326 227036 261332
rect 226982 239456 227038 239465
rect 226982 239391 227038 239400
rect 226614 235240 226670 235249
rect 226614 235175 226670 235184
rect 226522 181792 226578 181801
rect 226522 181727 226578 181736
rect 226430 146160 226486 146169
rect 226430 146095 226486 146104
rect 226628 138009 226656 235175
rect 226798 231296 226854 231305
rect 226798 231231 226854 231240
rect 226706 231160 226762 231169
rect 226706 231095 226762 231104
rect 226614 138000 226670 138009
rect 226614 137935 226670 137944
rect 226720 135289 226748 231095
rect 226812 151609 226840 231231
rect 226890 226128 226946 226137
rect 226890 226063 226946 226072
rect 226904 154329 226932 226063
rect 226996 168065 227024 239391
rect 227074 236736 227130 236745
rect 227074 236671 227130 236680
rect 227088 176225 227116 236671
rect 227166 234016 227222 234025
rect 227166 233951 227222 233960
rect 227180 192681 227208 233951
rect 227258 227080 227314 227089
rect 227258 227015 227314 227024
rect 227166 192672 227222 192681
rect 227166 192607 227222 192616
rect 227272 187241 227300 227015
rect 227258 187232 227314 187241
rect 227258 187167 227314 187176
rect 227074 176216 227130 176225
rect 227074 176151 227130 176160
rect 226982 168056 227038 168065
rect 226982 167991 227038 168000
rect 226890 154320 226946 154329
rect 226890 154255 226946 154264
rect 226798 151600 226854 151609
rect 226798 151535 226854 151544
rect 226706 135280 226762 135289
rect 226706 135215 226762 135224
rect 226522 125488 226578 125497
rect 226522 125423 226578 125432
rect 226536 124273 226564 125423
rect 226522 124264 226578 124273
rect 226522 124199 226578 124208
rect 226522 122768 226578 122777
rect 226522 122703 226578 122712
rect 226536 121553 226564 122703
rect 226522 121544 226578 121553
rect 226522 121479 226578 121488
rect 226522 117192 226578 117201
rect 226522 117127 226578 117136
rect 226536 116113 226564 117127
rect 226522 116104 226578 116113
rect 226522 116039 226578 116048
rect 226522 97880 226578 97889
rect 226522 97815 226578 97824
rect 226536 96937 226564 97815
rect 226522 96928 226578 96937
rect 226522 96863 226578 96872
rect 226522 92440 226578 92449
rect 226522 92375 226578 92384
rect 226536 91497 226564 92375
rect 226522 91488 226578 91497
rect 226522 91423 226578 91432
rect 226522 86864 226578 86873
rect 226522 86799 226578 86808
rect 226536 86057 226564 86799
rect 226522 86048 226578 86057
rect 226522 85983 226578 85992
rect 226522 73128 226578 73137
rect 226522 73063 226578 73072
rect 226536 72321 226564 73063
rect 226522 72312 226578 72321
rect 226522 72247 226578 72256
rect 227364 66881 227392 399910
rect 233240 399764 233292 399770
rect 233240 399706 233292 399712
rect 232044 399628 232096 399634
rect 232044 399570 232096 399576
rect 227904 398336 227956 398342
rect 227904 398278 227956 398284
rect 227812 398200 227864 398206
rect 227812 398142 227864 398148
rect 227718 398032 227774 398041
rect 227718 397967 227774 397976
rect 227442 229800 227498 229809
rect 227442 229735 227498 229744
rect 227456 200841 227484 229735
rect 227534 228440 227590 228449
rect 227534 228375 227590 228384
rect 227548 214577 227576 228375
rect 227626 227216 227682 227225
rect 227626 227151 227682 227160
rect 227534 214568 227590 214577
rect 227534 214503 227590 214512
rect 227442 200832 227498 200841
rect 227442 200767 227498 200776
rect 227640 198121 227668 227151
rect 227626 198112 227682 198121
rect 227626 198047 227682 198056
rect 227350 66872 227406 66881
rect 227350 66807 227406 66816
rect 227626 62112 227682 62121
rect 227626 62047 227682 62056
rect 227640 61441 227668 62047
rect 227626 61432 227682 61441
rect 227626 61367 227682 61376
rect 227732 58585 227760 397967
rect 227824 58993 227852 398142
rect 227810 58984 227866 58993
rect 227916 58954 227944 398278
rect 227996 398268 228048 398274
rect 227996 398210 228048 398216
rect 228008 59022 228036 398210
rect 228088 398132 228140 398138
rect 228088 398074 228140 398080
rect 227996 59016 228048 59022
rect 227996 58958 228048 58964
rect 227810 58919 227866 58928
rect 227904 58948 227956 58954
rect 227904 58890 227956 58896
rect 228100 58886 228128 398074
rect 228180 397996 228232 398002
rect 228180 397938 228232 397944
rect 228088 58880 228140 58886
rect 228088 58822 228140 58828
rect 227718 58576 227774 58585
rect 227718 58511 227774 58520
rect 228192 58342 228220 397938
rect 229100 397384 229152 397390
rect 229100 397326 229152 397332
rect 228272 396976 228324 396982
rect 228272 396918 228324 396924
rect 228284 58750 228312 396918
rect 228548 395820 228600 395826
rect 228548 395762 228600 395768
rect 228456 395752 228508 395758
rect 228456 395694 228508 395700
rect 228364 305652 228416 305658
rect 228364 305594 228416 305600
rect 228272 58744 228324 58750
rect 228272 58686 228324 58692
rect 228180 58336 228232 58342
rect 228180 58278 228232 58284
rect 228376 57866 228404 305594
rect 228468 162625 228496 395694
rect 228560 165345 228588 395762
rect 228732 319456 228784 319462
rect 228732 319398 228784 319404
rect 228640 264648 228692 264654
rect 228640 264590 228692 264596
rect 228546 165336 228602 165345
rect 228546 165271 228602 165280
rect 228454 162616 228510 162625
rect 228454 162551 228510 162560
rect 228652 77761 228680 264590
rect 228744 157185 228772 319398
rect 228824 261452 228876 261458
rect 228824 261394 228876 261400
rect 228836 209137 228864 261394
rect 228916 260636 228968 260642
rect 228916 260578 228968 260584
rect 228928 220017 228956 260578
rect 229006 242312 229062 242321
rect 229006 242247 229062 242256
rect 228914 220008 228970 220017
rect 228914 219943 228970 219952
rect 229020 211857 229048 242247
rect 229006 211848 229062 211857
rect 229006 211783 229062 211792
rect 228822 209128 228878 209137
rect 228822 209063 228878 209072
rect 228730 157176 228786 157185
rect 228730 157111 228786 157120
rect 228638 77752 228694 77761
rect 228638 77687 228694 77696
rect 229112 58478 229140 397326
rect 231952 396772 232004 396778
rect 231952 396714 232004 396720
rect 231860 396704 231912 396710
rect 231860 396646 231912 396652
rect 230572 396636 230624 396642
rect 230572 396578 230624 396584
rect 230480 396568 230532 396574
rect 230480 396510 230532 396516
rect 229192 396500 229244 396506
rect 229192 396442 229244 396448
rect 229204 58818 229232 396442
rect 229284 395548 229336 395554
rect 229284 395490 229336 395496
rect 229296 88777 229324 395490
rect 229376 264784 229428 264790
rect 229376 264726 229428 264732
rect 229282 88768 229338 88777
rect 229282 88703 229338 88712
rect 229388 59809 229416 264726
rect 229558 243536 229614 243545
rect 229558 243471 229614 243480
rect 229466 233880 229522 233889
rect 229466 233815 229522 233824
rect 229374 59800 229430 59809
rect 229374 59735 229430 59744
rect 229192 58812 229244 58818
rect 229192 58754 229244 58760
rect 229100 58472 229152 58478
rect 229100 58414 229152 58420
rect 228364 57860 228416 57866
rect 228364 57802 228416 57808
rect 229480 56914 229508 233815
rect 229572 189961 229600 243471
rect 229742 234696 229798 234705
rect 229742 234631 229798 234640
rect 229756 191865 229784 234631
rect 229742 191856 229798 191865
rect 229742 191791 229798 191800
rect 229558 189952 229614 189961
rect 229558 189887 229614 189896
rect 230492 58274 230520 396510
rect 230480 58268 230532 58274
rect 230480 58210 230532 58216
rect 230584 58138 230612 396578
rect 231124 395820 231176 395826
rect 231124 395762 231176 395768
rect 230664 264580 230716 264586
rect 230664 264522 230716 264528
rect 230676 129713 230704 264522
rect 230848 263424 230900 263430
rect 230848 263366 230900 263372
rect 230754 229936 230810 229945
rect 230754 229871 230810 229880
rect 230662 129704 230718 129713
rect 230662 129639 230718 129648
rect 230768 118833 230796 229871
rect 230860 178945 230888 263366
rect 230938 249248 230994 249257
rect 230938 249183 230994 249192
rect 230952 217297 230980 249183
rect 230938 217288 230994 217297
rect 230938 217223 230994 217232
rect 230846 178936 230902 178945
rect 230846 178871 230902 178880
rect 230754 118824 230810 118833
rect 230754 118759 230810 118768
rect 231136 105097 231164 395762
rect 231216 395548 231268 395554
rect 231216 395490 231268 395496
rect 231228 159905 231256 395490
rect 231308 260432 231360 260438
rect 231308 260374 231360 260380
rect 231320 206417 231348 260374
rect 231306 206408 231362 206417
rect 231306 206343 231362 206352
rect 231214 159896 231270 159905
rect 231214 159831 231270 159840
rect 231122 105088 231178 105097
rect 231122 105023 231178 105032
rect 230572 58132 230624 58138
rect 230572 58074 230624 58080
rect 231872 58070 231900 396646
rect 231964 58206 231992 396714
rect 232056 83201 232084 399570
rect 232504 396024 232556 396030
rect 232504 395966 232556 395972
rect 232136 378820 232188 378826
rect 232136 378762 232188 378768
rect 232042 83192 232098 83201
rect 232042 83127 232098 83136
rect 232148 80481 232176 378762
rect 232412 266076 232464 266082
rect 232412 266018 232464 266024
rect 232228 265940 232280 265946
rect 232228 265882 232280 265888
rect 232134 80472 232190 80481
rect 232134 80407 232190 80416
rect 232240 69601 232268 265882
rect 232320 264512 232372 264518
rect 232320 264454 232372 264460
rect 232332 107817 232360 264454
rect 232424 173505 232452 266018
rect 232410 173496 232466 173505
rect 232410 173431 232466 173440
rect 232318 107808 232374 107817
rect 232318 107743 232374 107752
rect 232516 73137 232544 395966
rect 233252 99657 233280 399706
rect 233424 399560 233476 399566
rect 233424 399502 233476 399508
rect 249156 399560 249208 399566
rect 249156 399502 249208 399508
rect 233332 399492 233384 399498
rect 233332 399434 233384 399440
rect 233344 102377 233372 399434
rect 233436 110673 233464 399502
rect 246304 399492 246356 399498
rect 246304 399434 246356 399440
rect 235998 398168 236054 398177
rect 235998 398103 236054 398112
rect 233976 396500 234028 396506
rect 233976 396442 234028 396448
rect 233884 395888 233936 395894
rect 233884 395830 233936 395836
rect 233516 266008 233568 266014
rect 233516 265950 233568 265956
rect 233422 110664 233478 110673
rect 233422 110599 233478 110608
rect 233330 102368 233386 102377
rect 233330 102303 233386 102312
rect 233238 99648 233294 99657
rect 233238 99583 233294 99592
rect 233528 94217 233556 265950
rect 233514 94208 233570 94217
rect 233514 94143 233570 94152
rect 233896 86873 233924 395830
rect 233988 184521 234016 396442
rect 235264 395752 235316 395758
rect 235264 395694 235316 395700
rect 234068 264512 234120 264518
rect 234068 264454 234120 264460
rect 233974 184512 234030 184521
rect 233974 184447 234030 184456
rect 234080 140729 234108 264454
rect 234066 140720 234122 140729
rect 234066 140655 234122 140664
rect 235276 125497 235304 395694
rect 235356 263424 235408 263430
rect 235356 263366 235408 263372
rect 235262 125488 235318 125497
rect 235262 125423 235318 125432
rect 233882 86864 233938 86873
rect 233882 86799 233938 86808
rect 232502 73128 232558 73137
rect 232502 73063 232558 73072
rect 232226 69592 232282 69601
rect 232226 69527 232282 69536
rect 235368 62121 235396 263366
rect 235538 232112 235594 232121
rect 235538 232047 235594 232056
rect 235446 226400 235502 226409
rect 235446 226335 235502 226344
rect 235460 99521 235488 226335
rect 235552 165753 235580 232047
rect 235630 226672 235686 226681
rect 235630 226607 235686 226616
rect 235644 218113 235672 226607
rect 235630 218104 235686 218113
rect 235630 218039 235686 218048
rect 235538 165744 235594 165753
rect 235538 165679 235594 165688
rect 235446 99512 235502 99521
rect 235446 99447 235502 99456
rect 235354 62112 235410 62121
rect 235354 62047 235410 62056
rect 232228 59628 232280 59634
rect 232228 59570 232280 59576
rect 233332 59628 233384 59634
rect 233332 59570 233384 59576
rect 232240 59514 232268 59570
rect 232240 59498 232452 59514
rect 232240 59492 232464 59498
rect 232240 59486 232412 59492
rect 232412 59434 232464 59440
rect 232228 59424 232280 59430
rect 232504 59424 232556 59430
rect 232280 59372 232504 59378
rect 232228 59366 232556 59372
rect 232240 59350 232544 59366
rect 233344 59362 233372 59570
rect 236012 59498 236040 398103
rect 236182 397352 236238 397361
rect 236182 397287 236238 397296
rect 239218 397352 239274 397361
rect 239218 397287 239274 397296
rect 241610 397352 241666 397361
rect 241610 397287 241666 397296
rect 242898 397352 242954 397361
rect 242898 397287 242954 397296
rect 244462 397352 244518 397361
rect 244462 397287 244518 397296
rect 236196 396914 236224 397287
rect 239232 397254 239260 397287
rect 238024 397248 238076 397254
rect 238024 397190 238076 397196
rect 239220 397248 239272 397254
rect 239220 397190 239272 397196
rect 236184 396908 236236 396914
rect 236184 396850 236236 396856
rect 237378 396808 237434 396817
rect 237378 396743 237434 396752
rect 236642 228032 236698 228041
rect 236642 227967 236698 227976
rect 236656 138145 236684 227967
rect 236734 226536 236790 226545
rect 236734 226471 236790 226480
rect 236748 205737 236776 226471
rect 236734 205728 236790 205737
rect 236734 205663 236790 205672
rect 236642 138136 236698 138145
rect 236642 138071 236698 138080
rect 237392 59566 237420 396743
rect 238036 59634 238064 397190
rect 241624 396846 241652 397287
rect 241612 396840 241664 396846
rect 240138 396808 240194 396817
rect 241612 396782 241664 396788
rect 240138 396743 240194 396752
rect 238116 396568 238168 396574
rect 238116 396510 238168 396516
rect 238128 195401 238156 396510
rect 238208 261452 238260 261458
rect 238208 261394 238260 261400
rect 238114 195392 238170 195401
rect 238114 195327 238170 195336
rect 238220 122777 238248 261394
rect 239402 228168 239458 228177
rect 239402 228103 239458 228112
rect 239416 178129 239444 228103
rect 239402 178120 239458 178129
rect 239402 178055 239458 178064
rect 238206 122768 238262 122777
rect 238206 122703 238262 122712
rect 240152 59906 240180 396743
rect 242256 396704 242308 396710
rect 242256 396646 242308 396652
rect 242164 396636 242216 396642
rect 242164 396578 242216 396584
rect 240876 261384 240928 261390
rect 240876 261326 240928 261332
rect 240782 227896 240838 227905
rect 240782 227831 240838 227840
rect 240796 64874 240824 227831
rect 240888 171057 240916 261326
rect 240874 171048 240930 171057
rect 240874 170983 240930 170992
rect 240704 64846 240824 64874
rect 240704 59906 240732 64846
rect 240140 59900 240192 59906
rect 240140 59842 240192 59848
rect 240692 59900 240744 59906
rect 240692 59842 240744 59848
rect 242176 59673 242204 396578
rect 242268 204241 242296 396646
rect 242912 395486 242940 397287
rect 244370 396808 244426 396817
rect 244370 396743 244426 396752
rect 242900 395480 242952 395486
rect 242900 395422 242952 395428
rect 242438 233336 242494 233345
rect 242438 233271 242494 233280
rect 242346 230344 242402 230353
rect 242346 230279 242402 230288
rect 242254 204232 242310 204241
rect 242254 204167 242310 204176
rect 242162 59664 242218 59673
rect 238024 59628 238076 59634
rect 242162 59599 242218 59608
rect 238024 59570 238076 59576
rect 237380 59560 237432 59566
rect 237380 59502 237432 59508
rect 236000 59492 236052 59498
rect 236000 59434 236052 59440
rect 233332 59356 233384 59362
rect 233332 59298 233384 59304
rect 231952 58200 232004 58206
rect 231952 58142 232004 58148
rect 231860 58064 231912 58070
rect 231860 58006 231912 58012
rect 229468 56908 229520 56914
rect 229468 56850 229520 56856
rect 226248 56840 226300 56846
rect 226248 56782 226300 56788
rect 225972 56704 226024 56710
rect 225418 56672 225474 56681
rect 225972 56646 226024 56652
rect 225418 56607 225474 56616
rect 227720 55684 227772 55690
rect 227720 55626 227772 55632
rect 226340 52896 226392 52902
rect 226340 52838 226392 52844
rect 224960 18896 225012 18902
rect 224960 18838 225012 18844
rect 224972 16574 225000 18838
rect 224972 16546 225184 16574
rect 223948 15632 224000 15638
rect 223948 15574 224000 15580
rect 223028 2848 223080 2854
rect 223028 2790 223080 2796
rect 223960 480 223988 15574
rect 225156 480 225184 16546
rect 226352 480 226380 52838
rect 227732 16574 227760 55626
rect 240140 53032 240192 53038
rect 240140 52974 240192 52980
rect 229100 52964 229152 52970
rect 229100 52906 229152 52912
rect 229112 16574 229140 52906
rect 233240 52828 233292 52834
rect 233240 52770 233292 52776
rect 233252 16574 233280 52770
rect 236000 52760 236052 52766
rect 236000 52702 236052 52708
rect 236012 16574 236040 52702
rect 238116 16584 238168 16590
rect 227732 16546 228772 16574
rect 229112 16546 229876 16574
rect 233252 16546 233464 16574
rect 236012 16546 237052 16574
rect 227536 15700 227588 15706
rect 227536 15642 227588 15648
rect 227548 480 227576 15642
rect 228744 480 228772 16546
rect 229848 480 229876 16546
rect 231032 15768 231084 15774
rect 231032 15710 231084 15716
rect 231044 480 231072 15710
rect 232228 5568 232280 5574
rect 232228 5510 232280 5516
rect 232240 480 232268 5510
rect 233436 480 233464 16546
rect 234620 15836 234672 15842
rect 234620 15778 234672 15784
rect 234632 480 234660 15778
rect 235816 5636 235868 5642
rect 235816 5578 235868 5584
rect 235828 480 235856 5578
rect 237024 480 237052 16546
rect 240152 16574 240180 52974
rect 242360 46918 242388 230279
rect 242452 71913 242480 233271
rect 242438 71904 242494 71913
rect 242438 71839 242494 71848
rect 244384 60217 244412 396743
rect 244476 395962 244504 397287
rect 245658 396808 245714 396817
rect 244924 396772 244976 396778
rect 245658 396743 245714 396752
rect 244924 396714 244976 396720
rect 244464 395956 244516 395962
rect 244464 395898 244516 395904
rect 244370 60208 244426 60217
rect 244370 60143 244426 60152
rect 244936 56817 244964 396714
rect 245672 59634 245700 396743
rect 246316 97889 246344 399434
rect 248602 397352 248658 397361
rect 248602 397287 248658 397296
rect 247130 396808 247186 396817
rect 247130 396743 247132 396752
rect 247184 396743 247186 396752
rect 247132 396714 247184 396720
rect 247682 396672 247738 396681
rect 247682 396607 247684 396616
rect 247736 396607 247738 396616
rect 247684 396578 247736 396584
rect 248616 395418 248644 397287
rect 249064 396160 249116 396166
rect 249064 396102 249116 396108
rect 248604 395412 248656 395418
rect 248604 395354 248656 395360
rect 246302 97880 246358 97889
rect 246302 97815 246358 97824
rect 245660 59628 245712 59634
rect 245660 59570 245712 59576
rect 249076 58410 249104 396102
rect 249168 92449 249196 399502
rect 265162 398168 265218 398177
rect 265162 398103 265218 398112
rect 300858 398168 300914 398177
rect 300858 398103 300914 398112
rect 315762 398168 315818 398177
rect 315762 398103 315818 398112
rect 325698 398168 325754 398177
rect 325698 398103 325754 398112
rect 250074 397352 250130 397361
rect 250074 397287 250130 397296
rect 252650 397352 252706 397361
rect 252650 397287 252706 397296
rect 253570 397352 253626 397361
rect 253570 397287 253626 397296
rect 256146 397352 256202 397361
rect 256146 397287 256202 397296
rect 260930 397352 260986 397361
rect 260930 397287 260986 397296
rect 262034 397352 262090 397361
rect 262034 397287 262090 397296
rect 263598 397352 263654 397361
rect 265176 397322 265204 398103
rect 271142 397352 271198 397361
rect 263598 397287 263654 397296
rect 265164 397316 265216 397322
rect 249890 396808 249946 396817
rect 249890 396743 249946 396752
rect 249154 92440 249210 92449
rect 249154 92375 249210 92384
rect 249904 59945 249932 396743
rect 250088 396030 250116 397287
rect 251270 396808 251326 396817
rect 251270 396743 251326 396752
rect 251178 396672 251234 396681
rect 251178 396607 251234 396616
rect 250076 396024 250128 396030
rect 250076 395966 250128 395972
rect 249890 59936 249946 59945
rect 249890 59871 249946 59880
rect 251192 59838 251220 396607
rect 251284 117201 251312 396743
rect 252664 396302 252692 397287
rect 253204 396704 253256 396710
rect 253204 396646 253256 396652
rect 252652 396296 252704 396302
rect 252652 396238 252704 396244
rect 253216 265470 253244 396646
rect 253584 395690 253612 397287
rect 254490 396808 254546 396817
rect 254490 396743 254546 396752
rect 255318 396808 255374 396817
rect 255318 396743 255374 396752
rect 254504 396710 254532 396743
rect 254492 396704 254544 396710
rect 254492 396646 254544 396652
rect 253572 395684 253624 395690
rect 253572 395626 253624 395632
rect 253204 265464 253256 265470
rect 253204 265406 253256 265412
rect 251270 117192 251326 117201
rect 251270 117127 251326 117136
rect 255332 60081 255360 396743
rect 256160 395894 256188 397287
rect 258078 396944 258134 396953
rect 258078 396879 258134 396888
rect 256698 396808 256754 396817
rect 256698 396743 256754 396752
rect 256148 395888 256200 395894
rect 256148 395830 256200 395836
rect 256712 264518 256740 396743
rect 256700 264512 256752 264518
rect 256700 264454 256752 264460
rect 255318 60072 255374 60081
rect 255318 60007 255374 60016
rect 251180 59832 251232 59838
rect 251180 59774 251232 59780
rect 249064 58404 249116 58410
rect 249064 58346 249116 58352
rect 258092 56953 258120 396879
rect 258170 396808 258226 396817
rect 258170 396743 258226 396752
rect 259458 396808 259514 396817
rect 259458 396743 259514 396752
rect 258184 268394 258212 396743
rect 258724 396296 258776 396302
rect 258724 396238 258776 396244
rect 258172 268388 258224 268394
rect 258172 268330 258224 268336
rect 258736 58614 258764 396238
rect 259472 262818 259500 396743
rect 259550 396672 259606 396681
rect 259550 396607 259606 396616
rect 259564 265810 259592 396607
rect 260944 395826 260972 397287
rect 262048 396166 262076 397287
rect 262218 396808 262274 396817
rect 262218 396743 262274 396752
rect 262036 396160 262088 396166
rect 262036 396102 262088 396108
rect 260932 395820 260984 395826
rect 260932 395762 260984 395768
rect 259552 265804 259604 265810
rect 259552 265746 259604 265752
rect 259460 262812 259512 262818
rect 259460 262754 259512 262760
rect 260102 230616 260158 230625
rect 260102 230551 260158 230560
rect 260116 126954 260144 230551
rect 260104 126948 260156 126954
rect 260104 126890 260156 126896
rect 262232 59158 262260 396743
rect 262864 396704 262916 396710
rect 262864 396646 262916 396652
rect 262876 264722 262904 396646
rect 263612 396438 263640 397287
rect 271142 397287 271198 397296
rect 273258 397352 273314 397361
rect 273258 397287 273314 397296
rect 273626 397352 273682 397361
rect 273626 397287 273682 397296
rect 274730 397352 274786 397361
rect 274730 397287 274786 397296
rect 276386 397352 276442 397361
rect 276386 397287 276442 397296
rect 278042 397352 278098 397361
rect 278042 397287 278098 397296
rect 290186 397352 290242 397361
rect 290186 397287 290242 397296
rect 293314 397352 293370 397361
rect 293314 397287 293370 397296
rect 298466 397352 298522 397361
rect 298466 397287 298522 397296
rect 300124 397316 300176 397322
rect 265164 397258 265216 397264
rect 263874 397216 263930 397225
rect 263874 397151 263930 397160
rect 263888 396710 263916 397151
rect 265254 396808 265310 396817
rect 264244 396772 264296 396778
rect 265254 396743 265256 396752
rect 264244 396714 264296 396720
rect 265308 396743 265310 396752
rect 266450 396808 266506 396817
rect 266450 396743 266506 396752
rect 267830 396808 267886 396817
rect 267830 396743 267886 396752
rect 269118 396808 269174 396817
rect 270590 396808 270646 396817
rect 269118 396743 269174 396752
rect 269764 396772 269816 396778
rect 265256 396714 265308 396720
rect 263876 396704 263928 396710
rect 263876 396646 263928 396652
rect 263600 396432 263652 396438
rect 263600 396374 263652 396380
rect 263600 396228 263652 396234
rect 263600 396170 263652 396176
rect 263612 395622 263640 396170
rect 263600 395616 263652 395622
rect 263600 395558 263652 395564
rect 262864 264716 262916 264722
rect 262864 264658 262916 264664
rect 262220 59152 262272 59158
rect 262220 59094 262272 59100
rect 264256 58682 264284 396714
rect 266358 396672 266414 396681
rect 266358 396607 266414 396616
rect 266372 261390 266400 396607
rect 266464 267034 266492 396743
rect 267738 396672 267794 396681
rect 267738 396607 267794 396616
rect 266452 267028 266504 267034
rect 266452 266970 266504 266976
rect 266360 261384 266412 261390
rect 266360 261326 266412 261332
rect 267752 59294 267780 396607
rect 267844 59906 267872 396743
rect 267832 59900 267884 59906
rect 267832 59842 267884 59848
rect 269132 59401 269160 396743
rect 270590 396743 270646 396752
rect 269764 396714 269816 396720
rect 269776 59537 269804 396714
rect 270604 261458 270632 396743
rect 271156 396506 271184 397287
rect 273272 397186 273300 397287
rect 273442 397216 273498 397225
rect 273260 397180 273312 397186
rect 273442 397151 273498 397160
rect 273260 397122 273312 397128
rect 272522 396808 272578 396817
rect 272522 396743 272524 396752
rect 272576 396743 272578 396752
rect 272524 396714 272576 396720
rect 271144 396500 271196 396506
rect 271144 396442 271196 396448
rect 273456 395758 273484 397151
rect 273640 396574 273668 397287
rect 274744 396642 274772 397287
rect 276110 396808 276166 396817
rect 276110 396743 276166 396752
rect 274732 396636 274784 396642
rect 274732 396578 274784 396584
rect 273628 396568 273680 396574
rect 273628 396510 273680 396516
rect 273444 395752 273496 395758
rect 273444 395694 273496 395700
rect 276124 265538 276152 396743
rect 276400 396234 276428 397287
rect 278056 397118 278084 397287
rect 278044 397112 278096 397118
rect 278044 397054 278096 397060
rect 277490 396808 277546 396817
rect 277490 396743 277546 396752
rect 278778 396808 278834 396817
rect 278778 396743 278834 396752
rect 280158 396808 280214 396817
rect 283562 396808 283618 396817
rect 280158 396743 280214 396752
rect 282184 396772 282236 396778
rect 276388 396228 276440 396234
rect 276388 396170 276440 396176
rect 276664 396228 276716 396234
rect 276664 396170 276716 396176
rect 276112 265532 276164 265538
rect 276112 265474 276164 265480
rect 270592 261452 270644 261458
rect 270592 261394 270644 261400
rect 269762 59528 269818 59537
rect 269762 59463 269818 59472
rect 269118 59392 269174 59401
rect 269118 59327 269174 59336
rect 267740 59288 267792 59294
rect 267740 59230 267792 59236
rect 264244 58676 264296 58682
rect 264244 58618 264296 58624
rect 258724 58608 258776 58614
rect 258724 58550 258776 58556
rect 258078 56944 258134 56953
rect 258078 56879 258134 56888
rect 244922 56808 244978 56817
rect 244922 56743 244978 56752
rect 276676 56642 276704 396170
rect 277504 56982 277532 396743
rect 278792 265742 278820 396743
rect 278780 265736 278832 265742
rect 278780 265678 278832 265684
rect 280172 264450 280200 396743
rect 283562 396743 283564 396752
rect 282184 396714 282236 396720
rect 283616 396743 283618 396752
rect 285954 396808 286010 396817
rect 285954 396743 286010 396752
rect 287058 396808 287114 396817
rect 287058 396743 287114 396752
rect 283564 396714 283616 396720
rect 280160 264444 280212 264450
rect 280160 264386 280212 264392
rect 282196 260574 282224 396714
rect 285968 396710 285996 396743
rect 284944 396704 284996 396710
rect 284944 396646 284996 396652
rect 285956 396704 286008 396710
rect 285956 396646 286008 396652
rect 284956 262206 284984 396646
rect 287072 263498 287100 396743
rect 290200 395350 290228 397287
rect 291844 396160 291896 396166
rect 291844 396102 291896 396108
rect 290188 395344 290240 395350
rect 290188 395286 290240 395292
rect 291856 263566 291884 396102
rect 293328 395554 293356 397287
rect 295338 396808 295394 396817
rect 295338 396743 295394 396752
rect 293316 395548 293368 395554
rect 293316 395490 293368 395496
rect 295352 264382 295380 396743
rect 298480 396234 298508 397287
rect 300124 397258 300176 397264
rect 298468 396228 298520 396234
rect 298468 396170 298520 396176
rect 295340 264376 295392 264382
rect 295340 264318 295392 264324
rect 291844 263560 291896 263566
rect 291844 263502 291896 263508
rect 287060 263492 287112 263498
rect 287060 263434 287112 263440
rect 284944 262200 284996 262206
rect 284944 262142 284996 262148
rect 282184 260568 282236 260574
rect 282184 260510 282236 260516
rect 281998 247072 282054 247081
rect 281998 247007 282054 247016
rect 282012 245614 282040 247007
rect 282000 245608 282052 245614
rect 282000 245550 282052 245556
rect 300136 57186 300164 397258
rect 300872 396166 300900 398103
rect 308586 397352 308642 397361
rect 308586 397287 308588 397296
rect 308640 397287 308642 397296
rect 310978 397352 311034 397361
rect 310978 397287 311034 397296
rect 313370 397352 313426 397361
rect 313370 397287 313426 397296
rect 308588 397258 308640 397264
rect 302238 396808 302294 396817
rect 302238 396743 302294 396752
rect 304998 396808 305054 396817
rect 304998 396743 305054 396752
rect 300860 396160 300912 396166
rect 300860 396102 300912 396108
rect 300124 57180 300176 57186
rect 300124 57122 300176 57128
rect 302252 57050 302280 396743
rect 304264 396092 304316 396098
rect 304264 396034 304316 396040
rect 304276 260506 304304 396034
rect 305012 264314 305040 396743
rect 307024 396704 307076 396710
rect 307024 396646 307076 396652
rect 305000 264308 305052 264314
rect 305000 264250 305052 264256
rect 307036 262138 307064 396646
rect 310992 396370 311020 397287
rect 310980 396364 311032 396370
rect 310980 396306 311032 396312
rect 313384 396098 313412 397287
rect 315776 396710 315804 398103
rect 317418 396808 317474 396817
rect 317418 396743 317474 396752
rect 320178 396808 320234 396817
rect 320178 396743 320234 396752
rect 322938 396808 322994 396817
rect 322938 396743 322994 396752
rect 315764 396704 315816 396710
rect 315764 396646 315816 396652
rect 313372 396092 313424 396098
rect 313372 396034 313424 396040
rect 307024 262132 307076 262138
rect 307024 262074 307076 262080
rect 317432 262070 317460 396743
rect 317420 262064 317472 262070
rect 317420 262006 317472 262012
rect 304264 260500 304316 260506
rect 304264 260442 304316 260448
rect 320192 260438 320220 396743
rect 320180 260432 320232 260438
rect 320180 260374 320232 260380
rect 322952 59430 322980 396743
rect 325712 265674 325740 398103
rect 342258 397352 342314 397361
rect 342258 397287 342314 397296
rect 342272 396302 342300 397287
rect 342350 396808 342406 396817
rect 342350 396743 342406 396752
rect 342260 396296 342312 396302
rect 342260 396238 342312 396244
rect 342364 301510 342392 396743
rect 342352 301504 342404 301510
rect 342352 301446 342404 301452
rect 325700 265668 325752 265674
rect 325700 265610 325752 265616
rect 322940 59424 322992 59430
rect 322940 59366 322992 59372
rect 356532 58721 356560 485823
rect 358818 478952 358874 478961
rect 358818 478887 358874 478896
rect 358084 456816 358136 456822
rect 358084 456758 358136 456764
rect 357438 414352 357494 414361
rect 357438 414287 357494 414296
rect 357452 237969 357480 414287
rect 357530 413128 357586 413137
rect 357530 413063 357586 413072
rect 357544 399702 357572 413063
rect 357532 399696 357584 399702
rect 357532 399638 357584 399644
rect 358096 260234 358124 456758
rect 358832 263430 358860 478887
rect 358910 418840 358966 418849
rect 358910 418775 358966 418784
rect 358820 263424 358872 263430
rect 358820 263366 358872 263372
rect 358084 260228 358136 260234
rect 358084 260170 358136 260176
rect 358924 260166 358952 418775
rect 359002 417208 359058 417217
rect 359002 417143 359058 417152
rect 359016 399566 359044 417143
rect 359094 415848 359150 415857
rect 359094 415783 359150 415792
rect 359004 399560 359056 399566
rect 359004 399502 359056 399508
rect 359108 399498 359136 415783
rect 359096 399492 359148 399498
rect 359096 399434 359148 399440
rect 360856 260370 360884 510614
rect 360844 260364 360896 260370
rect 360844 260306 360896 260312
rect 363616 260302 363644 563042
rect 367756 261934 367784 616830
rect 370516 262002 370544 700402
rect 382924 700392 382976 700398
rect 382924 700334 382976 700340
rect 381544 696992 381596 696998
rect 381544 696934 381596 696940
rect 377404 643136 377456 643142
rect 377404 643078 377456 643084
rect 376024 590708 376076 590714
rect 376024 590650 376076 590656
rect 374644 484424 374696 484430
rect 374644 484366 374696 484372
rect 371884 404388 371936 404394
rect 371884 404330 371936 404336
rect 370504 261996 370556 262002
rect 370504 261938 370556 261944
rect 367744 261928 367796 261934
rect 367744 261870 367796 261876
rect 371896 261594 371924 404330
rect 374656 261662 374684 484366
rect 376036 300150 376064 590650
rect 376024 300144 376076 300150
rect 376024 300086 376076 300092
rect 377416 261866 377444 643078
rect 378784 536852 378836 536858
rect 378784 536794 378836 536800
rect 378796 298790 378824 536794
rect 378784 298784 378836 298790
rect 378784 298726 378836 298732
rect 377404 261860 377456 261866
rect 377404 261802 377456 261808
rect 381556 261730 381584 696934
rect 382936 261798 382964 700334
rect 385696 263294 385724 700538
rect 397472 700534 397500 703520
rect 388444 700528 388496 700534
rect 388444 700470 388496 700476
rect 397460 700528 397512 700534
rect 397460 700470 397512 700476
rect 400864 700528 400916 700534
rect 400864 700470 400916 700476
rect 388456 263362 388484 700470
rect 399484 683188 399536 683194
rect 399484 683130 399536 683136
rect 396724 630692 396776 630698
rect 396724 630634 396776 630640
rect 395344 576904 395396 576910
rect 395344 576846 395396 576852
rect 393964 524476 394016 524482
rect 393964 524418 394016 524424
rect 392584 470620 392636 470626
rect 392584 470562 392636 470568
rect 389824 430636 389876 430642
rect 389824 430578 389876 430584
rect 388444 263356 388496 263362
rect 388444 263298 388496 263304
rect 385684 263288 385736 263294
rect 385684 263230 385736 263236
rect 389836 262886 389864 430578
rect 392596 262954 392624 470562
rect 393976 263022 394004 524418
rect 395356 263090 395384 576846
rect 396736 263226 396764 630634
rect 396724 263220 396776 263226
rect 396724 263162 396776 263168
rect 399496 263158 399524 683130
rect 399484 263152 399536 263158
rect 399484 263094 399536 263100
rect 395344 263084 395396 263090
rect 395344 263026 395396 263032
rect 393964 263016 394016 263022
rect 393964 262958 394016 262964
rect 392584 262948 392636 262954
rect 392584 262890 392636 262896
rect 389824 262880 389876 262886
rect 389824 262822 389876 262828
rect 382924 261792 382976 261798
rect 382924 261734 382976 261740
rect 381544 261724 381596 261730
rect 381544 261666 381596 261672
rect 374644 261656 374696 261662
rect 374644 261598 374696 261604
rect 371884 261588 371936 261594
rect 371884 261530 371936 261536
rect 400876 261526 400904 700470
rect 412652 294710 412680 703582
rect 413480 703474 413508 703582
rect 413622 703520 413734 704960
rect 429212 703582 429700 703610
rect 413664 703474 413692 703520
rect 413480 703446 413692 703474
rect 412640 294704 412692 294710
rect 412640 294646 412692 294652
rect 429212 284986 429240 703582
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 462332 700602 462360 703520
rect 462320 700596 462372 700602
rect 462320 700538 462372 700544
rect 478524 700534 478552 703520
rect 478512 700528 478564 700534
rect 478512 700470 478564 700476
rect 494808 700466 494836 703520
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 527192 700398 527220 703520
rect 543476 702434 543504 703520
rect 542372 702406 543504 702434
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 542372 294642 542400 702406
rect 559668 700330 559696 703520
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 697232 580226 697241
rect 580170 697167 580226 697176
rect 580184 696998 580212 697167
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 683904 580226 683913
rect 580170 683839 580226 683848
rect 580184 683194 580212 683839
rect 580172 683188 580224 683194
rect 580172 683130 580224 683136
rect 580172 670744 580224 670750
rect 580170 670712 580172 670721
rect 580224 670712 580226 670721
rect 580170 670647 580226 670656
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580184 643142 580212 643991
rect 580172 643136 580224 643142
rect 580172 643078 580224 643084
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580184 630698 580212 630799
rect 580172 630692 580224 630698
rect 580172 630634 580224 630640
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580184 616894 580212 617471
rect 580172 616888 580224 616894
rect 580172 616830 580224 616836
rect 579802 591016 579858 591025
rect 579802 590951 579858 590960
rect 579816 590714 579844 590951
rect 579804 590708 579856 590714
rect 579804 590650 579856 590656
rect 580170 577688 580226 577697
rect 580170 577623 580226 577632
rect 580184 576910 580212 577623
rect 580172 576904 580224 576910
rect 580172 576846 580224 576852
rect 579802 564360 579858 564369
rect 579802 564295 579858 564304
rect 579816 563106 579844 564295
rect 579804 563100 579856 563106
rect 579804 563042 579856 563048
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580184 536858 580212 537775
rect 580172 536852 580224 536858
rect 580172 536794 580224 536800
rect 580170 524512 580226 524521
rect 580170 524447 580172 524456
rect 580224 524447 580226 524456
rect 580172 524418 580224 524424
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 580184 510678 580212 511255
rect 580172 510672 580224 510678
rect 580172 510614 580224 510620
rect 580170 484664 580226 484673
rect 580170 484599 580226 484608
rect 580184 484430 580212 484599
rect 580172 484424 580224 484430
rect 580172 484366 580224 484372
rect 579986 471472 580042 471481
rect 579986 471407 580042 471416
rect 580000 470626 580028 471407
rect 579988 470620 580040 470626
rect 579988 470562 580040 470568
rect 580170 458144 580226 458153
rect 580170 458079 580226 458088
rect 580184 456822 580212 458079
rect 580172 456816 580224 456822
rect 580172 456758 580224 456764
rect 580170 431624 580226 431633
rect 580170 431559 580226 431568
rect 580184 430642 580212 431559
rect 580172 430636 580224 430642
rect 580172 430578 580224 430584
rect 580262 418296 580318 418305
rect 580262 418231 580318 418240
rect 580170 404968 580226 404977
rect 580170 404903 580226 404912
rect 580184 404394 580212 404903
rect 580172 404388 580224 404394
rect 580172 404330 580224 404336
rect 580170 378448 580226 378457
rect 580170 378383 580226 378392
rect 580184 378214 580212 378383
rect 580172 378208 580224 378214
rect 580172 378150 580224 378156
rect 579618 365120 579674 365129
rect 579618 365055 579674 365064
rect 579632 364410 579660 365055
rect 579620 364404 579672 364410
rect 579620 364346 579672 364352
rect 580172 351960 580224 351966
rect 580170 351928 580172 351937
rect 580224 351928 580226 351937
rect 580170 351863 580226 351872
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580184 324358 580212 325207
rect 580172 324352 580224 324358
rect 580172 324294 580224 324300
rect 579986 312080 580042 312089
rect 579986 312015 580042 312024
rect 580000 311914 580028 312015
rect 579988 311908 580040 311914
rect 579988 311850 580040 311856
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 580184 298178 580212 298687
rect 580172 298172 580224 298178
rect 580172 298114 580224 298120
rect 542360 294636 542412 294642
rect 542360 294578 542412 294584
rect 429200 284980 429252 284986
rect 429200 284922 429252 284928
rect 580170 272232 580226 272241
rect 580170 272167 580226 272176
rect 580184 271930 580212 272167
rect 580172 271924 580224 271930
rect 580172 271866 580224 271872
rect 580276 264246 580304 418231
rect 580264 264240 580316 264246
rect 580264 264182 580316 264188
rect 400864 261520 400916 261526
rect 400864 261462 400916 261468
rect 363604 260296 363656 260302
rect 363604 260238 363656 260244
rect 358912 260160 358964 260166
rect 358912 260102 358964 260108
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 357438 237960 357494 237969
rect 357438 237895 357494 237904
rect 396722 227760 396778 227769
rect 396722 227695 396778 227704
rect 396736 153202 396764 227695
rect 580262 226944 580318 226953
rect 580262 226879 580318 226888
rect 396724 153196 396776 153202
rect 396724 153138 396776 153144
rect 579620 153196 579672 153202
rect 579620 153138 579672 153144
rect 579632 152697 579660 153138
rect 579618 152688 579674 152697
rect 579618 152623 579674 152632
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580172 59968 580224 59974
rect 580172 59910 580224 59916
rect 580184 59673 580212 59910
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 356518 58712 356574 58721
rect 356518 58647 356574 58656
rect 347042 57352 347098 57361
rect 347042 57287 347098 57296
rect 302240 57044 302292 57050
rect 302240 56986 302292 56992
rect 277492 56976 277544 56982
rect 277492 56918 277544 56924
rect 276664 56636 276716 56642
rect 276664 56578 276716 56584
rect 313280 55208 313332 55214
rect 313280 55150 313332 55156
rect 309140 54460 309192 54466
rect 309140 54402 309192 54408
rect 302240 54392 302292 54398
rect 302240 54334 302292 54340
rect 299480 54324 299532 54330
rect 299480 54266 299532 54272
rect 251180 52420 251232 52426
rect 251180 52362 251232 52368
rect 247040 51672 247092 51678
rect 247040 51614 247092 51620
rect 242348 46912 242400 46918
rect 242348 46854 242400 46860
rect 242900 24132 242952 24138
rect 242900 24074 242952 24080
rect 240152 16546 240548 16574
rect 238116 16526 238168 16532
rect 238128 480 238156 16526
rect 239312 5704 239364 5710
rect 239312 5646 239364 5652
rect 239324 480 239352 5646
rect 240520 480 240548 16546
rect 241704 16516 241756 16522
rect 241704 16458 241756 16464
rect 241716 480 241744 16458
rect 242912 2786 242940 24074
rect 247052 16574 247080 51614
rect 247052 16546 247632 16574
rect 245200 16448 245252 16454
rect 245200 16390 245252 16396
rect 242992 5772 243044 5778
rect 242992 5714 243044 5720
rect 242900 2780 242952 2786
rect 242900 2722 242952 2728
rect 243004 2666 243032 5714
rect 244096 2780 244148 2786
rect 244096 2722 244148 2728
rect 242912 2638 243032 2666
rect 242912 480 242940 2638
rect 244108 480 244136 2722
rect 245212 480 245240 16390
rect 246396 5840 246448 5846
rect 246396 5782 246448 5788
rect 246408 480 246436 5782
rect 247604 480 247632 16546
rect 248788 16380 248840 16386
rect 248788 16322 248840 16328
rect 248800 480 248828 16322
rect 249984 5908 250036 5914
rect 249984 5850 250036 5856
rect 249996 480 250024 5850
rect 251192 480 251220 52362
rect 253940 52352 253992 52358
rect 253940 52294 253992 52300
rect 253952 16574 253980 52294
rect 280160 50244 280212 50250
rect 280160 50186 280212 50192
rect 269120 17944 269172 17950
rect 269120 17886 269172 17892
rect 266360 17196 266412 17202
rect 266360 17138 266412 17144
rect 262220 17128 262272 17134
rect 262220 17070 262272 17076
rect 262232 16574 262260 17070
rect 266372 16574 266400 17138
rect 269132 16574 269160 17886
rect 273260 17876 273312 17882
rect 273260 17818 273312 17824
rect 273272 16574 273300 17818
rect 276020 17808 276072 17814
rect 276020 17750 276072 17756
rect 253952 16546 254716 16574
rect 262232 16546 262996 16574
rect 266372 16546 266584 16574
rect 269132 16546 270080 16574
rect 273272 16546 273668 16574
rect 252376 16312 252428 16318
rect 252376 16254 252428 16260
rect 252388 480 252416 16254
rect 253480 5976 253532 5982
rect 253480 5918 253532 5924
rect 253492 480 253520 5918
rect 254688 480 254716 16546
rect 255872 16244 255924 16250
rect 255872 16186 255924 16192
rect 255884 480 255912 16186
rect 259460 16176 259512 16182
rect 259460 16118 259512 16124
rect 258264 11212 258316 11218
rect 258264 11154 258316 11160
rect 257068 6044 257120 6050
rect 257068 5986 257120 5992
rect 257080 480 257108 5986
rect 258276 480 258304 11154
rect 259472 480 259500 16118
rect 261760 11280 261812 11286
rect 261760 11222 261812 11228
rect 260656 6112 260708 6118
rect 260656 6054 260708 6060
rect 260668 480 260696 6054
rect 261772 480 261800 11222
rect 262968 480 262996 16546
rect 265348 11348 265400 11354
rect 265348 11290 265400 11296
rect 264152 6860 264204 6866
rect 264152 6802 264204 6808
rect 264164 480 264192 6802
rect 265360 480 265388 11290
rect 266556 480 266584 16546
rect 268844 11416 268896 11422
rect 268844 11358 268896 11364
rect 267740 6792 267792 6798
rect 267740 6734 267792 6740
rect 267752 480 267780 6734
rect 268856 480 268884 11358
rect 270052 480 270080 16546
rect 271236 6724 271288 6730
rect 271236 6666 271288 6672
rect 271248 480 271276 6666
rect 272432 3120 272484 3126
rect 272432 3062 272484 3068
rect 272444 480 272472 3062
rect 273640 480 273668 16546
rect 274824 6656 274876 6662
rect 274824 6598 274876 6604
rect 274836 480 274864 6598
rect 276032 5574 276060 17750
rect 280172 16574 280200 50186
rect 291200 49360 291252 49366
rect 291200 49302 291252 49308
rect 287060 17740 287112 17746
rect 287060 17682 287112 17688
rect 287072 16574 287100 17682
rect 291212 16574 291240 49302
rect 298100 17604 298152 17610
rect 298100 17546 298152 17552
rect 298112 16574 298140 17546
rect 280172 16546 280752 16574
rect 287072 16546 287836 16574
rect 291212 16546 291424 16574
rect 298112 16546 298508 16574
rect 279516 11552 279568 11558
rect 279516 11494 279568 11500
rect 276112 11484 276164 11490
rect 276112 11426 276164 11432
rect 276020 5568 276072 5574
rect 276020 5510 276072 5516
rect 276124 3482 276152 11426
rect 278320 6588 278372 6594
rect 278320 6530 278372 6536
rect 277124 5568 277176 5574
rect 277124 5510 277176 5516
rect 276032 3454 276152 3482
rect 276032 480 276060 3454
rect 277136 480 277164 5510
rect 278332 480 278360 6530
rect 279528 480 279556 11494
rect 280724 480 280752 16546
rect 286600 11620 286652 11626
rect 286600 11562 286652 11568
rect 281908 6520 281960 6526
rect 281908 6462 281960 6468
rect 281920 480 281948 6462
rect 285404 6452 285456 6458
rect 285404 6394 285456 6400
rect 284300 3188 284352 3194
rect 284300 3130 284352 3136
rect 283104 2848 283156 2854
rect 283104 2790 283156 2796
rect 283116 480 283144 2790
rect 284312 480 284340 3130
rect 285416 480 285444 6394
rect 286612 480 286640 11562
rect 287808 480 287836 16546
rect 290188 11688 290240 11694
rect 290188 11630 290240 11636
rect 288992 6384 289044 6390
rect 288992 6326 289044 6332
rect 289004 480 289032 6326
rect 290200 480 290228 11630
rect 291396 480 291424 16546
rect 293684 12436 293736 12442
rect 293684 12378 293736 12384
rect 292580 6316 292632 6322
rect 292580 6258 292632 6264
rect 292592 480 292620 6258
rect 293696 480 293724 12378
rect 297272 12368 297324 12374
rect 297272 12310 297324 12316
rect 296076 6248 296128 6254
rect 296076 6190 296128 6196
rect 294880 2916 294932 2922
rect 294880 2858 294932 2864
rect 294892 480 294920 2858
rect 296088 480 296116 6190
rect 297284 480 297312 12310
rect 298480 480 298508 16546
rect 299492 3482 299520 54266
rect 300860 17536 300912 17542
rect 300860 17478 300912 17484
rect 300872 16574 300900 17478
rect 302252 16574 302280 54334
rect 307760 17468 307812 17474
rect 307760 17410 307812 17416
rect 300872 16546 302004 16574
rect 302252 16546 303200 16574
rect 299572 12300 299624 12306
rect 299572 12242 299624 12248
rect 299584 5574 299612 12242
rect 299572 5568 299624 5574
rect 299572 5510 299624 5516
rect 300768 5568 300820 5574
rect 300768 5510 300820 5516
rect 299492 3454 299704 3482
rect 299676 480 299704 3454
rect 300780 480 300808 5510
rect 301976 480 302004 16546
rect 303172 480 303200 16546
rect 304356 12232 304408 12238
rect 304356 12174 304408 12180
rect 304368 480 304396 12174
rect 307772 3398 307800 17410
rect 309152 16574 309180 54402
rect 311900 49156 311952 49162
rect 311900 49098 311952 49104
rect 311912 16574 311940 49098
rect 313292 16574 313320 55150
rect 316040 55140 316092 55146
rect 316040 55082 316092 55088
rect 309152 16546 310284 16574
rect 311912 16546 312676 16574
rect 313292 16546 313872 16574
rect 307944 12164 307996 12170
rect 307944 12106 307996 12112
rect 306748 3392 306800 3398
rect 306748 3334 306800 3340
rect 307760 3392 307812 3398
rect 307760 3334 307812 3340
rect 305552 3324 305604 3330
rect 305552 3266 305604 3272
rect 305564 480 305592 3266
rect 306760 480 306788 3334
rect 307956 480 307984 12106
rect 309048 3392 309100 3398
rect 309048 3334 309100 3340
rect 309060 480 309088 3334
rect 310256 480 310284 16546
rect 311440 12096 311492 12102
rect 311440 12038 311492 12044
rect 311452 480 311480 12038
rect 312648 480 312676 16546
rect 313844 480 313872 16546
rect 315028 12028 315080 12034
rect 315028 11970 315080 11976
rect 315040 480 315068 11970
rect 316052 3398 316080 55082
rect 320180 55072 320232 55078
rect 320180 55014 320232 55020
rect 318800 18828 318852 18834
rect 318800 18770 318852 18776
rect 316132 17400 316184 17406
rect 316132 17342 316184 17348
rect 316144 16574 316172 17342
rect 318812 16574 318840 18770
rect 320192 16574 320220 55014
rect 324320 55004 324372 55010
rect 324320 54946 324372 54952
rect 322940 49224 322992 49230
rect 322940 49166 322992 49172
rect 322952 16574 322980 49166
rect 324332 16574 324360 54946
rect 327080 54936 327132 54942
rect 327080 54878 327132 54884
rect 325700 18760 325752 18766
rect 325700 18702 325752 18708
rect 325712 16574 325740 18702
rect 327092 16574 327120 54878
rect 335360 52284 335412 52290
rect 335360 52226 335412 52232
rect 329840 49292 329892 49298
rect 329840 49234 329892 49240
rect 329852 16574 329880 49234
rect 332600 17332 332652 17338
rect 332600 17274 332652 17280
rect 316144 16546 316264 16574
rect 318812 16546 319760 16574
rect 320192 16546 320956 16574
rect 322952 16546 323348 16574
rect 324332 16546 324452 16574
rect 325712 16546 326844 16574
rect 327092 16546 328040 16574
rect 329852 16546 330432 16574
rect 316040 3392 316092 3398
rect 316040 3334 316092 3340
rect 316236 480 316264 16546
rect 318524 11960 318576 11966
rect 318524 11902 318576 11908
rect 317328 3392 317380 3398
rect 317328 3334 317380 3340
rect 317340 480 317368 3334
rect 318536 480 318564 11902
rect 319732 480 319760 16546
rect 320928 480 320956 16546
rect 322112 11892 322164 11898
rect 322112 11834 322164 11840
rect 322124 480 322152 11834
rect 323320 480 323348 16546
rect 324424 480 324452 16546
rect 325608 11824 325660 11830
rect 325608 11766 325660 11772
rect 325620 480 325648 11766
rect 326816 480 326844 16546
rect 328012 480 328040 16546
rect 329196 11756 329248 11762
rect 329196 11698 329248 11704
rect 329208 480 329236 11698
rect 330404 480 330432 16546
rect 331588 7064 331640 7070
rect 331588 7006 331640 7012
rect 331600 480 331628 7006
rect 332612 3398 332640 17274
rect 332692 17264 332744 17270
rect 332692 17206 332744 17212
rect 332600 3392 332652 3398
rect 332600 3334 332652 3340
rect 332704 480 332732 17206
rect 335372 16574 335400 52226
rect 339500 52216 339552 52222
rect 339500 52158 339552 52164
rect 339512 16574 339540 52158
rect 342260 52148 342312 52154
rect 342260 52090 342312 52096
rect 340880 49088 340932 49094
rect 340880 49030 340932 49036
rect 340892 16574 340920 49030
rect 342272 16574 342300 52090
rect 346400 52080 346452 52086
rect 346400 52022 346452 52028
rect 343640 17672 343692 17678
rect 343640 17614 343692 17620
rect 343652 16574 343680 17614
rect 346412 16574 346440 52022
rect 335372 16546 336320 16574
rect 339512 16546 339908 16574
rect 340892 16546 341012 16574
rect 342272 16546 343404 16574
rect 343652 16546 344600 16574
rect 346412 16546 346992 16574
rect 335084 7132 335136 7138
rect 335084 7074 335136 7080
rect 333888 3392 333940 3398
rect 333888 3334 333940 3340
rect 333900 480 333928 3334
rect 335096 480 335124 7074
rect 336292 480 336320 16546
rect 338672 7200 338724 7206
rect 338672 7142 338724 7148
rect 337476 2984 337528 2990
rect 337476 2926 337528 2932
rect 337488 480 337516 2926
rect 338684 480 338712 7142
rect 339880 480 339908 16546
rect 340984 480 341012 16546
rect 342168 7268 342220 7274
rect 342168 7210 342220 7216
rect 342180 480 342208 7210
rect 343376 480 343404 16546
rect 344572 480 344600 16546
rect 345756 7336 345808 7342
rect 345756 7278 345808 7284
rect 345768 480 345796 7278
rect 346964 480 346992 16546
rect 347056 3398 347084 57287
rect 401600 57248 401652 57254
rect 401600 57190 401652 57196
rect 429842 57216 429898 57225
rect 357532 52012 357584 52018
rect 357532 51954 357584 51960
rect 356336 7472 356388 7478
rect 356336 7414 356388 7420
rect 352840 7404 352892 7410
rect 352840 7346 352892 7352
rect 348056 4004 348108 4010
rect 348056 3946 348108 3952
rect 347044 3392 347096 3398
rect 347044 3334 347096 3340
rect 348068 480 348096 3946
rect 351644 3936 351696 3942
rect 351644 3878 351696 3884
rect 349252 3392 349304 3398
rect 349252 3334 349304 3340
rect 349264 480 349292 3334
rect 350448 3052 350500 3058
rect 350448 2994 350500 3000
rect 350460 480 350488 2994
rect 351656 480 351684 3878
rect 352852 480 352880 7346
rect 354036 3868 354088 3874
rect 354036 3810 354088 3816
rect 354048 480 354076 3810
rect 355232 3800 355284 3806
rect 355232 3742 355284 3748
rect 355244 480 355272 3742
rect 356348 480 356376 7414
rect 357544 480 357572 51954
rect 364340 51944 364392 51950
rect 364340 51886 364392 51892
rect 360200 50312 360252 50318
rect 360200 50254 360252 50260
rect 360212 16574 360240 50254
rect 361580 18692 361632 18698
rect 361580 18634 361632 18640
rect 361592 16574 361620 18634
rect 364352 16574 364380 51886
rect 401612 16574 401640 57190
rect 429842 57151 429898 57160
rect 417424 55752 417476 55758
rect 417424 55694 417476 55700
rect 405740 54868 405792 54874
rect 405740 54810 405792 54816
rect 405752 16574 405780 54810
rect 412640 54800 412692 54806
rect 412640 54742 412692 54748
rect 407764 53780 407816 53786
rect 407764 53722 407816 53728
rect 360212 16546 361160 16574
rect 361592 16546 362356 16574
rect 364352 16546 364656 16574
rect 401612 16546 402560 16574
rect 405752 16546 406056 16574
rect 359924 7540 359976 7546
rect 359924 7482 359976 7488
rect 358728 3732 358780 3738
rect 358728 3674 358780 3680
rect 358740 480 358768 3674
rect 359936 480 359964 7482
rect 361132 480 361160 16546
rect 362328 480 362356 16546
rect 363512 8288 363564 8294
rect 363512 8230 363564 8236
rect 363524 480 363552 8230
rect 364628 480 364656 16546
rect 396540 13796 396592 13802
rect 396540 13738 396592 13744
rect 393044 13048 393096 13054
rect 393044 12990 393096 12996
rect 389456 12980 389508 12986
rect 389456 12922 389508 12928
rect 385960 12912 386012 12918
rect 385960 12854 386012 12860
rect 382372 12844 382424 12850
rect 382372 12786 382424 12792
rect 378876 12776 378928 12782
rect 378876 12718 378928 12724
rect 374000 12708 374052 12714
rect 374000 12650 374052 12656
rect 368204 12640 368256 12646
rect 368204 12582 368256 12588
rect 367008 8220 367060 8226
rect 367008 8162 367060 8168
rect 365812 3664 365864 3670
rect 365812 3606 365864 3612
rect 365824 480 365852 3606
rect 367020 480 367048 8162
rect 368216 480 368244 12582
rect 370596 8152 370648 8158
rect 370596 8094 370648 8100
rect 369400 6180 369452 6186
rect 369400 6122 369452 6128
rect 368478 5808 368534 5817
rect 368478 5743 368534 5752
rect 368492 2990 368520 5743
rect 368480 2984 368532 2990
rect 368480 2926 368532 2932
rect 369412 480 369440 6122
rect 370608 480 370636 8094
rect 374012 3602 374040 12650
rect 374092 8084 374144 8090
rect 374092 8026 374144 8032
rect 372896 3596 372948 3602
rect 372896 3538 372948 3544
rect 374000 3596 374052 3602
rect 374000 3538 374052 3544
rect 371700 2984 371752 2990
rect 371700 2926 371752 2932
rect 371712 480 371740 2926
rect 372908 480 372936 3538
rect 374104 480 374132 8026
rect 377680 8016 377732 8022
rect 377680 7958 377732 7964
rect 375288 3596 375340 3602
rect 375288 3538 375340 3544
rect 375300 480 375328 3538
rect 376484 3528 376536 3534
rect 376484 3470 376536 3476
rect 376496 480 376524 3470
rect 377692 480 377720 7958
rect 378888 480 378916 12718
rect 381176 7948 381228 7954
rect 381176 7890 381228 7896
rect 379980 3460 380032 3466
rect 379980 3402 380032 3408
rect 379992 480 380020 3402
rect 381188 480 381216 7890
rect 382384 480 382412 12786
rect 384764 7880 384816 7886
rect 384764 7822 384816 7828
rect 383566 5944 383622 5953
rect 383566 5879 383622 5888
rect 383580 480 383608 5879
rect 384776 480 384804 7822
rect 385972 480 386000 12854
rect 388260 7812 388312 7818
rect 388260 7754 388312 7760
rect 387156 3256 387208 3262
rect 387156 3198 387208 3204
rect 387168 480 387196 3198
rect 388272 480 388300 7754
rect 389468 480 389496 12922
rect 391848 7744 391900 7750
rect 391848 7686 391900 7692
rect 390652 4140 390704 4146
rect 390652 4082 390704 4088
rect 390664 480 390692 4082
rect 391860 480 391888 7686
rect 393056 480 393084 12990
rect 395344 7676 395396 7682
rect 395344 7618 395396 7624
rect 394238 6080 394294 6089
rect 394238 6015 394294 6024
rect 394252 480 394280 6015
rect 395356 480 395384 7618
rect 396552 480 396580 13738
rect 398840 13728 398892 13734
rect 398840 13670 398892 13676
rect 397734 6896 397790 6905
rect 397734 6831 397790 6840
rect 397748 480 397776 6831
rect 398852 3534 398880 13670
rect 398932 7608 398984 7614
rect 398932 7550 398984 7556
rect 398840 3528 398892 3534
rect 398840 3470 398892 3476
rect 398944 480 398972 7550
rect 400128 3528 400180 3534
rect 400128 3470 400180 3476
rect 400140 480 400168 3470
rect 401324 2168 401376 2174
rect 401324 2110 401376 2116
rect 401336 480 401364 2110
rect 402532 480 402560 16546
rect 403624 13660 403676 13666
rect 403624 13602 403676 13608
rect 403636 480 403664 13602
rect 404820 4072 404872 4078
rect 404820 4014 404872 4020
rect 404832 480 404860 4014
rect 406028 480 406056 16546
rect 407212 13592 407264 13598
rect 407212 13534 407264 13540
rect 407224 480 407252 13534
rect 407776 3058 407804 53722
rect 412652 16574 412680 54742
rect 414664 53712 414716 53718
rect 414664 53654 414716 53660
rect 412652 16546 413140 16574
rect 410800 13524 410852 13530
rect 410800 13466 410852 13472
rect 408406 3904 408462 3913
rect 408406 3839 408462 3848
rect 407764 3052 407816 3058
rect 407764 2994 407816 3000
rect 408420 480 408448 3839
rect 409604 3052 409656 3058
rect 409604 2994 409656 3000
rect 409616 480 409644 2994
rect 410812 480 410840 13466
rect 411902 3088 411958 3097
rect 411902 3023 411958 3032
rect 411916 480 411944 3023
rect 413112 480 413140 16546
rect 414296 13456 414348 13462
rect 414296 13398 414348 13404
rect 414308 480 414336 13398
rect 414676 3534 414704 53654
rect 417436 16574 417464 55694
rect 421564 53644 421616 53650
rect 421564 53586 421616 53592
rect 417436 16546 417556 16574
rect 417424 13388 417476 13394
rect 417424 13330 417476 13336
rect 415490 3768 415546 3777
rect 415490 3703 415546 3712
rect 414664 3528 414716 3534
rect 414664 3470 414716 3476
rect 415504 480 415532 3703
rect 416688 3528 416740 3534
rect 416688 3470 416740 3476
rect 416700 480 416728 3470
rect 417436 2938 417464 13330
rect 417528 3126 417556 16546
rect 421380 13320 421432 13326
rect 421380 13262 421432 13268
rect 418986 3224 419042 3233
rect 418986 3159 419042 3168
rect 417516 3120 417568 3126
rect 417516 3062 417568 3068
rect 417436 2910 417924 2938
rect 417896 480 417924 2910
rect 419000 480 419028 3159
rect 420184 3120 420236 3126
rect 420184 3062 420236 3068
rect 420196 480 420224 3062
rect 421392 480 421420 13262
rect 421576 3806 421604 53586
rect 425704 53508 425756 53514
rect 425704 53450 425756 53456
rect 423772 13252 423824 13258
rect 423772 13194 423824 13200
rect 421564 3800 421616 3806
rect 421564 3742 421616 3748
rect 423680 3800 423732 3806
rect 423680 3742 423732 3748
rect 422574 3632 422630 3641
rect 422574 3567 422630 3576
rect 422588 480 422616 3567
rect 423692 1986 423720 3742
rect 423784 3534 423812 13194
rect 425716 3534 425744 53450
rect 428464 13184 428516 13190
rect 428464 13126 428516 13132
rect 426162 6760 426218 6769
rect 426162 6695 426218 6704
rect 423772 3528 423824 3534
rect 423772 3470 423824 3476
rect 424968 3528 425020 3534
rect 424968 3470 425020 3476
rect 425704 3528 425756 3534
rect 425704 3470 425756 3476
rect 423692 1958 423812 1986
rect 423784 480 423812 1958
rect 424980 480 425008 3470
rect 426176 480 426204 6695
rect 427268 3528 427320 3534
rect 427268 3470 427320 3476
rect 427280 480 427308 3470
rect 428476 480 428504 13126
rect 429658 4040 429714 4049
rect 429658 3975 429714 3984
rect 429672 480 429700 3975
rect 429856 3466 429884 57151
rect 450544 56568 450596 56574
rect 450544 56510 450596 56516
rect 447784 56500 447836 56506
rect 447784 56442 447836 56448
rect 434720 55820 434772 55826
rect 434720 55762 434772 55768
rect 430580 54732 430632 54738
rect 430580 54674 430632 54680
rect 430592 16574 430620 54674
rect 432604 51060 432656 51066
rect 432604 51002 432656 51008
rect 430592 16546 430896 16574
rect 429844 3460 429896 3466
rect 429844 3402 429896 3408
rect 430868 480 430896 16546
rect 432052 13116 432104 13122
rect 432052 13058 432104 13064
rect 432064 480 432092 13058
rect 432616 3806 432644 51002
rect 434732 16574 434760 55762
rect 438860 54664 438912 54670
rect 438860 54606 438912 54612
rect 436744 51876 436796 51882
rect 436744 51818 436796 51824
rect 434732 16546 435588 16574
rect 434444 8356 434496 8362
rect 434444 8298 434496 8304
rect 433246 6488 433302 6497
rect 433246 6423 433302 6432
rect 432604 3800 432656 3806
rect 432604 3742 432656 3748
rect 433260 480 433288 6423
rect 434456 480 434484 8298
rect 435560 480 435588 16546
rect 436650 6352 436706 6361
rect 436650 6287 436706 6296
rect 436664 3210 436692 6287
rect 436756 4146 436784 51818
rect 438872 16574 438900 54606
rect 443644 53576 443696 53582
rect 443644 53518 443696 53524
rect 440240 20120 440292 20126
rect 440240 20062 440292 20068
rect 440252 16574 440280 20062
rect 438872 16546 439176 16574
rect 440252 16546 440372 16574
rect 437940 8424 437992 8430
rect 437940 8366 437992 8372
rect 436744 4140 436796 4146
rect 436744 4082 436796 4088
rect 436664 3182 436784 3210
rect 436756 480 436784 3182
rect 437952 480 437980 8366
rect 439148 480 439176 16546
rect 440344 480 440372 16546
rect 441528 8492 441580 8498
rect 441528 8434 441580 8440
rect 441540 480 441568 8434
rect 442632 4140 442684 4146
rect 442632 4082 442684 4088
rect 442644 480 442672 4082
rect 443656 3670 443684 53518
rect 445760 50992 445812 50998
rect 445760 50934 445812 50940
rect 445772 16574 445800 50934
rect 445772 16546 446260 16574
rect 445024 8560 445076 8566
rect 445024 8502 445076 8508
rect 443644 3664 443696 3670
rect 443644 3606 443696 3612
rect 443826 3496 443882 3505
rect 443826 3431 443882 3440
rect 443840 480 443868 3431
rect 445036 480 445064 8502
rect 446232 480 446260 16546
rect 447416 4208 447468 4214
rect 447416 4150 447468 4156
rect 447428 480 447456 4150
rect 447796 3738 447824 56442
rect 448520 50924 448572 50930
rect 448520 50866 448572 50872
rect 447784 3732 447836 3738
rect 447784 3674 447836 3680
rect 448532 3534 448560 50866
rect 448612 8628 448664 8634
rect 448612 8570 448664 8576
rect 448520 3528 448572 3534
rect 448520 3470 448572 3476
rect 448624 480 448652 8570
rect 450556 3670 450584 56510
rect 454684 56432 454736 56438
rect 454684 56374 454736 56380
rect 452660 53440 452712 53446
rect 452660 53382 452712 53388
rect 452672 16574 452700 53382
rect 454040 20052 454092 20058
rect 454040 19994 454092 20000
rect 454052 16574 454080 19994
rect 452672 16546 453344 16574
rect 454052 16546 454540 16574
rect 452108 8696 452160 8702
rect 452108 8638 452160 8644
rect 450912 4276 450964 4282
rect 450912 4218 450964 4224
rect 450544 3664 450596 3670
rect 450544 3606 450596 3612
rect 449808 3528 449860 3534
rect 449808 3470 449860 3476
rect 449820 480 449848 3470
rect 450924 480 450952 4218
rect 452120 480 452148 8638
rect 453316 480 453344 16546
rect 454512 480 454540 16546
rect 454696 3738 454724 56374
rect 461584 56364 461636 56370
rect 461584 56306 461636 56312
rect 456800 50856 456852 50862
rect 456800 50798 456852 50804
rect 456812 16574 456840 50798
rect 460940 18624 460992 18630
rect 460940 18566 460992 18572
rect 456812 16546 456932 16574
rect 455696 8764 455748 8770
rect 455696 8706 455748 8712
rect 454684 3732 454736 3738
rect 454684 3674 454736 3680
rect 455708 480 455736 8706
rect 456904 480 456932 16546
rect 459192 8832 459244 8838
rect 459192 8774 459244 8780
rect 458088 4344 458140 4350
rect 458088 4286 458140 4292
rect 458100 480 458128 4286
rect 459204 480 459232 8774
rect 460952 6914 460980 18566
rect 461596 16574 461624 56306
rect 479524 56296 479576 56302
rect 479524 56238 479576 56244
rect 468484 56228 468536 56234
rect 468484 56170 468536 56176
rect 463700 50788 463752 50794
rect 463700 50730 463752 50736
rect 463712 16574 463740 50730
rect 467840 19984 467892 19990
rect 467840 19926 467892 19932
rect 467852 16574 467880 19926
rect 461596 16546 461716 16574
rect 463712 16546 464016 16574
rect 467852 16546 468432 16574
rect 460952 6886 461624 6914
rect 460388 3800 460440 3806
rect 460388 3742 460440 3748
rect 460400 480 460428 3742
rect 461596 480 461624 6886
rect 461688 3806 461716 16546
rect 462780 8900 462832 8906
rect 462780 8842 462832 8848
rect 461676 3800 461728 3806
rect 461676 3742 461728 3748
rect 462792 480 462820 8842
rect 463988 480 464016 16546
rect 467472 13932 467524 13938
rect 467472 13874 467524 13880
rect 466276 9648 466328 9654
rect 466276 9590 466328 9596
rect 465170 3360 465226 3369
rect 465170 3295 465226 3304
rect 465184 480 465212 3295
rect 466288 480 466316 9590
rect 467484 480 467512 13874
rect 468404 3482 468432 16546
rect 468496 3874 468524 56170
rect 475384 54596 475436 54602
rect 475384 54538 475436 54544
rect 472624 53372 472676 53378
rect 472624 53314 472676 53320
rect 471060 14000 471112 14006
rect 471060 13942 471112 13948
rect 469864 9580 469916 9586
rect 469864 9522 469916 9528
rect 468484 3868 468536 3874
rect 468484 3810 468536 3816
rect 468404 3454 468708 3482
rect 468680 480 468708 3454
rect 469876 480 469904 9522
rect 471072 480 471100 13942
rect 472254 6624 472310 6633
rect 472254 6559 472310 6568
rect 472268 480 472296 6559
rect 472636 3942 472664 53314
rect 473360 14068 473412 14074
rect 473360 14010 473412 14016
rect 472624 3936 472676 3942
rect 472624 3878 472676 3884
rect 473372 3398 473400 14010
rect 473452 9512 473504 9518
rect 473452 9454 473504 9460
rect 473360 3392 473412 3398
rect 473360 3334 473412 3340
rect 473464 480 473492 9454
rect 475396 4010 475424 54538
rect 478144 14136 478196 14142
rect 478144 14078 478196 14084
rect 475752 9444 475804 9450
rect 475752 9386 475804 9392
rect 475384 4004 475436 4010
rect 475384 3946 475436 3952
rect 474556 3392 474608 3398
rect 474556 3334 474608 3340
rect 474568 480 474596 3334
rect 475764 480 475792 9386
rect 476948 9376 477000 9382
rect 476948 9318 477000 9324
rect 476960 480 476988 9318
rect 478156 480 478184 14078
rect 479536 4146 479564 56238
rect 483020 56160 483072 56166
rect 483020 56102 483072 56108
rect 483032 16574 483060 56102
rect 500960 56092 501012 56098
rect 500960 56034 501012 56040
rect 500972 16574 501000 56034
rect 507860 56024 507912 56030
rect 507860 55966 507912 55972
rect 502340 53304 502392 53310
rect 502340 53246 502392 53252
rect 502352 16574 502380 53246
rect 507872 16574 507900 55966
rect 519544 55956 519596 55962
rect 519544 55898 519596 55904
rect 512644 53236 512696 53242
rect 512644 53178 512696 53184
rect 483032 16546 484072 16574
rect 500972 16546 501828 16574
rect 502352 16546 503024 16574
rect 507872 16546 508912 16574
rect 481640 14204 481692 14210
rect 481640 14146 481692 14152
rect 479524 4140 479576 4146
rect 479524 4082 479576 4088
rect 480536 4140 480588 4146
rect 480536 4082 480588 4088
rect 479340 2100 479392 2106
rect 479340 2042 479392 2048
rect 479352 480 479380 2042
rect 480548 480 480576 4082
rect 481652 3602 481680 14146
rect 481732 9308 481784 9314
rect 481732 9250 481784 9256
rect 481548 3596 481600 3602
rect 481548 3538 481600 3544
rect 481640 3596 481692 3602
rect 481640 3538 481692 3544
rect 481560 3398 481588 3538
rect 481548 3392 481600 3398
rect 481548 3334 481600 3340
rect 481744 480 481772 9250
rect 482836 3596 482888 3602
rect 482836 3538 482888 3544
rect 482848 480 482876 3538
rect 484044 480 484072 16546
rect 497096 15156 497148 15162
rect 497096 15098 497148 15104
rect 493508 14408 493560 14414
rect 493508 14350 493560 14356
rect 489920 14340 489972 14346
rect 489920 14282 489972 14288
rect 486424 14272 486476 14278
rect 486424 14214 486476 14220
rect 485228 9240 485280 9246
rect 485228 9182 485280 9188
rect 485240 480 485268 9182
rect 486436 480 486464 14214
rect 488816 9172 488868 9178
rect 488816 9114 488868 9120
rect 487620 3392 487672 3398
rect 487620 3334 487672 3340
rect 487632 480 487660 3334
rect 488828 480 488856 9114
rect 489932 480 489960 14282
rect 492312 9104 492364 9110
rect 492312 9046 492364 9052
rect 491116 3664 491168 3670
rect 491116 3606 491168 3612
rect 491128 480 491156 3606
rect 492324 480 492352 9046
rect 493520 480 493548 14350
rect 495900 9036 495952 9042
rect 495900 8978 495952 8984
rect 494704 3732 494756 3738
rect 494704 3674 494756 3680
rect 494716 480 494744 3674
rect 495912 480 495940 8978
rect 497108 480 497136 15098
rect 500592 15088 500644 15094
rect 500592 15030 500644 15036
rect 499396 8968 499448 8974
rect 499396 8910 499448 8916
rect 498200 3800 498252 3806
rect 498200 3742 498252 3748
rect 498212 480 498240 3742
rect 499408 480 499436 8910
rect 500604 480 500632 15030
rect 501800 480 501828 16546
rect 502996 480 503024 16546
rect 504180 15020 504232 15026
rect 504180 14962 504232 14968
rect 504192 480 504220 14962
rect 507676 14952 507728 14958
rect 507676 14894 507728 14900
rect 506480 3936 506532 3942
rect 506480 3878 506532 3884
rect 505376 3868 505428 3874
rect 505376 3810 505428 3816
rect 505388 480 505416 3810
rect 506492 480 506520 3878
rect 507688 480 507716 14894
rect 508884 480 508912 16546
rect 511264 14884 511316 14890
rect 511264 14826 511316 14832
rect 510068 4004 510120 4010
rect 510068 3946 510120 3952
rect 510080 480 510108 3946
rect 511276 480 511304 14826
rect 512460 4412 512512 4418
rect 512460 4354 512512 4360
rect 512472 480 512500 4354
rect 512656 3534 512684 53178
rect 519556 16574 519584 55898
rect 526444 54528 526496 54534
rect 526444 54470 526496 54476
rect 520280 53168 520332 53174
rect 520280 53110 520332 53116
rect 520292 16574 520320 53110
rect 519556 16546 519676 16574
rect 520292 16546 520780 16574
rect 514760 14816 514812 14822
rect 514760 14758 514812 14764
rect 512644 3528 512696 3534
rect 512644 3470 512696 3476
rect 513564 3528 513616 3534
rect 513564 3470 513616 3476
rect 513576 480 513604 3470
rect 514772 480 514800 14758
rect 518348 14748 518400 14754
rect 518348 14690 518400 14696
rect 515956 4480 516008 4486
rect 515956 4422 516008 4428
rect 515968 480 515996 4422
rect 517152 3596 517204 3602
rect 517152 3538 517204 3544
rect 517164 480 517192 3538
rect 518360 480 518388 14690
rect 519544 4548 519596 4554
rect 519544 4490 519596 4496
rect 519556 480 519584 4490
rect 519648 2922 519676 16546
rect 519636 2916 519688 2922
rect 519636 2858 519688 2864
rect 520752 480 520780 16546
rect 521844 14680 521896 14686
rect 521844 14622 521896 14628
rect 521856 480 521884 14622
rect 525432 14612 525484 14618
rect 525432 14554 525484 14560
rect 523040 4616 523092 4622
rect 523040 4558 523092 4564
rect 523052 480 523080 4558
rect 524236 2916 524288 2922
rect 524236 2858 524288 2864
rect 524248 480 524276 2858
rect 525444 480 525472 14554
rect 526456 3534 526484 54470
rect 530584 53100 530636 53106
rect 530584 53042 530636 53048
rect 529020 14544 529072 14550
rect 529020 14486 529072 14492
rect 526628 4684 526680 4690
rect 526628 4626 526680 4632
rect 526444 3528 526496 3534
rect 526444 3470 526496 3476
rect 526640 480 526668 4626
rect 527824 3528 527876 3534
rect 527824 3470 527876 3476
rect 527836 480 527864 3470
rect 529032 480 529060 14486
rect 530124 4752 530176 4758
rect 530124 4694 530176 4700
rect 530136 480 530164 4694
rect 530596 3534 530624 53042
rect 535460 51808 535512 51814
rect 535460 51750 535512 51756
rect 533344 50720 533396 50726
rect 533344 50662 533396 50668
rect 532516 14476 532568 14482
rect 532516 14418 532568 14424
rect 530584 3528 530636 3534
rect 530584 3470 530636 3476
rect 531320 3528 531372 3534
rect 531320 3470 531372 3476
rect 531332 480 531360 3470
rect 532528 480 532556 14418
rect 533356 3534 533384 50662
rect 535472 16574 535500 51750
rect 542360 51740 542412 51746
rect 542360 51682 542412 51688
rect 537484 50652 537536 50658
rect 537484 50594 537536 50600
rect 535472 16546 536144 16574
rect 534908 10192 534960 10198
rect 534908 10134 534960 10140
rect 533712 5500 533764 5506
rect 533712 5442 533764 5448
rect 533344 3528 533396 3534
rect 533344 3470 533396 3476
rect 533724 480 533752 5442
rect 534920 480 534948 10134
rect 536116 480 536144 16546
rect 537208 5432 537260 5438
rect 537208 5374 537260 5380
rect 537220 480 537248 5374
rect 537496 3670 537524 50594
rect 539600 50516 539652 50522
rect 539600 50458 539652 50464
rect 538404 10260 538456 10266
rect 538404 10202 538456 10208
rect 537484 3664 537536 3670
rect 537484 3606 537536 3612
rect 538416 480 538444 10202
rect 539612 480 539640 50458
rect 542372 16574 542400 51682
rect 544384 50584 544436 50590
rect 544384 50526 544436 50532
rect 542372 16546 543228 16574
rect 541992 11008 542044 11014
rect 541992 10950 542044 10956
rect 540796 5364 540848 5370
rect 540796 5306 540848 5312
rect 540808 480 540836 5306
rect 542004 480 542032 10950
rect 543200 480 543228 16546
rect 544292 5296 544344 5302
rect 544292 5238 544344 5244
rect 544304 2666 544332 5238
rect 544396 3602 544424 50526
rect 546500 50448 546552 50454
rect 546500 50390 546552 50396
rect 546512 16574 546540 50390
rect 564440 50380 564492 50386
rect 564440 50322 564492 50328
rect 560300 49020 560352 49026
rect 560300 48962 560352 48968
rect 560312 16574 560340 48962
rect 546512 16546 546724 16574
rect 560312 16546 560892 16574
rect 545488 10940 545540 10946
rect 545488 10882 545540 10888
rect 544384 3596 544436 3602
rect 544384 3538 544436 3544
rect 544304 2638 544424 2666
rect 544396 480 544424 2638
rect 545500 480 545528 10882
rect 546696 480 546724 16546
rect 547880 10872 547932 10878
rect 547880 10814 547932 10820
rect 547892 3398 547920 10814
rect 552664 10804 552716 10810
rect 552664 10746 552716 10752
rect 547972 5228 548024 5234
rect 547972 5170 548024 5176
rect 547880 3392 547932 3398
rect 547880 3334 547932 3340
rect 547984 2666 548012 5170
rect 551468 5160 551520 5166
rect 551468 5102 551520 5108
rect 550272 3664 550324 3670
rect 550272 3606 550324 3612
rect 549076 3392 549128 3398
rect 549076 3334 549128 3340
rect 547892 2638 548012 2666
rect 547892 480 547920 2638
rect 549088 480 549116 3334
rect 550284 480 550312 3606
rect 551480 480 551508 5102
rect 552676 480 552704 10746
rect 556160 10736 556212 10742
rect 556160 10678 556212 10684
rect 554964 5092 555016 5098
rect 554964 5034 555016 5040
rect 553768 3528 553820 3534
rect 553768 3470 553820 3476
rect 553780 480 553808 3470
rect 554976 480 555004 5034
rect 556172 480 556200 10678
rect 559748 10668 559800 10674
rect 559748 10610 559800 10616
rect 558552 5024 558604 5030
rect 558552 4966 558604 4972
rect 557356 3596 557408 3602
rect 557356 3538 557408 3544
rect 557368 480 557396 3538
rect 558564 480 558592 4966
rect 559760 480 559788 10610
rect 560864 480 560892 16546
rect 563244 10600 563296 10606
rect 563244 10542 563296 10548
rect 562048 4956 562100 4962
rect 562048 4898 562100 4904
rect 562060 480 562088 4898
rect 563256 480 563284 10542
rect 564452 480 564480 50322
rect 579988 46912 580040 46918
rect 579988 46854 580040 46860
rect 580000 46345 580028 46854
rect 579986 46336 580042 46345
rect 579986 46271 580042 46280
rect 580276 33153 580304 226879
rect 580354 225720 580410 225729
rect 580354 225655 580410 225664
rect 580368 86193 580396 225655
rect 580354 86184 580410 86193
rect 580354 86119 580410 86128
rect 580356 55888 580408 55894
rect 580356 55830 580408 55836
rect 580262 33144 580318 33153
rect 580262 33079 580318 33088
rect 580080 20664 580132 20670
rect 580080 20606 580132 20612
rect 580092 19825 580120 20606
rect 580078 19816 580134 19825
rect 580078 19751 580134 19760
rect 568028 16108 568080 16114
rect 568028 16050 568080 16056
rect 566832 10532 566884 10538
rect 566832 10474 566884 10480
rect 565634 5128 565690 5137
rect 565634 5063 565690 5072
rect 565648 480 565676 5063
rect 566844 480 566872 10474
rect 568040 480 568068 16050
rect 571524 16040 571576 16046
rect 571524 15982 571576 15988
rect 570328 10464 570380 10470
rect 570328 10406 570380 10412
rect 569132 4888 569184 4894
rect 569132 4830 569184 4836
rect 569144 480 569172 4830
rect 570340 480 570368 10406
rect 571536 480 571564 15982
rect 575112 15972 575164 15978
rect 575112 15914 575164 15920
rect 572720 10396 572772 10402
rect 572720 10338 572772 10344
rect 572732 3534 572760 10338
rect 572810 4992 572866 5001
rect 572810 4927 572866 4936
rect 572720 3528 572772 3534
rect 572720 3470 572772 3476
rect 572824 2530 572852 4927
rect 573916 3528 573968 3534
rect 573916 3470 573968 3476
rect 572732 2502 572852 2530
rect 572732 480 572760 2502
rect 573928 480 573956 3470
rect 575124 480 575152 15914
rect 578608 15904 578660 15910
rect 578608 15846 578660 15852
rect 577412 10328 577464 10334
rect 577412 10270 577464 10276
rect 576306 4856 576362 4865
rect 576306 4791 576362 4800
rect 576320 480 576348 4791
rect 577424 480 577452 10270
rect 578620 480 578648 15846
rect 580368 6633 580396 55830
rect 580354 6624 580410 6633
rect 580354 6559 580410 6568
rect 582194 6216 582250 6225
rect 582194 6151 582250 6160
rect 581000 4820 581052 4826
rect 581000 4762 581052 4768
rect 581012 480 581040 4762
rect 582208 480 582236 6151
rect 583392 3460 583444 3466
rect 583392 3402 583444 3408
rect 583404 480 583432 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13514 -960 13626 480
rect 14710 -960 14822 480
rect 15906 -960 16018 480
rect 17010 -960 17122 480
rect 18206 -960 18318 480
rect 19402 -960 19514 480
rect 20598 -960 20710 480
rect 21794 -960 21906 480
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 27682 -960 27794 480
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 34766 -960 34878 480
rect 35962 -960 36074 480
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 43046 -960 43158 480
rect 44242 -960 44354 480
rect 45438 -960 45550 480
rect 46634 -960 46746 480
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 52522 -960 52634 480
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58410 -960 58522 480
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 70278 -960 70390 480
rect 71474 -960 71586 480
rect 72578 -960 72690 480
rect 73774 -960 73886 480
rect 74970 -960 75082 480
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 130538 -960 130650 480
rect 131734 -960 131846 480
rect 132930 -960 133042 480
rect 134126 -960 134238 480
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 141210 -960 141322 480
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 148294 -960 148406 480
rect 149490 -960 149602 480
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 156574 -960 156686 480
rect 157770 -960 157882 480
rect 158874 -960 158986 480
rect 160070 -960 160182 480
rect 161266 -960 161378 480
rect 162462 -960 162574 480
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 174238 -960 174350 480
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177826 -960 177938 480
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184910 -960 185022 480
rect 186106 -960 186218 480
rect 187302 -960 187414 480
rect 188498 -960 188610 480
rect 189694 -960 189806 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197882 -960 197994 480
rect 199078 -960 199190 480
rect 200274 -960 200386 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206162 -960 206274 480
rect 207358 -960 207470 480
rect 208554 -960 208666 480
rect 209750 -960 209862 480
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 213338 -960 213450 480
rect 214442 -960 214554 480
rect 215638 -960 215750 480
rect 216834 -960 216946 480
rect 218030 -960 218142 480
rect 219226 -960 219338 480
rect 220422 -960 220534 480
rect 221526 -960 221638 480
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 226310 -960 226422 480
rect 227506 -960 227618 480
rect 228702 -960 228814 480
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232198 -960 232310 480
rect 233394 -960 233506 480
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 240478 -960 240590 480
rect 241674 -960 241786 480
rect 242870 -960 242982 480
rect 244066 -960 244178 480
rect 245170 -960 245282 480
rect 246366 -960 246478 480
rect 247562 -960 247674 480
rect 248758 -960 248870 480
rect 249954 -960 250066 480
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255842 -960 255954 480
rect 257038 -960 257150 480
rect 258234 -960 258346 480
rect 259430 -960 259542 480
rect 260626 -960 260738 480
rect 261730 -960 261842 480
rect 262926 -960 263038 480
rect 264122 -960 264234 480
rect 265318 -960 265430 480
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268814 -960 268926 480
rect 270010 -960 270122 480
rect 271206 -960 271318 480
rect 272402 -960 272514 480
rect 273598 -960 273710 480
rect 274794 -960 274906 480
rect 275990 -960 276102 480
rect 277094 -960 277206 480
rect 278290 -960 278402 480
rect 279486 -960 279598 480
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283074 -960 283186 480
rect 284270 -960 284382 480
rect 285374 -960 285486 480
rect 286570 -960 286682 480
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 290158 -960 290270 480
rect 291354 -960 291466 480
rect 292550 -960 292662 480
rect 293654 -960 293766 480
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 297242 -960 297354 480
rect 298438 -960 298550 480
rect 299634 -960 299746 480
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 303130 -960 303242 480
rect 304326 -960 304438 480
rect 305522 -960 305634 480
rect 306718 -960 306830 480
rect 307914 -960 308026 480
rect 309018 -960 309130 480
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312606 -960 312718 480
rect 313802 -960 313914 480
rect 314998 -960 315110 480
rect 316194 -960 316306 480
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 319690 -960 319802 480
rect 320886 -960 320998 480
rect 322082 -960 322194 480
rect 323278 -960 323390 480
rect 324382 -960 324494 480
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327970 -960 328082 480
rect 329166 -960 329278 480
rect 330362 -960 330474 480
rect 331558 -960 331670 480
rect 332662 -960 332774 480
rect 333858 -960 333970 480
rect 335054 -960 335166 480
rect 336250 -960 336362 480
rect 337446 -960 337558 480
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340942 -960 341054 480
rect 342138 -960 342250 480
rect 343334 -960 343446 480
rect 344530 -960 344642 480
rect 345726 -960 345838 480
rect 346922 -960 347034 480
rect 348026 -960 348138 480
rect 349222 -960 349334 480
rect 350418 -960 350530 480
rect 351614 -960 351726 480
rect 352810 -960 352922 480
rect 354006 -960 354118 480
rect 355202 -960 355314 480
rect 356306 -960 356418 480
rect 357502 -960 357614 480
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 -960 361202 480
rect 362286 -960 362398 480
rect 363482 -960 363594 480
rect 364586 -960 364698 480
rect 365782 -960 365894 480
rect 366978 -960 367090 480
rect 368174 -960 368286 480
rect 369370 -960 369482 480
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372866 -960 372978 480
rect 374062 -960 374174 480
rect 375258 -960 375370 480
rect 376454 -960 376566 480
rect 377650 -960 377762 480
rect 378846 -960 378958 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384734 -960 384846 480
rect 385930 -960 386042 480
rect 387126 -960 387238 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395314 -960 395426 480
rect 396510 -960 396622 480
rect 397706 -960 397818 480
rect 398902 -960 399014 480
rect 400098 -960 400210 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404790 -960 404902 480
rect 405986 -960 406098 480
rect 407182 -960 407294 480
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410770 -960 410882 480
rect 411874 -960 411986 480
rect 413070 -960 413182 480
rect 414266 -960 414378 480
rect 415462 -960 415574 480
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418958 -960 419070 480
rect 420154 -960 420266 480
rect 421350 -960 421462 480
rect 422546 -960 422658 480
rect 423742 -960 423854 480
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429630 -960 429742 480
rect 430826 -960 430938 480
rect 432022 -960 432134 480
rect 433218 -960 433330 480
rect 434414 -960 434526 480
rect 435518 -960 435630 480
rect 436714 -960 436826 480
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446190 -960 446302 480
rect 447386 -960 447498 480
rect 448582 -960 448694 480
rect 449778 -960 449890 480
rect 450882 -960 450994 480
rect 452078 -960 452190 480
rect 453274 -960 453386 480
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 461554 -960 461666 480
rect 462750 -960 462862 480
rect 463946 -960 464058 480
rect 465142 -960 465254 480
rect 466246 -960 466358 480
rect 467442 -960 467554 480
rect 468638 -960 468750 480
rect 469834 -960 469946 480
rect 471030 -960 471142 480
rect 472226 -960 472338 480
rect 473422 -960 473534 480
rect 474526 -960 474638 480
rect 475722 -960 475834 480
rect 476918 -960 477030 480
rect 478114 -960 478226 480
rect 479310 -960 479422 480
rect 480506 -960 480618 480
rect 481702 -960 481814 480
rect 482806 -960 482918 480
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488786 -960 488898 480
rect 489890 -960 490002 480
rect 491086 -960 491198 480
rect 492282 -960 492394 480
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495870 -960 495982 480
rect 497066 -960 497178 480
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 501758 -960 501870 480
rect 502954 -960 503066 480
rect 504150 -960 504262 480
rect 505346 -960 505458 480
rect 506450 -960 506562 480
rect 507646 -960 507758 480
rect 508842 -960 508954 480
rect 510038 -960 510150 480
rect 511234 -960 511346 480
rect 512430 -960 512542 480
rect 513534 -960 513646 480
rect 514730 -960 514842 480
rect 515926 -960 516038 480
rect 517122 -960 517234 480
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520710 -960 520822 480
rect 521814 -960 521926 480
rect 523010 -960 523122 480
rect 524206 -960 524318 480
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527794 -960 527906 480
rect 528990 -960 529102 480
rect 530094 -960 530206 480
rect 531290 -960 531402 480
rect 532486 -960 532598 480
rect 533682 -960 533794 480
rect 534878 -960 534990 480
rect 536074 -960 536186 480
rect 537178 -960 537290 480
rect 538374 -960 538486 480
rect 539570 -960 539682 480
rect 540766 -960 540878 480
rect 541962 -960 542074 480
rect 543158 -960 543270 480
rect 544354 -960 544466 480
rect 545458 -960 545570 480
rect 546654 -960 546766 480
rect 547850 -960 547962 480
rect 549046 -960 549158 480
rect 550242 -960 550354 480
rect 551438 -960 551550 480
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554934 -960 555046 480
rect 556130 -960 556242 480
rect 557326 -960 557438 480
rect 558522 -960 558634 480
rect 559718 -960 559830 480
rect 560822 -960 560934 480
rect 562018 -960 562130 480
rect 563214 -960 563326 480
rect 564410 -960 564522 480
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 2778 684256 2834 684312
rect 3514 671200 3570 671256
rect 3422 658144 3478 658200
rect 3422 632068 3424 632088
rect 3424 632068 3476 632088
rect 3476 632068 3478 632088
rect 3422 632032 3478 632068
rect 3146 619112 3202 619168
rect 3238 606056 3294 606112
rect 3330 579944 3386 580000
rect 3422 566888 3478 566944
rect 3422 553832 3478 553888
rect 3422 527856 3478 527912
rect 3422 514820 3478 514856
rect 3422 514800 3424 514820
rect 3424 514800 3476 514820
rect 3476 514800 3478 514820
rect 3054 501744 3110 501800
rect 3422 475632 3478 475688
rect 3238 462576 3294 462632
rect 3146 449520 3202 449576
rect 3422 423544 3478 423600
rect 3146 410488 3202 410544
rect 3422 397468 3424 397488
rect 3424 397468 3476 397488
rect 3476 397468 3478 397488
rect 3422 397432 3478 397468
rect 3422 371320 3478 371376
rect 3146 358400 3202 358456
rect 3330 345344 3386 345400
rect 3422 319232 3478 319288
rect 3238 306176 3294 306232
rect 3422 293120 3478 293176
rect 3054 267144 3110 267200
rect 58714 489912 58770 489968
rect 53654 488824 53710 488880
rect 53562 484744 53618 484800
rect 53378 484608 53434 484664
rect 3422 254088 3478 254144
rect 3422 249056 3478 249112
rect 4066 241032 4122 241088
rect 4158 235184 4214 235240
rect 21362 233688 21418 233744
rect 18602 233552 18658 233608
rect 14462 231920 14518 231976
rect 11702 231104 11758 231160
rect 7562 230968 7618 231024
rect 4802 230832 4858 230888
rect 3606 228520 3662 228576
rect 3422 228248 3478 228304
rect 2778 214920 2834 214976
rect 3146 188808 3202 188864
rect 3330 162832 3386 162888
rect 3330 136720 3386 136776
rect 3146 110608 3202 110664
rect 3238 97552 3294 97608
rect 3330 84632 3386 84688
rect 3330 71576 3386 71632
rect 3514 227024 3570 227080
rect 3698 227160 3754 227216
rect 3606 201864 3662 201920
rect 3698 149776 3754 149832
rect 15842 230696 15898 230752
rect 3514 58520 3570 58576
rect 12346 57568 12402 57624
rect 10966 57432 11022 57488
rect 9586 57296 9642 57352
rect 4066 57160 4122 57216
rect 3422 45464 3478 45520
rect 2870 32408 2926 32464
rect 3422 19352 3478 19408
rect 3422 6432 3478 6488
rect 570 3304 626 3360
rect 15106 57024 15162 57080
rect 13726 56888 13782 56944
rect 17222 226752 17278 226808
rect 25502 229472 25558 229528
rect 22742 228384 22798 228440
rect 17866 56752 17922 56808
rect 29642 229336 29698 229392
rect 55034 487872 55090 487928
rect 54942 487464 54998 487520
rect 53746 487192 53802 487248
rect 56874 487328 56930 487384
rect 56506 485968 56562 486024
rect 55126 484880 55182 484936
rect 56414 483928 56470 483984
rect 55678 226480 55734 226536
rect 55770 226344 55826 226400
rect 55862 207304 55918 207360
rect 55954 189488 56010 189544
rect 56046 177520 56102 177576
rect 56230 222264 56286 222320
rect 56414 216280 56470 216336
rect 56322 147736 56378 147792
rect 56690 435376 56746 435432
rect 56598 407496 56654 407552
rect 56138 73208 56194 73264
rect 56782 225936 56838 225992
rect 56782 171536 56838 171592
rect 58622 485016 58678 485072
rect 57518 484200 57574 484256
rect 57426 432384 57482 432440
rect 57334 430616 57390 430672
rect 57242 429392 57298 429448
rect 57058 237904 57114 237960
rect 57334 239400 57390 239456
rect 57242 186496 57298 186552
rect 57150 117952 57206 118008
rect 57058 108976 57114 109032
rect 57242 82184 57298 82240
rect 57150 79192 57206 79248
rect 56874 64232 56930 64288
rect 57610 436328 57666 436384
rect 57518 210296 57574 210352
rect 57518 195336 57574 195392
rect 57518 192480 57574 192536
rect 57518 183504 57574 183560
rect 57426 162560 57482 162616
rect 57426 156712 57482 156768
rect 57426 153720 57482 153776
rect 57426 150728 57482 150784
rect 57426 144744 57482 144800
rect 57702 433336 57758 433392
rect 57886 427896 57942 427952
rect 57794 409944 57850 410000
rect 58346 242120 58402 242176
rect 58254 236544 58310 236600
rect 58162 232600 58218 232656
rect 57794 227704 57850 227760
rect 57702 226208 57758 226264
rect 57610 135768 57666 135824
rect 57610 126948 57666 126984
rect 57610 126928 57612 126948
rect 57612 126928 57664 126948
rect 57664 126928 57666 126948
rect 57610 120944 57666 121000
rect 57886 226072 57942 226128
rect 57794 219272 57850 219328
rect 57886 198328 57942 198384
rect 57794 168544 57850 168600
rect 57794 159704 57850 159760
rect 57794 141752 57850 141808
rect 57794 132776 57850 132832
rect 58162 129784 58218 129840
rect 57702 114960 57758 115016
rect 57610 111968 57666 112024
rect 57610 105984 57666 106040
rect 57610 102992 57666 103048
rect 57610 100000 57666 100056
rect 58254 94152 58310 94208
rect 57518 91160 57574 91216
rect 57610 88168 57666 88224
rect 58438 201320 58494 201376
rect 58622 232736 58678 232792
rect 58622 227296 58678 227352
rect 58530 165552 58586 165608
rect 58346 85176 58402 85232
rect 57610 70216 57666 70272
rect 57334 61376 57390 61432
rect 56506 57704 56562 57760
rect 56506 57296 56562 57352
rect 59082 490048 59138 490104
rect 58990 488688 59046 488744
rect 58898 488552 58954 488608
rect 58714 204312 58770 204368
rect 58898 180512 58954 180568
rect 58806 97008 58862 97064
rect 58990 174528 59046 174584
rect 59174 488960 59230 489016
rect 59082 123936 59138 123992
rect 103978 491408 104034 491464
rect 101678 491272 101734 491328
rect 99194 487736 99250 487792
rect 101678 486512 101734 486568
rect 103978 486512 104034 486568
rect 99194 485968 99250 486024
rect 60002 485152 60058 485208
rect 88338 485152 88394 485208
rect 59266 484472 59322 484528
rect 59174 76200 59230 76256
rect 59450 484064 59506 484120
rect 59358 408176 59414 408232
rect 59450 213288 59506 213344
rect 108762 490184 108818 490240
rect 178314 488960 178370 489016
rect 130842 487872 130898 487928
rect 126334 487600 126390 487656
rect 126334 486648 126390 486704
rect 130842 486648 130898 486704
rect 108762 486512 108818 486568
rect 178314 485560 178370 485616
rect 104898 485016 104954 485072
rect 85394 398112 85450 398168
rect 113638 398112 113694 398168
rect 78310 397296 78366 397352
rect 79966 397296 80022 397352
rect 80426 397296 80482 397352
rect 83278 397296 83334 397352
rect 60002 229880 60058 229936
rect 61106 226616 61162 226672
rect 60186 226344 60242 226400
rect 61106 226208 61162 226264
rect 61290 226888 61346 226944
rect 61750 226344 61806 226400
rect 77206 396752 77262 396808
rect 75918 396616 75974 396672
rect 73618 234640 73674 234696
rect 67546 233416 67602 233472
rect 64786 233280 64842 233336
rect 63406 230288 63462 230344
rect 62762 227704 62818 227760
rect 66350 229200 66406 229256
rect 65338 227840 65394 227896
rect 72698 232056 72754 232112
rect 69294 230560 69350 230616
rect 70306 229608 70362 229664
rect 70306 228520 70362 228576
rect 71226 227976 71282 228032
rect 70306 227704 70362 227760
rect 74538 229744 74594 229800
rect 74262 228112 74318 228168
rect 82726 396752 82782 396808
rect 78586 247016 78642 247072
rect 76562 234776 76618 234832
rect 75918 227296 75974 227352
rect 74538 227160 74594 227216
rect 80610 236272 80666 236328
rect 86498 397296 86554 397352
rect 87694 397332 87696 397352
rect 87696 397332 87748 397352
rect 87748 397332 87750 397352
rect 87694 397296 87750 397332
rect 88706 397296 88762 397352
rect 92294 397296 92350 397352
rect 93490 397296 93546 397352
rect 96526 397296 96582 397352
rect 98918 397296 98974 397352
rect 100114 397296 100170 397352
rect 101586 397296 101642 397352
rect 101862 397296 101918 397352
rect 102874 397296 102930 397352
rect 103702 397296 103758 397352
rect 105910 397296 105966 397352
rect 107198 397296 107254 397352
rect 109774 397296 109830 397352
rect 111614 397296 111670 397352
rect 85486 396752 85542 396808
rect 96434 397160 96490 397216
rect 89626 396752 89682 396808
rect 91006 396752 91062 396808
rect 93766 396752 93822 396808
rect 95146 396752 95202 396808
rect 86222 257896 86278 257952
rect 86222 236272 86278 236328
rect 85486 232464 85542 232520
rect 89718 396616 89774 396672
rect 91098 396616 91154 396672
rect 91098 232600 91154 232656
rect 98458 397160 98514 397216
rect 97906 396752 97962 396808
rect 101954 396752 102010 396808
rect 104806 397160 104862 397216
rect 101126 233824 101182 233880
rect 102046 233824 102102 233880
rect 104070 233824 104126 233880
rect 106002 396752 106058 396808
rect 104806 238040 104862 238096
rect 104714 233824 104770 233880
rect 107382 396752 107438 396808
rect 108854 396752 108910 396808
rect 106002 232600 106058 232656
rect 111522 396752 111578 396808
rect 108946 396616 109002 396672
rect 113178 397160 113234 397216
rect 113086 396752 113142 396808
rect 108946 244840 109002 244896
rect 114466 397296 114522 397352
rect 115846 397296 115902 397352
rect 118146 397296 118202 397352
rect 117226 396752 117282 396808
rect 117134 396616 117190 396672
rect 113086 243480 113142 243536
rect 114926 233824 114982 233880
rect 115846 233824 115902 233880
rect 118606 396752 118662 396808
rect 119894 396752 119950 396808
rect 117226 242256 117282 242312
rect 118606 249192 118662 249248
rect 121366 396752 121422 396808
rect 124126 396752 124182 396808
rect 124126 250416 124182 250472
rect 124126 240760 124182 240816
rect 122654 236680 122710 236736
rect 136454 397296 136510 397352
rect 138478 397296 138534 397352
rect 126886 396752 126942 396808
rect 129646 396752 129702 396808
rect 131026 396752 131082 396808
rect 133786 396752 133842 396808
rect 125138 232736 125194 232792
rect 128358 230424 128414 230480
rect 127530 229880 127586 229936
rect 129186 230424 129242 230480
rect 131118 230424 131174 230480
rect 140778 396752 140834 396808
rect 144826 396752 144882 396808
rect 146206 396752 146262 396808
rect 132130 230424 132186 230480
rect 135258 230424 135314 230480
rect 135994 230424 136050 230480
rect 138018 230424 138074 230480
rect 141422 255856 141478 255912
rect 138202 245656 138258 245712
rect 138202 240760 138258 240816
rect 138938 230424 138994 230480
rect 141422 245656 141478 245712
rect 142158 230424 142214 230480
rect 142986 230424 143042 230480
rect 146206 232736 146262 232792
rect 150714 397296 150770 397352
rect 147678 396752 147734 396808
rect 154486 396752 154542 396808
rect 155958 396752 156014 396808
rect 158626 396752 158682 396808
rect 161386 396752 161442 396808
rect 164146 396752 164202 396808
rect 166906 396752 166962 396808
rect 146942 255856 146998 255912
rect 146298 230424 146354 230480
rect 146850 230424 146906 230480
rect 153198 230424 153254 230480
rect 155958 249056 156014 249112
rect 153842 230424 153898 230480
rect 156050 235184 156106 235240
rect 158626 240760 158682 240816
rect 164606 233688 164662 233744
rect 161662 233552 161718 233608
rect 161018 230968 161074 231024
rect 158074 230832 158130 230888
rect 160190 229744 160246 229800
rect 160098 229608 160154 229664
rect 160098 228248 160154 228304
rect 158810 226752 158866 226808
rect 164054 231104 164110 231160
rect 163042 229880 163098 229936
rect 166998 231920 167054 231976
rect 165986 229472 166042 229528
rect 169942 230696 169998 230752
rect 167918 229608 167974 229664
rect 168562 227024 168618 227080
rect 171874 229336 171930 229392
rect 170954 228384 171010 228440
rect 174174 233824 174230 233880
rect 183466 397296 183522 397352
rect 183190 396752 183246 396808
rect 175186 233824 175242 233880
rect 179786 229744 179842 229800
rect 181166 226752 181222 226808
rect 183742 230152 183798 230208
rect 182730 229880 182786 229936
rect 182086 226752 182142 226808
rect 184754 230016 184810 230072
rect 187974 233824 188030 233880
rect 188986 233824 189042 233880
rect 190918 233824 190974 233880
rect 191746 233824 191802 233880
rect 196714 487736 196770 487792
rect 196530 236680 196586 236736
rect 196806 483384 196862 483440
rect 196714 230152 196770 230208
rect 197910 486920 197966 486976
rect 197358 479168 197414 479224
rect 196806 229744 196862 229800
rect 197358 239400 197414 239456
rect 198646 486648 198702 486704
rect 198278 486376 198334 486432
rect 198094 485832 198150 485888
rect 197910 239400 197966 239456
rect 198462 486104 198518 486160
rect 198370 485560 198426 485616
rect 198278 231104 198334 231160
rect 198554 483928 198610 483984
rect 198462 236816 198518 236872
rect 198370 230016 198426 230072
rect 198830 419328 198886 419384
rect 198738 417696 198794 417752
rect 198646 236680 198702 236736
rect 199014 416336 199070 416392
rect 198922 413616 198978 413672
rect 199382 414840 199438 414896
rect 198830 242120 198886 242176
rect 198738 236544 198794 236600
rect 198554 229880 198610 229936
rect 198094 229744 198150 229800
rect 199382 228248 199438 228304
rect 202878 487600 202934 487656
rect 202142 486512 202198 486568
rect 201774 233824 201830 233880
rect 203522 486240 203578 486296
rect 202786 233824 202842 233880
rect 202142 231240 202198 231296
rect 203522 235184 203578 235240
rect 205638 234776 205694 234832
rect 205638 231920 205694 231976
rect 209778 485288 209834 485344
rect 211342 230424 211398 230480
rect 213182 230424 213238 230480
rect 266082 490048 266138 490104
rect 217782 488960 217838 489016
rect 263598 488960 263654 489016
rect 217690 487600 217746 487656
rect 217322 487192 217378 487248
rect 216586 485288 216642 485344
rect 215574 233824 215630 233880
rect 217414 486784 217470 486840
rect 217322 484472 217378 484528
rect 216678 435920 216734 435976
rect 216678 433744 216734 433800
rect 216678 432792 216734 432848
rect 216678 429936 216734 429992
rect 217230 428168 217286 428224
rect 216678 409944 216734 410000
rect 217138 408040 217194 408096
rect 217322 408312 217378 408368
rect 216586 233824 216642 233880
rect 217138 233824 217194 233880
rect 217598 485832 217654 485888
rect 217506 431024 217562 431080
rect 256146 487600 256202 487656
rect 217874 487464 217930 487520
rect 218242 486920 218298 486976
rect 218058 484472 218114 484528
rect 217966 436872 218022 436928
rect 217874 398112 217930 398168
rect 217690 235864 217746 235920
rect 217414 227024 217470 227080
rect 218150 483520 218206 483576
rect 218058 397976 218114 398032
rect 218978 486784 219034 486840
rect 218610 486648 218666 486704
rect 218426 486376 218482 486432
rect 218334 483656 218390 483712
rect 218242 399472 218298 399528
rect 218150 231648 218206 231704
rect 218518 485152 218574 485208
rect 218426 267688 218482 267744
rect 218426 258304 218482 258360
rect 218426 257896 218482 257952
rect 218426 248376 218482 248432
rect 218426 247968 218482 248024
rect 218426 238856 218482 238912
rect 218702 485968 218758 486024
rect 218610 398248 218666 398304
rect 218610 393352 218666 393408
rect 218334 231376 218390 231432
rect 218518 238448 218574 238504
rect 218518 235048 218574 235104
rect 218426 230968 218482 231024
rect 217966 229880 218022 229936
rect 77390 226616 77446 226672
rect 62118 226480 62174 226536
rect 75550 226480 75606 226536
rect 68558 226344 68614 226400
rect 218794 485016 218850 485072
rect 218886 483248 218942 483304
rect 219990 486512 220046 486568
rect 219806 486240 219862 486296
rect 219346 486104 219402 486160
rect 219254 485696 219310 485752
rect 219162 483792 219218 483848
rect 219070 483248 219126 483304
rect 219070 383560 219126 383616
rect 219070 374176 219126 374232
rect 218978 373904 219034 373960
rect 218978 364384 219034 364440
rect 218978 364248 219034 364304
rect 218978 354728 219034 354784
rect 218978 354592 219034 354648
rect 218978 345072 219034 345128
rect 219070 344528 219126 344584
rect 219070 335416 219126 335472
rect 219070 325624 219126 325680
rect 219070 316240 219126 316296
rect 218978 315968 219034 316024
rect 218978 306448 219034 306504
rect 218978 306312 219034 306368
rect 218978 296792 219034 296848
rect 218978 296656 219034 296712
rect 218978 287136 219034 287192
rect 218978 287000 219034 287056
rect 218978 277480 219034 277536
rect 218978 277344 219034 277400
rect 218978 267824 219034 267880
rect 218886 231784 218942 231840
rect 218794 228656 218850 228712
rect 219070 230016 219126 230072
rect 219622 485968 219678 486024
rect 219714 485152 219770 485208
rect 219622 484200 219678 484256
rect 219438 484064 219494 484120
rect 219530 483792 219586 483848
rect 219622 483656 219678 483712
rect 219714 403144 219770 403200
rect 219346 392808 219402 392864
rect 219346 383832 219402 383888
rect 219346 335008 219402 335064
rect 219346 325896 219402 325952
rect 219254 231512 219310 231568
rect 219162 228520 219218 228576
rect 219898 483520 219954 483576
rect 219898 402872 219954 402928
rect 219806 233960 219862 234016
rect 219346 227160 219402 227216
rect 316038 489912 316094 489968
rect 276202 488824 276258 488880
rect 266082 486784 266138 486840
rect 301042 488688 301098 488744
rect 256146 485832 256202 485888
rect 263598 485832 263654 485888
rect 276202 485832 276258 485888
rect 303434 488552 303490 488608
rect 318706 487328 318762 487384
rect 316038 486512 316094 486568
rect 340142 487192 340198 487248
rect 315946 486376 316002 486432
rect 318706 486376 318762 486432
rect 340142 486376 340198 486432
rect 303434 485832 303490 485888
rect 301042 485016 301098 485072
rect 356518 485832 356574 485888
rect 315946 483792 316002 483848
rect 220082 399880 220138 399936
rect 220082 235864 220138 235920
rect 219898 228384 219954 228440
rect 223210 230016 223266 230072
rect 224590 229200 224646 229256
rect 61934 226208 61990 226264
rect 218702 226208 218758 226264
rect 220542 226208 220598 226264
rect 223578 226208 223634 226264
rect 224590 226208 224646 226264
rect 59542 138760 59598 138816
rect 59266 67224 59322 67280
rect 224406 60288 224462 60344
rect 222658 60152 222714 60208
rect 58898 57840 58954 57896
rect 58622 57024 58678 57080
rect 55678 3576 55734 3632
rect 60002 57432 60058 57488
rect 60922 57160 60978 57216
rect 59726 3596 59782 3632
rect 59726 3576 59728 3596
rect 59728 3576 59780 3596
rect 59780 3576 59782 3596
rect 62118 57704 62174 57760
rect 61842 57180 61898 57216
rect 62670 57568 62726 57624
rect 62946 57432 63002 57488
rect 62394 57296 62450 57352
rect 61842 57160 61844 57180
rect 61844 57160 61896 57180
rect 61896 57160 61898 57180
rect 59358 3304 59414 3360
rect 63590 56888 63646 56944
rect 63774 56888 63830 56944
rect 63222 56752 63278 56808
rect 63406 56788 63408 56808
rect 63408 56788 63460 56808
rect 63460 56788 63462 56808
rect 63406 56752 63462 56788
rect 64142 56616 64198 56672
rect 65522 56908 65578 56944
rect 65522 56888 65524 56908
rect 65524 56888 65576 56908
rect 65576 56888 65578 56908
rect 65614 56788 65616 56808
rect 65616 56788 65668 56808
rect 65668 56788 65670 56808
rect 65614 56752 65670 56788
rect 66902 57160 66958 57216
rect 103058 57432 103114 57488
rect 103518 57432 103574 57488
rect 116858 57024 116914 57080
rect 117502 56616 117558 56672
rect 118330 57160 118386 57216
rect 118606 56888 118662 56944
rect 118606 56772 118662 56808
rect 118606 56752 118608 56772
rect 118608 56752 118660 56772
rect 118660 56752 118662 56772
rect 118790 56752 118846 56808
rect 118974 57024 119030 57080
rect 120998 57296 121054 57352
rect 123482 56616 123538 56672
rect 126334 56888 126390 56944
rect 129186 57024 129242 57080
rect 129922 56888 129978 56944
rect 131946 57432 132002 57488
rect 132866 57432 132922 57488
rect 132498 56888 132554 56944
rect 132682 56888 132738 56944
rect 133050 57024 133106 57080
rect 134798 57024 134854 57080
rect 136822 56772 136878 56808
rect 136822 56752 136824 56772
rect 136824 56752 136876 56772
rect 136876 56752 136878 56772
rect 137926 56888 137982 56944
rect 140410 57432 140466 57488
rect 142066 57160 142122 57216
rect 142250 57160 142306 57216
rect 142894 57024 142950 57080
rect 143906 57568 143962 57624
rect 146298 57296 146354 57352
rect 151726 5752 151782 5808
rect 158626 6840 158682 6896
rect 157246 6024 157302 6080
rect 155866 5888 155922 5944
rect 160466 57432 160522 57488
rect 161110 3848 161166 3904
rect 162582 3712 162638 3768
rect 163870 3576 163926 3632
rect 166354 57044 166410 57080
rect 166354 57024 166356 57044
rect 166356 57024 166408 57044
rect 166408 57024 166410 57044
rect 165250 6704 165306 6760
rect 166630 6432 166686 6488
rect 168654 57060 168656 57080
rect 168656 57060 168708 57080
rect 168708 57060 168710 57080
rect 168654 57024 168710 57060
rect 168010 6296 168066 6352
rect 171046 57568 171102 57624
rect 169666 3440 169722 3496
rect 171598 57568 171654 57624
rect 175186 3304 175242 3360
rect 180706 56772 180762 56808
rect 180706 56752 180708 56772
rect 180708 56752 180760 56772
rect 180760 56752 180762 56772
rect 180798 56652 180800 56672
rect 180800 56652 180852 56672
rect 180852 56652 180854 56672
rect 180798 56616 180854 56652
rect 199658 5072 199714 5128
rect 203522 57160 203578 57216
rect 201406 4936 201462 4992
rect 202786 4800 202842 4856
rect 204074 6160 204130 6216
rect 204718 59744 204774 59800
rect 206190 58656 206246 58712
rect 204442 56752 204498 56808
rect 207018 57704 207074 57760
rect 206742 57568 206798 57624
rect 209042 59608 209098 59664
rect 209962 57704 210018 57760
rect 209686 57432 209742 57488
rect 210514 57840 210570 57896
rect 208766 56888 208822 56944
rect 211894 60016 211950 60072
rect 211434 57840 211490 57896
rect 211158 56616 211214 56672
rect 210422 6568 210478 6624
rect 213182 3984 213238 4040
rect 214654 58520 214710 58576
rect 218150 59200 218206 59256
rect 218702 58928 218758 58984
rect 213550 3168 213606 3224
rect 213458 3032 213514 3088
rect 219254 59064 219310 59120
rect 219622 58928 219678 58984
rect 219622 58520 219678 58576
rect 219254 57704 219310 57760
rect 218978 57024 219034 57080
rect 220174 59200 220230 59256
rect 220450 57840 220506 57896
rect 221646 59336 221702 59392
rect 221830 58248 221886 58304
rect 222750 59472 222806 59528
rect 223578 60016 223634 60072
rect 224406 59744 224462 59800
rect 223578 59064 223634 59120
rect 223946 59064 224002 59120
rect 223486 57704 223542 57760
rect 224314 59064 224370 59120
rect 224406 58248 224462 58304
rect 225326 244840 225382 244896
rect 225234 64096 225290 64152
rect 225418 240760 225474 240816
rect 225326 60424 225382 60480
rect 225326 60288 225382 60344
rect 225234 60152 225290 60208
rect 225142 57432 225198 57488
rect 225510 238040 225566 238096
rect 225786 232736 225842 232792
rect 225694 232600 225750 232656
rect 225602 232464 225658 232520
rect 225878 231376 225934 231432
rect 225786 65592 225842 65648
rect 225970 228248 226026 228304
rect 226246 250416 226302 250472
rect 226338 231512 226394 231568
rect 226338 222672 226394 222728
rect 226338 204176 226394 204232
rect 226338 203496 226394 203552
rect 226246 148824 226302 148880
rect 226246 147736 226302 147792
rect 226154 143520 226210 143576
rect 226154 143384 226210 143440
rect 226062 132368 226118 132424
rect 225970 65592 226026 65648
rect 225878 65456 225934 65512
rect 226062 65456 226118 65512
rect 225970 65320 226026 65376
rect 225786 65184 225842 65240
rect 225694 62736 225750 62792
rect 225694 60424 225750 60480
rect 225602 57568 225658 57624
rect 225878 62736 225934 62792
rect 226062 60016 226118 60072
rect 226982 239400 227038 239456
rect 226614 235184 226670 235240
rect 226522 181736 226578 181792
rect 226430 146104 226486 146160
rect 226798 231240 226854 231296
rect 226706 231104 226762 231160
rect 226614 137944 226670 138000
rect 226890 226072 226946 226128
rect 227074 236680 227130 236736
rect 227166 233960 227222 234016
rect 227258 227024 227314 227080
rect 227166 192616 227222 192672
rect 227258 187176 227314 187232
rect 227074 176160 227130 176216
rect 226982 168000 227038 168056
rect 226890 154264 226946 154320
rect 226798 151544 226854 151600
rect 226706 135224 226762 135280
rect 226522 125432 226578 125488
rect 226522 124208 226578 124264
rect 226522 122712 226578 122768
rect 226522 121488 226578 121544
rect 226522 117136 226578 117192
rect 226522 116048 226578 116104
rect 226522 97824 226578 97880
rect 226522 96872 226578 96928
rect 226522 92384 226578 92440
rect 226522 91432 226578 91488
rect 226522 86808 226578 86864
rect 226522 85992 226578 86048
rect 226522 73072 226578 73128
rect 226522 72256 226578 72312
rect 227718 397976 227774 398032
rect 227442 229744 227498 229800
rect 227534 228384 227590 228440
rect 227626 227160 227682 227216
rect 227534 214512 227590 214568
rect 227442 200776 227498 200832
rect 227626 198056 227682 198112
rect 227350 66816 227406 66872
rect 227626 62056 227682 62112
rect 227626 61376 227682 61432
rect 227810 58928 227866 58984
rect 227718 58520 227774 58576
rect 228546 165280 228602 165336
rect 228454 162560 228510 162616
rect 229006 242256 229062 242312
rect 228914 219952 228970 220008
rect 229006 211792 229062 211848
rect 228822 209072 228878 209128
rect 228730 157120 228786 157176
rect 228638 77696 228694 77752
rect 229282 88712 229338 88768
rect 229558 243480 229614 243536
rect 229466 233824 229522 233880
rect 229374 59744 229430 59800
rect 229742 234640 229798 234696
rect 229742 191800 229798 191856
rect 229558 189896 229614 189952
rect 230754 229880 230810 229936
rect 230662 129648 230718 129704
rect 230938 249192 230994 249248
rect 230938 217232 230994 217288
rect 230846 178880 230902 178936
rect 230754 118768 230810 118824
rect 231306 206352 231362 206408
rect 231214 159840 231270 159896
rect 231122 105032 231178 105088
rect 232042 83136 232098 83192
rect 232134 80416 232190 80472
rect 232410 173440 232466 173496
rect 232318 107752 232374 107808
rect 235998 398112 236054 398168
rect 233422 110608 233478 110664
rect 233330 102312 233386 102368
rect 233238 99592 233294 99648
rect 233514 94152 233570 94208
rect 233974 184456 234030 184512
rect 234066 140664 234122 140720
rect 235262 125432 235318 125488
rect 233882 86808 233938 86864
rect 232502 73072 232558 73128
rect 232226 69536 232282 69592
rect 235538 232056 235594 232112
rect 235446 226344 235502 226400
rect 235630 226616 235686 226672
rect 235630 218048 235686 218104
rect 235538 165688 235594 165744
rect 235446 99456 235502 99512
rect 235354 62056 235410 62112
rect 236182 397296 236238 397352
rect 239218 397296 239274 397352
rect 241610 397296 241666 397352
rect 242898 397296 242954 397352
rect 244462 397296 244518 397352
rect 237378 396752 237434 396808
rect 236642 227976 236698 228032
rect 236734 226480 236790 226536
rect 236734 205672 236790 205728
rect 236642 138080 236698 138136
rect 240138 396752 240194 396808
rect 238114 195336 238170 195392
rect 239402 228112 239458 228168
rect 239402 178064 239458 178120
rect 238206 122712 238262 122768
rect 240782 227840 240838 227896
rect 240874 170992 240930 171048
rect 244370 396752 244426 396808
rect 242438 233280 242494 233336
rect 242346 230288 242402 230344
rect 242254 204176 242310 204232
rect 242162 59608 242218 59664
rect 225418 56616 225474 56672
rect 242438 71848 242494 71904
rect 245658 396752 245714 396808
rect 244370 60152 244426 60208
rect 248602 397296 248658 397352
rect 247130 396772 247186 396808
rect 247130 396752 247132 396772
rect 247132 396752 247184 396772
rect 247184 396752 247186 396772
rect 247682 396636 247738 396672
rect 247682 396616 247684 396636
rect 247684 396616 247736 396636
rect 247736 396616 247738 396636
rect 246302 97824 246358 97880
rect 265162 398112 265218 398168
rect 300858 398112 300914 398168
rect 315762 398112 315818 398168
rect 325698 398112 325754 398168
rect 250074 397296 250130 397352
rect 252650 397296 252706 397352
rect 253570 397296 253626 397352
rect 256146 397296 256202 397352
rect 260930 397296 260986 397352
rect 262034 397296 262090 397352
rect 263598 397296 263654 397352
rect 249890 396752 249946 396808
rect 249154 92384 249210 92440
rect 251270 396752 251326 396808
rect 251178 396616 251234 396672
rect 249890 59880 249946 59936
rect 254490 396752 254546 396808
rect 255318 396752 255374 396808
rect 251270 117136 251326 117192
rect 258078 396888 258134 396944
rect 256698 396752 256754 396808
rect 255318 60016 255374 60072
rect 258170 396752 258226 396808
rect 259458 396752 259514 396808
rect 259550 396616 259606 396672
rect 262218 396752 262274 396808
rect 260102 230560 260158 230616
rect 271142 397296 271198 397352
rect 273258 397296 273314 397352
rect 273626 397296 273682 397352
rect 274730 397296 274786 397352
rect 276386 397296 276442 397352
rect 278042 397296 278098 397352
rect 290186 397296 290242 397352
rect 293314 397296 293370 397352
rect 298466 397296 298522 397352
rect 263874 397160 263930 397216
rect 265254 396772 265310 396808
rect 265254 396752 265256 396772
rect 265256 396752 265308 396772
rect 265308 396752 265310 396772
rect 266450 396752 266506 396808
rect 267830 396752 267886 396808
rect 269118 396752 269174 396808
rect 266358 396616 266414 396672
rect 267738 396616 267794 396672
rect 270590 396752 270646 396808
rect 273442 397160 273498 397216
rect 272522 396772 272578 396808
rect 272522 396752 272524 396772
rect 272524 396752 272576 396772
rect 272576 396752 272578 396772
rect 276110 396752 276166 396808
rect 277490 396752 277546 396808
rect 278778 396752 278834 396808
rect 280158 396752 280214 396808
rect 269762 59472 269818 59528
rect 269118 59336 269174 59392
rect 258078 56888 258134 56944
rect 244922 56752 244978 56808
rect 283562 396772 283618 396808
rect 283562 396752 283564 396772
rect 283564 396752 283616 396772
rect 283616 396752 283618 396772
rect 285954 396752 286010 396808
rect 287058 396752 287114 396808
rect 295338 396752 295394 396808
rect 281998 247016 282054 247072
rect 308586 397316 308642 397352
rect 308586 397296 308588 397316
rect 308588 397296 308640 397316
rect 308640 397296 308642 397316
rect 310978 397296 311034 397352
rect 313370 397296 313426 397352
rect 302238 396752 302294 396808
rect 304998 396752 305054 396808
rect 317418 396752 317474 396808
rect 320178 396752 320234 396808
rect 322938 396752 322994 396808
rect 342258 397296 342314 397352
rect 342350 396752 342406 396808
rect 358818 478896 358874 478952
rect 357438 414296 357494 414352
rect 357530 413072 357586 413128
rect 358910 418784 358966 418840
rect 359002 417152 359058 417208
rect 359094 415792 359150 415848
rect 580170 697176 580226 697232
rect 580170 683848 580226 683904
rect 580170 670692 580172 670712
rect 580172 670692 580224 670712
rect 580224 670692 580226 670712
rect 580170 670656 580226 670692
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 579802 590960 579858 591016
rect 580170 577632 580226 577688
rect 579802 564304 579858 564360
rect 580170 537784 580226 537840
rect 580170 524476 580226 524512
rect 580170 524456 580172 524476
rect 580172 524456 580224 524476
rect 580224 524456 580226 524476
rect 580170 511264 580226 511320
rect 580170 484608 580226 484664
rect 579986 471416 580042 471472
rect 580170 458088 580226 458144
rect 580170 431568 580226 431624
rect 580262 418240 580318 418296
rect 580170 404912 580226 404968
rect 580170 378392 580226 378448
rect 579618 365064 579674 365120
rect 580170 351908 580172 351928
rect 580172 351908 580224 351928
rect 580224 351908 580226 351928
rect 580170 351872 580226 351908
rect 580170 325216 580226 325272
rect 579986 312024 580042 312080
rect 580170 298696 580226 298752
rect 580170 272176 580226 272232
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 357438 237904 357494 237960
rect 396722 227704 396778 227760
rect 580262 226888 580318 226944
rect 579618 152632 579674 152688
rect 580170 125976 580226 126032
rect 580170 59608 580226 59664
rect 356518 58656 356574 58712
rect 347042 57296 347098 57352
rect 429842 57160 429898 57216
rect 368478 5752 368534 5808
rect 383566 5888 383622 5944
rect 394238 6024 394294 6080
rect 397734 6840 397790 6896
rect 408406 3848 408462 3904
rect 411902 3032 411958 3088
rect 415490 3712 415546 3768
rect 418986 3168 419042 3224
rect 422574 3576 422630 3632
rect 426162 6704 426218 6760
rect 429658 3984 429714 4040
rect 433246 6432 433302 6488
rect 436650 6296 436706 6352
rect 443826 3440 443882 3496
rect 465170 3304 465226 3360
rect 472254 6568 472310 6624
rect 579986 46280 580042 46336
rect 580354 225664 580410 225720
rect 580354 86128 580410 86184
rect 580262 33088 580318 33144
rect 580078 19760 580134 19816
rect 565634 5072 565690 5128
rect 572810 4936 572866 4992
rect 576306 4800 576362 4856
rect 580354 6568 580410 6624
rect 582194 6160 582250 6216
<< metal3 >>
rect -960 697220 480 697460
rect 580165 697234 580231 697237
rect 583520 697234 584960 697324
rect 580165 697232 584960 697234
rect 580165 697176 580170 697232
rect 580226 697176 584960 697232
rect 580165 697174 584960 697176
rect 580165 697171 580231 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 2773 684314 2839 684317
rect -960 684312 2839 684314
rect -960 684256 2778 684312
rect 2834 684256 2839 684312
rect -960 684254 2839 684256
rect -960 684164 480 684254
rect 2773 684251 2839 684254
rect 580165 683906 580231 683909
rect 583520 683906 584960 683996
rect 580165 683904 584960 683906
rect 580165 683848 580170 683904
rect 580226 683848 584960 683904
rect 580165 683846 584960 683848
rect 580165 683843 580231 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 3509 671258 3575 671261
rect -960 671256 3575 671258
rect -960 671200 3514 671256
rect 3570 671200 3575 671256
rect -960 671198 3575 671200
rect -960 671108 480 671198
rect 3509 671195 3575 671198
rect 580165 670714 580231 670717
rect 583520 670714 584960 670804
rect 580165 670712 584960 670714
rect 580165 670656 580170 670712
rect 580226 670656 584960 670712
rect 580165 670654 584960 670656
rect 580165 670651 580231 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 3417 658202 3483 658205
rect -960 658200 3483 658202
rect -960 658144 3422 658200
rect 3478 658144 3483 658200
rect -960 658142 3483 658144
rect -960 658052 480 658142
rect 3417 658139 3483 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 3417 632090 3483 632093
rect -960 632088 3483 632090
rect -960 632032 3422 632088
rect 3478 632032 3483 632088
rect -960 632030 3483 632032
rect -960 631940 480 632030
rect 3417 632027 3483 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 3141 619170 3207 619173
rect -960 619168 3207 619170
rect -960 619112 3146 619168
rect 3202 619112 3207 619168
rect -960 619110 3207 619112
rect -960 619020 480 619110
rect 3141 619107 3207 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 3233 606114 3299 606117
rect -960 606112 3299 606114
rect -960 606056 3238 606112
rect 3294 606056 3299 606112
rect -960 606054 3299 606056
rect -960 605964 480 606054
rect 3233 606051 3299 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 579797 591018 579863 591021
rect 583520 591018 584960 591108
rect 579797 591016 584960 591018
rect 579797 590960 579802 591016
rect 579858 590960 584960 591016
rect 579797 590958 584960 590960
rect 579797 590955 579863 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 3325 580002 3391 580005
rect -960 580000 3391 580002
rect -960 579944 3330 580000
rect 3386 579944 3391 580000
rect -960 579942 3391 579944
rect -960 579852 480 579942
rect 3325 579939 3391 579942
rect 580165 577690 580231 577693
rect 583520 577690 584960 577780
rect 580165 577688 584960 577690
rect 580165 577632 580170 577688
rect 580226 577632 584960 577688
rect 580165 577630 584960 577632
rect 580165 577627 580231 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3417 566946 3483 566949
rect -960 566944 3483 566946
rect -960 566888 3422 566944
rect 3478 566888 3483 566944
rect -960 566886 3483 566888
rect -960 566796 480 566886
rect 3417 566883 3483 566886
rect 579797 564362 579863 564365
rect 583520 564362 584960 564452
rect 579797 564360 584960 564362
rect 579797 564304 579802 564360
rect 579858 564304 584960 564360
rect 579797 564302 584960 564304
rect 579797 564299 579863 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 3417 553890 3483 553893
rect -960 553888 3483 553890
rect -960 553832 3422 553888
rect 3478 553832 3483 553888
rect -960 553830 3483 553832
rect -960 553740 480 553830
rect 3417 553827 3483 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 3417 527914 3483 527917
rect -960 527912 3483 527914
rect -960 527856 3422 527912
rect 3478 527856 3483 527912
rect -960 527854 3483 527856
rect -960 527764 480 527854
rect 3417 527851 3483 527854
rect 580165 524514 580231 524517
rect 583520 524514 584960 524604
rect 580165 524512 584960 524514
rect 580165 524456 580170 524512
rect 580226 524456 584960 524512
rect 580165 524454 584960 524456
rect 580165 524451 580231 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 3417 514858 3483 514861
rect -960 514856 3483 514858
rect -960 514800 3422 514856
rect 3478 514800 3483 514856
rect -960 514798 3483 514800
rect -960 514708 480 514798
rect 3417 514795 3483 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 3049 501802 3115 501805
rect -960 501800 3115 501802
rect -960 501744 3054 501800
rect 3110 501744 3115 501800
rect -960 501742 3115 501744
rect -960 501652 480 501742
rect 3049 501739 3115 501742
rect 583520 497844 584960 498084
rect 103973 491466 104039 491469
rect 218646 491466 218652 491468
rect 103973 491464 218652 491466
rect 103973 491408 103978 491464
rect 104034 491408 218652 491464
rect 103973 491406 218652 491408
rect 103973 491403 104039 491406
rect 218646 491404 218652 491406
rect 218716 491404 218722 491468
rect 101673 491330 101739 491333
rect 218830 491330 218836 491332
rect 101673 491328 218836 491330
rect 101673 491272 101678 491328
rect 101734 491272 218836 491328
rect 101673 491270 218836 491272
rect 101673 491267 101739 491270
rect 218830 491268 218836 491270
rect 218900 491268 218906 491332
rect 108757 490242 108823 490245
rect 219198 490242 219204 490244
rect 108757 490240 219204 490242
rect 108757 490184 108762 490240
rect 108818 490184 219204 490240
rect 108757 490182 219204 490184
rect 108757 490179 108823 490182
rect 219198 490180 219204 490182
rect 219268 490180 219274 490244
rect 59077 490106 59143 490109
rect 266077 490106 266143 490109
rect 59077 490104 266143 490106
rect 59077 490048 59082 490104
rect 59138 490048 266082 490104
rect 266138 490048 266143 490104
rect 59077 490046 266143 490048
rect 59077 490043 59143 490046
rect 266077 490043 266143 490046
rect 58709 489970 58775 489973
rect 316033 489970 316099 489973
rect 58709 489968 316099 489970
rect 58709 489912 58714 489968
rect 58770 489912 316038 489968
rect 316094 489912 316099 489968
rect 58709 489910 316099 489912
rect 58709 489907 58775 489910
rect 316033 489907 316099 489910
rect 59169 489018 59235 489021
rect 178309 489018 178375 489021
rect 59169 489016 178375 489018
rect 59169 488960 59174 489016
rect 59230 488960 178314 489016
rect 178370 488960 178375 489016
rect 59169 488958 178375 488960
rect 59169 488955 59235 488958
rect 178309 488955 178375 488958
rect 217777 489018 217843 489021
rect 263593 489018 263659 489021
rect 217777 489016 263659 489018
rect 217777 488960 217782 489016
rect 217838 488960 263598 489016
rect 263654 488960 263659 489016
rect 217777 488958 263659 488960
rect 217777 488955 217843 488958
rect 263593 488955 263659 488958
rect 53649 488882 53715 488885
rect 276197 488882 276263 488885
rect 53649 488880 276263 488882
rect -960 488596 480 488836
rect 53649 488824 53654 488880
rect 53710 488824 276202 488880
rect 276258 488824 276263 488880
rect 53649 488822 276263 488824
rect 53649 488819 53715 488822
rect 276197 488819 276263 488822
rect 58985 488746 59051 488749
rect 301037 488746 301103 488749
rect 58985 488744 301103 488746
rect 58985 488688 58990 488744
rect 59046 488688 301042 488744
rect 301098 488688 301103 488744
rect 58985 488686 301103 488688
rect 58985 488683 59051 488686
rect 301037 488683 301103 488686
rect 58893 488610 58959 488613
rect 303429 488610 303495 488613
rect 58893 488608 303495 488610
rect 58893 488552 58898 488608
rect 58954 488552 303434 488608
rect 303490 488552 303495 488608
rect 58893 488550 303495 488552
rect 58893 488547 58959 488550
rect 303429 488547 303495 488550
rect 55029 487930 55095 487933
rect 130837 487930 130903 487933
rect 55029 487928 130903 487930
rect 55029 487872 55034 487928
rect 55090 487872 130842 487928
rect 130898 487872 130903 487928
rect 55029 487870 130903 487872
rect 55029 487867 55095 487870
rect 130837 487867 130903 487870
rect 99189 487794 99255 487797
rect 196709 487794 196775 487797
rect 99189 487792 196775 487794
rect 99189 487736 99194 487792
rect 99250 487736 196714 487792
rect 196770 487736 196775 487792
rect 99189 487734 196775 487736
rect 99189 487731 99255 487734
rect 196709 487731 196775 487734
rect 126329 487658 126395 487661
rect 202873 487658 202939 487661
rect 126329 487656 202939 487658
rect 126329 487600 126334 487656
rect 126390 487600 202878 487656
rect 202934 487600 202939 487656
rect 126329 487598 202939 487600
rect 126329 487595 126395 487598
rect 202873 487595 202939 487598
rect 217685 487658 217751 487661
rect 256141 487658 256207 487661
rect 217685 487656 256207 487658
rect 217685 487600 217690 487656
rect 217746 487600 256146 487656
rect 256202 487600 256207 487656
rect 217685 487598 256207 487600
rect 217685 487595 217751 487598
rect 256141 487595 256207 487598
rect 54937 487522 55003 487525
rect 145598 487522 145604 487524
rect 54937 487520 145604 487522
rect 54937 487464 54942 487520
rect 54998 487464 145604 487520
rect 54937 487462 145604 487464
rect 54937 487459 55003 487462
rect 145598 487460 145604 487462
rect 145668 487460 145674 487524
rect 217869 487522 217935 487525
rect 271086 487522 271092 487524
rect 217869 487520 271092 487522
rect 217869 487464 217874 487520
rect 217930 487464 271092 487520
rect 217869 487462 271092 487464
rect 217869 487459 217935 487462
rect 271086 487460 271092 487462
rect 271156 487460 271162 487524
rect 56869 487386 56935 487389
rect 318701 487386 318767 487389
rect 56869 487384 318767 487386
rect 56869 487328 56874 487384
rect 56930 487328 318706 487384
rect 318762 487328 318767 487384
rect 56869 487326 318767 487328
rect 56869 487323 56935 487326
rect 318701 487323 318767 487326
rect 53741 487250 53807 487253
rect 111190 487250 111196 487252
rect 53741 487248 111196 487250
rect 53741 487192 53746 487248
rect 53802 487192 111196 487248
rect 53741 487190 111196 487192
rect 53741 487187 53807 487190
rect 111190 487188 111196 487190
rect 111260 487188 111266 487252
rect 217317 487250 217383 487253
rect 340137 487250 340203 487253
rect 217317 487248 340203 487250
rect 217317 487192 217322 487248
rect 217378 487192 340142 487248
rect 340198 487192 340203 487248
rect 217317 487190 340203 487192
rect 217317 487187 217383 487190
rect 340137 487187 340203 487190
rect 90950 487052 90956 487116
rect 91020 487114 91026 487116
rect 217542 487114 217548 487116
rect 91020 487054 217548 487114
rect 91020 487052 91026 487054
rect 217542 487052 217548 487054
rect 217612 487052 217618 487116
rect 138606 486916 138612 486980
rect 138676 486978 138682 486980
rect 197905 486978 197971 486981
rect 138676 486976 197971 486978
rect 138676 486920 197910 486976
rect 197966 486920 197971 486976
rect 138676 486918 197971 486920
rect 138676 486916 138682 486918
rect 197905 486915 197971 486918
rect 218237 486978 218303 486981
rect 326654 486978 326660 486980
rect 218237 486976 326660 486978
rect 218237 486920 218242 486976
rect 218298 486920 326660 486976
rect 218237 486918 326660 486920
rect 218237 486915 218303 486918
rect 326654 486916 326660 486918
rect 326724 486916 326730 486980
rect 150934 486780 150940 486844
rect 151004 486842 151010 486844
rect 217409 486842 217475 486845
rect 151004 486840 217475 486842
rect 151004 486784 217414 486840
rect 217470 486784 217475 486840
rect 151004 486782 217475 486784
rect 151004 486780 151010 486782
rect 217409 486779 217475 486782
rect 218973 486842 219039 486845
rect 266077 486844 266143 486845
rect 248638 486842 248644 486844
rect 218973 486840 248644 486842
rect 218973 486784 218978 486840
rect 219034 486784 248644 486840
rect 218973 486782 248644 486784
rect 218973 486779 219039 486782
rect 248638 486780 248644 486782
rect 248708 486780 248714 486844
rect 266077 486840 266124 486844
rect 266188 486842 266194 486844
rect 266077 486784 266082 486840
rect 266077 486780 266124 486784
rect 266188 486782 266234 486842
rect 266188 486780 266194 486782
rect 266077 486779 266143 486780
rect 126094 486644 126100 486708
rect 126164 486706 126170 486708
rect 126329 486706 126395 486709
rect 126164 486704 126395 486706
rect 126164 486648 126334 486704
rect 126390 486648 126395 486704
rect 126164 486646 126395 486648
rect 126164 486644 126170 486646
rect 126329 486643 126395 486646
rect 130837 486708 130903 486709
rect 130837 486704 130884 486708
rect 130948 486706 130954 486708
rect 130837 486648 130842 486704
rect 130837 486644 130884 486648
rect 130948 486646 130994 486706
rect 130948 486644 130954 486646
rect 143574 486644 143580 486708
rect 143644 486706 143650 486708
rect 198641 486706 198707 486709
rect 143644 486704 198707 486706
rect 143644 486648 198646 486704
rect 198702 486648 198707 486704
rect 143644 486646 198707 486648
rect 143644 486644 143650 486646
rect 130837 486643 130903 486644
rect 198641 486643 198707 486646
rect 218605 486706 218671 486709
rect 283782 486706 283788 486708
rect 218605 486704 283788 486706
rect 218605 486648 218610 486704
rect 218666 486648 283788 486704
rect 218605 486646 283788 486648
rect 218605 486643 218671 486646
rect 283782 486644 283788 486646
rect 283852 486644 283858 486708
rect 101070 486508 101076 486572
rect 101140 486570 101146 486572
rect 101673 486570 101739 486573
rect 101140 486568 101739 486570
rect 101140 486512 101678 486568
rect 101734 486512 101739 486568
rect 101140 486510 101739 486512
rect 101140 486508 101146 486510
rect 101673 486507 101739 486510
rect 103830 486508 103836 486572
rect 103900 486570 103906 486572
rect 103973 486570 104039 486573
rect 103900 486568 104039 486570
rect 103900 486512 103978 486568
rect 104034 486512 104039 486568
rect 103900 486510 104039 486512
rect 103900 486508 103906 486510
rect 103973 486507 104039 486510
rect 108614 486508 108620 486572
rect 108684 486570 108690 486572
rect 108757 486570 108823 486573
rect 108684 486568 108823 486570
rect 108684 486512 108762 486568
rect 108818 486512 108823 486568
rect 108684 486510 108823 486512
rect 108684 486508 108690 486510
rect 108757 486507 108823 486510
rect 123702 486508 123708 486572
rect 123772 486570 123778 486572
rect 202137 486570 202203 486573
rect 123772 486568 202203 486570
rect 123772 486512 202142 486568
rect 202198 486512 202203 486568
rect 123772 486510 202203 486512
rect 123772 486508 123778 486510
rect 202137 486507 202203 486510
rect 219985 486570 220051 486573
rect 288566 486570 288572 486572
rect 219985 486568 288572 486570
rect 219985 486512 219990 486568
rect 220046 486512 288572 486568
rect 219985 486510 288572 486512
rect 219985 486507 220051 486510
rect 288566 486508 288572 486510
rect 288636 486508 288642 486572
rect 316033 486570 316099 486573
rect 315990 486568 316099 486570
rect 315990 486512 316038 486568
rect 316094 486512 316099 486568
rect 315990 486507 316099 486512
rect 315990 486437 316050 486507
rect 116158 486372 116164 486436
rect 116228 486434 116234 486436
rect 198273 486434 198339 486437
rect 116228 486432 198339 486434
rect 116228 486376 198278 486432
rect 198334 486376 198339 486432
rect 116228 486374 198339 486376
rect 116228 486372 116234 486374
rect 198273 486371 198339 486374
rect 218421 486434 218487 486437
rect 305862 486434 305868 486436
rect 218421 486432 305868 486434
rect 218421 486376 218426 486432
rect 218482 486376 305868 486432
rect 218421 486374 305868 486376
rect 218421 486371 218487 486374
rect 305862 486372 305868 486374
rect 305932 486372 305938 486436
rect 315941 486432 316050 486437
rect 315941 486376 315946 486432
rect 316002 486376 316050 486432
rect 315941 486374 316050 486376
rect 318701 486434 318767 486437
rect 339718 486434 339724 486436
rect 318701 486432 339724 486434
rect 318701 486376 318706 486432
rect 318762 486376 339724 486432
rect 318701 486374 339724 486376
rect 315941 486371 316007 486374
rect 318701 486371 318767 486374
rect 339718 486372 339724 486374
rect 339788 486372 339794 486436
rect 340137 486434 340203 486437
rect 350758 486434 350764 486436
rect 340137 486432 350764 486434
rect 340137 486376 340142 486432
rect 340198 486376 350764 486432
rect 340137 486374 350764 486376
rect 340137 486371 340203 486374
rect 350758 486372 350764 486374
rect 350828 486372 350834 486436
rect 118550 486236 118556 486300
rect 118620 486298 118626 486300
rect 203517 486298 203583 486301
rect 118620 486296 203583 486298
rect 118620 486240 203522 486296
rect 203578 486240 203583 486296
rect 118620 486238 203583 486240
rect 118620 486236 118626 486238
rect 203517 486235 203583 486238
rect 219801 486298 219867 486301
rect 313590 486298 313596 486300
rect 219801 486296 313596 486298
rect 219801 486240 219806 486296
rect 219862 486240 313596 486296
rect 219801 486238 313596 486240
rect 219801 486235 219867 486238
rect 313590 486236 313596 486238
rect 313660 486236 313666 486300
rect 106222 486100 106228 486164
rect 106292 486162 106298 486164
rect 198457 486162 198523 486165
rect 106292 486160 198523 486162
rect 106292 486104 198462 486160
rect 198518 486104 198523 486160
rect 106292 486102 198523 486104
rect 106292 486100 106298 486102
rect 198457 486099 198523 486102
rect 219341 486162 219407 486165
rect 318374 486162 318380 486164
rect 219341 486160 318380 486162
rect 219341 486104 219346 486160
rect 219402 486104 318380 486160
rect 219341 486102 318380 486104
rect 219341 486099 219407 486102
rect 318374 486100 318380 486102
rect 318444 486100 318450 486164
rect 56501 486026 56567 486029
rect 93342 486026 93348 486028
rect 56501 486024 93348 486026
rect 56501 485968 56506 486024
rect 56562 485968 93348 486024
rect 56501 485966 93348 485968
rect 56501 485963 56567 485966
rect 93342 485964 93348 485966
rect 93412 485964 93418 486028
rect 98494 485964 98500 486028
rect 98564 486026 98570 486028
rect 99189 486026 99255 486029
rect 98564 486024 99255 486026
rect 98564 485968 99194 486024
rect 99250 485968 99255 486024
rect 98564 485966 99255 485968
rect 98564 485964 98570 485966
rect 99189 485963 99255 485966
rect 114318 485964 114324 486028
rect 114388 486026 114394 486028
rect 218697 486026 218763 486029
rect 114388 486024 218763 486026
rect 114388 485968 218702 486024
rect 218758 485968 218763 486024
rect 114388 485966 218763 485968
rect 114388 485964 114394 485966
rect 218697 485963 218763 485966
rect 219617 486026 219683 486029
rect 323342 486026 323348 486028
rect 219617 486024 323348 486026
rect 219617 485968 219622 486024
rect 219678 485968 323348 486024
rect 219617 485966 323348 485968
rect 219617 485963 219683 485966
rect 323342 485964 323348 485966
rect 323412 485964 323418 486028
rect 88742 485828 88748 485892
rect 88812 485890 88818 485892
rect 88812 485830 156706 485890
rect 88812 485828 88818 485830
rect 156646 485754 156706 485830
rect 158478 485828 158484 485892
rect 158548 485890 158554 485892
rect 198089 485890 198155 485893
rect 158548 485888 198155 485890
rect 158548 485832 198094 485888
rect 198150 485832 198155 485888
rect 158548 485830 198155 485832
rect 158548 485828 158554 485830
rect 198089 485827 198155 485830
rect 217593 485890 217659 485893
rect 256141 485892 256207 485893
rect 263593 485892 263659 485893
rect 253422 485890 253428 485892
rect 217593 485888 253428 485890
rect 217593 485832 217598 485888
rect 217654 485832 253428 485888
rect 217593 485830 253428 485832
rect 217593 485827 217659 485830
rect 253422 485828 253428 485830
rect 253492 485828 253498 485892
rect 256141 485888 256188 485892
rect 256252 485890 256258 485892
rect 263542 485890 263548 485892
rect 256141 485832 256146 485888
rect 256141 485828 256188 485832
rect 256252 485830 256298 485890
rect 263502 485830 263548 485890
rect 263612 485888 263659 485892
rect 263654 485832 263659 485888
rect 256252 485828 256258 485830
rect 263542 485828 263548 485830
rect 263612 485828 263659 485832
rect 256141 485827 256207 485828
rect 263593 485827 263659 485828
rect 276197 485892 276263 485893
rect 303429 485892 303495 485893
rect 276197 485888 276244 485892
rect 276308 485890 276314 485892
rect 276197 485832 276202 485888
rect 276197 485828 276244 485832
rect 276308 485830 276354 485890
rect 303429 485888 303476 485892
rect 303540 485890 303546 485892
rect 303429 485832 303434 485888
rect 276308 485828 276314 485830
rect 303429 485828 303476 485832
rect 303540 485830 303586 485890
rect 303540 485828 303546 485830
rect 338430 485828 338436 485892
rect 338500 485890 338506 485892
rect 356513 485890 356579 485893
rect 338500 485888 356579 485890
rect 338500 485832 356518 485888
rect 356574 485832 356579 485888
rect 338500 485830 356579 485832
rect 338500 485828 338506 485830
rect 276197 485827 276263 485828
rect 303429 485827 303495 485828
rect 356513 485827 356579 485830
rect 156646 485694 161490 485754
rect 161430 485482 161490 485694
rect 166022 485692 166028 485756
rect 166092 485754 166098 485756
rect 219249 485754 219315 485757
rect 166092 485752 219315 485754
rect 166092 485696 219254 485752
rect 219310 485696 219315 485752
rect 166092 485694 219315 485696
rect 166092 485692 166098 485694
rect 219249 485691 219315 485694
rect 178309 485620 178375 485621
rect 178309 485616 178356 485620
rect 178420 485618 178426 485620
rect 198365 485618 198431 485621
rect 260966 485618 260972 485620
rect 178309 485560 178314 485616
rect 178309 485556 178356 485560
rect 178420 485558 178466 485618
rect 198365 485616 260972 485618
rect 198365 485560 198370 485616
rect 198426 485560 260972 485616
rect 198365 485558 260972 485560
rect 178420 485556 178426 485558
rect 178309 485555 178375 485556
rect 198365 485555 198431 485558
rect 260966 485556 260972 485558
rect 261036 485556 261042 485620
rect 219014 485482 219020 485484
rect 161430 485422 219020 485482
rect 219014 485420 219020 485422
rect 219084 485420 219090 485484
rect 136030 485284 136036 485348
rect 136100 485346 136106 485348
rect 209773 485346 209839 485349
rect 136100 485344 209839 485346
rect 136100 485288 209778 485344
rect 209834 485288 209839 485344
rect 136100 485286 209839 485288
rect 136100 485284 136106 485286
rect 209773 485283 209839 485286
rect 216581 485346 216647 485349
rect 216581 485344 296730 485346
rect 216581 485288 216586 485344
rect 216642 485288 296730 485344
rect 216581 485286 296730 485288
rect 216581 485283 216647 485286
rect 59997 485210 60063 485213
rect 88333 485210 88399 485213
rect 59997 485208 88399 485210
rect 59997 485152 60002 485208
rect 60058 485152 88338 485208
rect 88394 485152 88399 485208
rect 59997 485150 88399 485152
rect 59997 485147 60063 485150
rect 88333 485147 88399 485150
rect 128486 485148 128492 485212
rect 128556 485210 128562 485212
rect 218513 485210 218579 485213
rect 128556 485208 218579 485210
rect 128556 485152 218518 485208
rect 218574 485152 218579 485208
rect 128556 485150 218579 485152
rect 128556 485148 128562 485150
rect 218513 485147 218579 485150
rect 219709 485210 219775 485213
rect 251030 485210 251036 485212
rect 219709 485208 251036 485210
rect 219709 485152 219714 485208
rect 219770 485152 251036 485208
rect 219709 485150 251036 485152
rect 219709 485147 219775 485150
rect 251030 485148 251036 485150
rect 251100 485148 251106 485212
rect 296670 485210 296730 485286
rect 308254 485210 308260 485212
rect 296670 485150 308260 485210
rect 308254 485148 308260 485150
rect 308324 485148 308330 485212
rect 58617 485074 58683 485077
rect 104893 485074 104959 485077
rect 58617 485072 104959 485074
rect 58617 485016 58622 485072
rect 58678 485016 104898 485072
rect 104954 485016 104959 485072
rect 58617 485014 104959 485016
rect 58617 485011 58683 485014
rect 104893 485011 104959 485014
rect 120942 485012 120948 485076
rect 121012 485074 121018 485076
rect 218789 485074 218855 485077
rect 301037 485076 301103 485077
rect 121012 485072 218855 485074
rect 121012 485016 218794 485072
rect 218850 485016 218855 485072
rect 121012 485014 218855 485016
rect 121012 485012 121018 485014
rect 218789 485011 218855 485014
rect 219934 485012 219940 485076
rect 220004 485074 220010 485076
rect 295926 485074 295932 485076
rect 220004 485014 295932 485074
rect 220004 485012 220010 485014
rect 295926 485012 295932 485014
rect 295996 485012 296002 485076
rect 301037 485072 301084 485076
rect 301148 485074 301154 485076
rect 301037 485016 301042 485072
rect 301037 485012 301084 485016
rect 301148 485014 301194 485074
rect 301148 485012 301154 485014
rect 301037 485011 301103 485012
rect 55121 484938 55187 484941
rect 268510 484938 268516 484940
rect 55121 484936 268516 484938
rect 55121 484880 55126 484936
rect 55182 484880 268516 484936
rect 55121 484878 268516 484880
rect 55121 484875 55187 484878
rect 268510 484876 268516 484878
rect 268580 484876 268586 484940
rect 53557 484802 53623 484805
rect 278446 484802 278452 484804
rect 53557 484800 278452 484802
rect 53557 484744 53562 484800
rect 53618 484744 278452 484800
rect 53557 484742 278452 484744
rect 53557 484739 53623 484742
rect 278446 484740 278452 484742
rect 278516 484740 278522 484804
rect 53373 484666 53439 484669
rect 311014 484666 311020 484668
rect 53373 484664 311020 484666
rect 53373 484608 53378 484664
rect 53434 484608 311020 484664
rect 53373 484606 311020 484608
rect 53373 484603 53439 484606
rect 311014 484604 311020 484606
rect 311084 484604 311090 484668
rect 580165 484666 580231 484669
rect 583520 484666 584960 484756
rect 580165 484664 584960 484666
rect 580165 484608 580170 484664
rect 580226 484608 584960 484664
rect 580165 484606 584960 484608
rect 580165 484603 580231 484606
rect 59261 484530 59327 484533
rect 179638 484530 179644 484532
rect 59261 484528 179644 484530
rect 59261 484472 59266 484528
rect 59322 484472 179644 484528
rect 59261 484470 179644 484472
rect 59261 484467 59327 484470
rect 179638 484468 179644 484470
rect 179708 484468 179714 484532
rect 190862 484468 190868 484532
rect 190932 484530 190938 484532
rect 217317 484530 217383 484533
rect 190932 484528 217383 484530
rect 190932 484472 217322 484528
rect 217378 484472 217383 484528
rect 190932 484470 217383 484472
rect 190932 484468 190938 484470
rect 217317 484467 217383 484470
rect 218053 484530 218119 484533
rect 298502 484530 298508 484532
rect 218053 484528 298508 484530
rect 218053 484472 218058 484528
rect 218114 484472 298508 484528
rect 218053 484470 298508 484472
rect 218053 484467 218119 484470
rect 298502 484468 298508 484470
rect 298572 484468 298578 484532
rect 583520 484516 584960 484606
rect 57513 484258 57579 484261
rect 219617 484260 219683 484261
rect 155902 484258 155908 484260
rect 57513 484256 155908 484258
rect 57513 484200 57518 484256
rect 57574 484200 155908 484256
rect 57513 484198 155908 484200
rect 57513 484195 57579 484198
rect 155902 484196 155908 484198
rect 155972 484196 155978 484260
rect 219566 484258 219572 484260
rect 219526 484198 219572 484258
rect 219636 484256 219683 484260
rect 219678 484200 219683 484256
rect 219566 484196 219572 484198
rect 219636 484196 219683 484200
rect 219617 484195 219683 484196
rect 59445 484122 59511 484125
rect 161054 484122 161060 484124
rect 59445 484120 161060 484122
rect 59445 484064 59450 484120
rect 59506 484064 161060 484120
rect 59445 484062 161060 484064
rect 59445 484059 59511 484062
rect 161054 484060 161060 484062
rect 161124 484060 161130 484124
rect 219433 484122 219499 484125
rect 273478 484122 273484 484124
rect 219433 484120 273484 484122
rect 219433 484064 219438 484120
rect 219494 484064 273484 484120
rect 219433 484062 273484 484064
rect 219433 484059 219499 484062
rect 273478 484060 273484 484062
rect 273548 484060 273554 484124
rect 56409 483986 56475 483989
rect 163262 483986 163268 483988
rect 56409 483984 163268 483986
rect 56409 483928 56414 483984
rect 56470 483928 163268 483984
rect 56409 483926 163268 483928
rect 56409 483923 56475 483926
rect 163262 483924 163268 483926
rect 163332 483924 163338 483988
rect 198549 483986 198615 483989
rect 258390 483986 258396 483988
rect 198549 483984 258396 483986
rect 198549 483928 198554 483984
rect 198610 483928 258396 483984
rect 198549 483926 258396 483928
rect 198549 483923 198615 483926
rect 258390 483924 258396 483926
rect 258460 483924 258466 483988
rect 133638 483788 133644 483852
rect 133708 483850 133714 483852
rect 219157 483850 219223 483853
rect 133708 483848 219223 483850
rect 133708 483792 219162 483848
rect 219218 483792 219223 483848
rect 133708 483790 219223 483792
rect 133708 483788 133714 483790
rect 219157 483787 219223 483790
rect 219525 483850 219591 483853
rect 280928 483850 280934 483852
rect 219525 483848 280934 483850
rect 219525 483792 219530 483848
rect 219586 483792 280934 483848
rect 219525 483790 280934 483792
rect 219525 483787 219591 483790
rect 280928 483788 280934 483790
rect 280998 483788 281004 483852
rect 315941 483850 316007 483853
rect 316166 483850 316172 483852
rect 315896 483848 316172 483850
rect 315896 483792 315946 483848
rect 316002 483792 316172 483848
rect 315896 483790 316172 483792
rect 315941 483787 316007 483790
rect 316166 483788 316172 483790
rect 316236 483788 316242 483852
rect 122790 483654 142170 483714
rect 96176 483380 96182 483444
rect 96246 483442 96252 483444
rect 122790 483442 122850 483654
rect 96246 483382 122850 483442
rect 96246 483380 96252 483382
rect 141056 483380 141062 483444
rect 141126 483380 141132 483444
rect 142110 483442 142170 483654
rect 153568 483652 153574 483716
rect 153638 483714 153644 483716
rect 218329 483714 218395 483717
rect 153638 483712 218395 483714
rect 153638 483656 218334 483712
rect 218390 483656 218395 483712
rect 153638 483654 218395 483656
rect 153638 483652 153644 483654
rect 218329 483651 218395 483654
rect 219617 483714 219683 483717
rect 286096 483714 286102 483716
rect 219617 483712 286102 483714
rect 219617 483656 219622 483712
rect 219678 483656 286102 483712
rect 219617 483654 286102 483656
rect 219617 483651 219683 483654
rect 286096 483652 286102 483654
rect 286166 483652 286172 483716
rect 148400 483516 148406 483580
rect 148470 483578 148476 483580
rect 218145 483578 218211 483581
rect 148470 483576 218211 483578
rect 148470 483520 218150 483576
rect 218206 483520 218211 483576
rect 148470 483518 218211 483520
rect 148470 483516 148476 483518
rect 218145 483515 218211 483518
rect 219893 483578 219959 483581
rect 290992 483578 290998 483580
rect 219893 483576 290998 483578
rect 219893 483520 219898 483576
rect 219954 483520 290998 483576
rect 219893 483518 290998 483520
rect 219893 483515 219959 483518
rect 290992 483516 290998 483518
rect 291062 483516 291068 483580
rect 196801 483442 196867 483445
rect 142110 483440 196867 483442
rect 142110 483384 196806 483440
rect 196862 483384 196867 483440
rect 142110 483382 196867 483384
rect 141064 483306 141124 483380
rect 196801 483379 196867 483382
rect 219750 483380 219756 483444
rect 219820 483442 219826 483444
rect 293576 483442 293582 483444
rect 219820 483382 293582 483442
rect 219820 483380 219826 483382
rect 293576 483380 293582 483382
rect 293646 483380 293652 483444
rect 321048 483380 321054 483444
rect 321118 483380 321124 483444
rect 218881 483306 218947 483309
rect 141064 483304 218947 483306
rect 141064 483248 218886 483304
rect 218942 483248 218947 483304
rect 141064 483246 218947 483248
rect 218881 483243 218947 483246
rect 219065 483306 219131 483309
rect 321056 483306 321116 483380
rect 219065 483304 321116 483306
rect 219065 483248 219070 483304
rect 219126 483248 321116 483304
rect 219065 483246 321116 483248
rect 219065 483243 219131 483246
rect 218094 480252 218100 480316
rect 218164 480314 218170 480316
rect 219382 480314 219388 480316
rect 218164 480254 219388 480314
rect 218164 480252 218170 480254
rect 219382 480252 219388 480254
rect 219452 480252 219458 480316
rect 218462 479844 218468 479908
rect 218532 479906 218538 479908
rect 219198 479906 219204 479908
rect 218532 479846 219204 479906
rect 218532 479844 218538 479846
rect 219198 479844 219204 479846
rect 219268 479844 219274 479908
rect 197353 479226 197419 479229
rect 196942 479224 197419 479226
rect 196942 479220 197358 479224
rect 196604 479168 197358 479220
rect 197414 479168 197419 479224
rect 196604 479166 197419 479168
rect 196604 479160 197002 479166
rect 197353 479163 197419 479166
rect 356562 478954 356622 479190
rect 358813 478954 358879 478957
rect 356562 478952 358879 478954
rect 356562 478896 358818 478952
rect 358874 478896 358879 478952
rect 356562 478894 358879 478896
rect 358813 478891 358879 478894
rect -960 475690 480 475780
rect 3417 475690 3483 475693
rect -960 475688 3483 475690
rect -960 475632 3422 475688
rect 3478 475632 3483 475688
rect -960 475630 3483 475632
rect -960 475540 480 475630
rect 3417 475627 3483 475630
rect 579981 471474 580047 471477
rect 583520 471474 584960 471564
rect 579981 471472 584960 471474
rect 579981 471416 579986 471472
rect 580042 471416 584960 471472
rect 579981 471414 584960 471416
rect 579981 471411 580047 471414
rect 583520 471324 584960 471414
rect 218462 470732 218468 470796
rect 218532 470794 218538 470796
rect 219198 470794 219204 470796
rect 218532 470734 219204 470794
rect 218532 470732 218538 470734
rect 219198 470732 219204 470734
rect 219268 470732 219274 470796
rect 218462 470460 218468 470524
rect 218532 470522 218538 470524
rect 219382 470522 219388 470524
rect 218532 470462 219388 470522
rect 218532 470460 218538 470462
rect 219382 470460 219388 470462
rect 219452 470460 219458 470524
rect -960 462634 480 462724
rect 3233 462634 3299 462637
rect -960 462632 3299 462634
rect -960 462576 3238 462632
rect 3294 462576 3299 462632
rect -960 462574 3299 462576
rect -960 462484 480 462574
rect 3233 462571 3299 462574
rect 218462 460940 218468 461004
rect 218532 461002 218538 461004
rect 219382 461002 219388 461004
rect 218532 460942 219388 461002
rect 218532 460940 218538 460942
rect 219382 460940 219388 460942
rect 219452 460940 219458 461004
rect 218462 460804 218468 460868
rect 218532 460866 218538 460868
rect 219382 460866 219388 460868
rect 218532 460806 219388 460866
rect 218532 460804 218538 460806
rect 219382 460804 219388 460806
rect 219452 460804 219458 460868
rect 580165 458146 580231 458149
rect 583520 458146 584960 458236
rect 580165 458144 584960 458146
rect 580165 458088 580170 458144
rect 580226 458088 584960 458144
rect 580165 458086 584960 458088
rect 580165 458083 580231 458086
rect 583520 457996 584960 458086
rect 218462 451284 218468 451348
rect 218532 451346 218538 451348
rect 219382 451346 219388 451348
rect 218532 451286 219388 451346
rect 218532 451284 218538 451286
rect 219382 451284 219388 451286
rect 219452 451284 219458 451348
rect 218462 451148 218468 451212
rect 218532 451210 218538 451212
rect 219382 451210 219388 451212
rect 218532 451150 219388 451210
rect 218532 451148 218538 451150
rect 219382 451148 219388 451150
rect 219452 451148 219458 451212
rect -960 449578 480 449668
rect 3141 449578 3207 449581
rect -960 449576 3207 449578
rect -960 449520 3146 449576
rect 3202 449520 3207 449576
rect -960 449518 3207 449520
rect -960 449428 480 449518
rect 3141 449515 3207 449518
rect 583520 444668 584960 444908
rect 218462 441628 218468 441692
rect 218532 441690 218538 441692
rect 219382 441690 219388 441692
rect 218532 441630 219388 441690
rect 218532 441628 218538 441630
rect 219382 441628 219388 441630
rect 219452 441628 219458 441692
rect 218462 441492 218468 441556
rect 218532 441554 218538 441556
rect 219382 441554 219388 441556
rect 218532 441494 219388 441554
rect 218532 441492 218538 441494
rect 219382 441492 219388 441494
rect 219452 441492 219458 441556
rect 217961 436930 218027 436933
rect 217961 436928 219450 436930
rect -960 436508 480 436748
rect 57605 436386 57671 436389
rect 60002 436386 60062 436894
rect 217961 436872 217966 436928
rect 218022 436924 219450 436928
rect 218022 436872 220064 436924
rect 217961 436870 220064 436872
rect 217961 436867 218027 436870
rect 219390 436864 220064 436870
rect 57605 436384 60062 436386
rect 57605 436328 57610 436384
rect 57666 436328 60062 436384
rect 57605 436326 60062 436328
rect 57605 436323 57671 436326
rect 216673 435978 216739 435981
rect 216673 435976 219450 435978
rect 56685 435434 56751 435437
rect 60002 435434 60062 435942
rect 216673 435920 216678 435976
rect 216734 435972 219450 435976
rect 216734 435920 220064 435972
rect 216673 435918 220064 435920
rect 216673 435915 216739 435918
rect 219390 435912 220064 435918
rect 56685 435432 60062 435434
rect 56685 435376 56690 435432
rect 56746 435376 60062 435432
rect 56685 435374 60062 435376
rect 56685 435371 56751 435374
rect 216673 433802 216739 433805
rect 216673 433800 219450 433802
rect 57697 433394 57763 433397
rect 60002 433394 60062 433766
rect 216673 433744 216678 433800
rect 216734 433796 219450 433800
rect 216734 433744 220064 433796
rect 216673 433742 220064 433744
rect 216673 433739 216739 433742
rect 219390 433736 220064 433742
rect 57697 433392 60062 433394
rect 57697 433336 57702 433392
rect 57758 433336 60062 433392
rect 57697 433334 60062 433336
rect 57697 433331 57763 433334
rect 216673 432850 216739 432853
rect 216673 432848 219450 432850
rect 57421 432442 57487 432445
rect 60002 432442 60062 432814
rect 216673 432792 216678 432848
rect 216734 432844 219450 432848
rect 216734 432792 220064 432844
rect 216673 432790 220064 432792
rect 216673 432787 216739 432790
rect 219390 432784 220064 432790
rect 57421 432440 60062 432442
rect 57421 432384 57426 432440
rect 57482 432384 60062 432440
rect 57421 432382 60062 432384
rect 57421 432379 57487 432382
rect 218462 431972 218468 432036
rect 218532 432034 218538 432036
rect 219382 432034 219388 432036
rect 218532 431974 219388 432034
rect 218532 431972 218538 431974
rect 219382 431972 219388 431974
rect 219452 431972 219458 432036
rect 218462 431836 218468 431900
rect 218532 431898 218538 431900
rect 219382 431898 219388 431900
rect 218532 431838 219388 431898
rect 218532 431836 218538 431838
rect 219382 431836 219388 431838
rect 219452 431836 219458 431900
rect 580165 431626 580231 431629
rect 583520 431626 584960 431716
rect 580165 431624 584960 431626
rect 580165 431568 580170 431624
rect 580226 431568 584960 431624
rect 580165 431566 584960 431568
rect 580165 431563 580231 431566
rect 583520 431476 584960 431566
rect 217501 431082 217567 431085
rect 217501 431080 219450 431082
rect 57329 430674 57395 430677
rect 60002 430674 60062 431046
rect 217501 431024 217506 431080
rect 217562 431076 219450 431080
rect 217562 431024 220064 431076
rect 217501 431022 220064 431024
rect 217501 431019 217567 431022
rect 219390 431016 220064 431022
rect 57329 430672 60062 430674
rect 57329 430616 57334 430672
rect 57390 430616 60062 430672
rect 57329 430614 60062 430616
rect 57329 430611 57395 430614
rect 216673 429994 216739 429997
rect 216673 429992 219450 429994
rect 57237 429450 57303 429453
rect 60002 429450 60062 429958
rect 216673 429936 216678 429992
rect 216734 429988 219450 429992
rect 216734 429936 220064 429988
rect 216673 429934 220064 429936
rect 216673 429931 216739 429934
rect 219390 429928 220064 429934
rect 57237 429448 60062 429450
rect 57237 429392 57242 429448
rect 57298 429392 60062 429448
rect 57237 429390 60062 429392
rect 57237 429387 57303 429390
rect 217225 428226 217291 428229
rect 217225 428224 219450 428226
rect 57881 427954 57947 427957
rect 60002 427954 60062 428190
rect 217225 428168 217230 428224
rect 217286 428220 219450 428224
rect 217286 428168 220064 428220
rect 217225 428166 220064 428168
rect 217225 428163 217291 428166
rect 219390 428160 220064 428166
rect 57881 427952 60062 427954
rect 57881 427896 57886 427952
rect 57942 427896 60062 427952
rect 57881 427894 60062 427896
rect 57881 427891 57947 427894
rect -960 423602 480 423692
rect 3417 423602 3483 423605
rect -960 423600 3483 423602
rect -960 423544 3422 423600
rect 3478 423544 3483 423600
rect -960 423542 3483 423544
rect -960 423452 480 423542
rect 3417 423539 3483 423542
rect 218462 422316 218468 422380
rect 218532 422378 218538 422380
rect 219382 422378 219388 422380
rect 218532 422318 219388 422378
rect 218532 422316 218538 422318
rect 219382 422316 219388 422318
rect 219452 422316 219458 422380
rect 218462 422180 218468 422244
rect 218532 422242 218538 422244
rect 219382 422242 219388 422244
rect 218532 422182 219388 422242
rect 218532 422180 218538 422182
rect 219382 422180 219388 422182
rect 219452 422180 219458 422244
rect 198825 419386 198891 419389
rect 197126 419384 198891 419386
rect 197126 419380 198830 419384
rect 196604 419328 198830 419380
rect 198886 419328 198891 419384
rect 196604 419326 198891 419328
rect 196604 419320 197186 419326
rect 198825 419323 198891 419326
rect 356562 418842 356622 419350
rect 358905 418842 358971 418845
rect 356562 418840 358971 418842
rect 356562 418784 358910 418840
rect 358966 418784 358971 418840
rect 356562 418782 358971 418784
rect 358905 418779 358971 418782
rect 580257 418298 580323 418301
rect 583520 418298 584960 418388
rect 580257 418296 584960 418298
rect 580257 418240 580262 418296
rect 580318 418240 584960 418296
rect 580257 418238 584960 418240
rect 580257 418235 580323 418238
rect 583520 418148 584960 418238
rect 198733 417754 198799 417757
rect 197126 417752 198799 417754
rect 197126 417748 198738 417752
rect 196604 417696 198738 417748
rect 198794 417696 198799 417752
rect 196604 417694 198799 417696
rect 196604 417688 197186 417694
rect 198733 417691 198799 417694
rect 356562 417210 356622 417718
rect 358997 417210 359063 417213
rect 356562 417208 359063 417210
rect 356562 417152 359002 417208
rect 359058 417152 359063 417208
rect 356562 417150 359063 417152
rect 358997 417147 359063 417150
rect 199009 416394 199075 416397
rect 197126 416392 199075 416394
rect 197126 416388 199014 416392
rect 196604 416336 199014 416388
rect 199070 416336 199075 416392
rect 196604 416334 199075 416336
rect 196604 416328 197186 416334
rect 199009 416331 199075 416334
rect 356562 415850 356622 416358
rect 359089 415850 359155 415853
rect 356562 415848 359155 415850
rect 356562 415792 359094 415848
rect 359150 415792 359155 415848
rect 356562 415790 359155 415792
rect 359089 415787 359155 415790
rect 199377 414898 199443 414901
rect 197126 414896 199443 414898
rect 197126 414892 199382 414896
rect 196604 414840 199382 414892
rect 199438 414840 199443 414896
rect 196604 414838 199443 414840
rect 196604 414832 197186 414838
rect 199377 414835 199443 414838
rect 356562 414354 356622 414862
rect 357433 414354 357499 414357
rect 356562 414352 357499 414354
rect 356562 414296 357438 414352
rect 357494 414296 357499 414352
rect 356562 414294 357499 414296
rect 357433 414291 357499 414294
rect 198917 413674 198983 413677
rect 197126 413672 198983 413674
rect 197126 413668 198922 413672
rect 196604 413616 198922 413668
rect 198978 413616 198983 413672
rect 196604 413614 198983 413616
rect 196604 413608 197186 413614
rect 198917 413611 198983 413614
rect 356562 413130 356622 413638
rect 357525 413130 357591 413133
rect 356562 413128 357591 413130
rect 356562 413072 357530 413128
rect 357586 413072 357591 413128
rect 356562 413070 357591 413072
rect 357525 413067 357591 413070
rect 218462 412660 218468 412724
rect 218532 412722 218538 412724
rect 219382 412722 219388 412724
rect 218532 412662 219388 412722
rect 218532 412660 218538 412662
rect 219382 412660 219388 412662
rect 219452 412660 219458 412724
rect 218462 412524 218468 412588
rect 218532 412586 218538 412588
rect 219382 412586 219388 412588
rect 218532 412526 219388 412586
rect 218532 412524 218538 412526
rect 219382 412524 219388 412526
rect 219452 412524 219458 412588
rect -960 410546 480 410636
rect 3141 410546 3207 410549
rect -960 410544 3207 410546
rect -960 410488 3146 410544
rect 3202 410488 3207 410544
rect -960 410486 3207 410488
rect -960 410396 480 410486
rect 3141 410483 3207 410486
rect 57789 410002 57855 410005
rect 216673 410002 216739 410005
rect 57789 410000 60062 410002
rect 57789 409944 57794 410000
rect 57850 409944 60062 410000
rect 57789 409942 60062 409944
rect 216673 410000 219450 410002
rect 216673 409944 216678 410000
rect 216734 409996 219450 410000
rect 216734 409944 220064 409996
rect 216673 409942 220064 409944
rect 57789 409939 57855 409942
rect 216673 409939 216739 409942
rect 219390 409936 220064 409942
rect 217317 408370 217383 408373
rect 217317 408368 219450 408370
rect 59353 408234 59419 408237
rect 60002 408234 60062 408334
rect 217317 408312 217322 408368
rect 217378 408364 219450 408368
rect 217378 408312 220064 408364
rect 217317 408310 220064 408312
rect 217317 408307 217383 408310
rect 219390 408304 220064 408310
rect 59353 408232 60062 408234
rect 59353 408176 59358 408232
rect 59414 408176 60062 408232
rect 59353 408174 60062 408176
rect 59353 408171 59419 408174
rect 217133 408098 217199 408101
rect 217133 408096 220094 408098
rect 56593 407554 56659 407557
rect 60002 407554 60062 408062
rect 217133 408040 217138 408096
rect 217194 408040 220094 408096
rect 217133 408038 220094 408040
rect 217133 408035 217199 408038
rect 56593 407552 60062 407554
rect 56593 407496 56598 407552
rect 56654 407496 60062 407552
rect 56593 407494 60062 407496
rect 56593 407491 56659 407494
rect 580165 404970 580231 404973
rect 583520 404970 584960 405060
rect 580165 404968 584960 404970
rect 580165 404912 580170 404968
rect 580226 404912 584960 404968
rect 580165 404910 584960 404912
rect 580165 404907 580231 404910
rect 583520 404820 584960 404910
rect 219566 403276 219572 403340
rect 219636 403338 219642 403340
rect 219636 403278 220002 403338
rect 219636 403276 219642 403278
rect 219566 403140 219572 403204
rect 219636 403202 219642 403204
rect 219709 403202 219775 403205
rect 219636 403200 219775 403202
rect 219636 403144 219714 403200
rect 219770 403144 219775 403200
rect 219636 403142 219775 403144
rect 219636 403140 219642 403142
rect 219709 403139 219775 403142
rect 218462 403004 218468 403068
rect 218532 403066 218538 403068
rect 219382 403066 219388 403068
rect 218532 403006 219388 403066
rect 218532 403004 218538 403006
rect 219382 403004 219388 403006
rect 219452 403004 219458 403068
rect 219942 402933 220002 403278
rect 218462 402868 218468 402932
rect 218532 402930 218538 402932
rect 219382 402930 219388 402932
rect 218532 402870 219388 402930
rect 218532 402868 218538 402870
rect 219382 402868 219388 402870
rect 219452 402868 219458 402932
rect 219893 402928 220002 402933
rect 219893 402872 219898 402928
rect 219954 402872 220002 402928
rect 219893 402870 220002 402872
rect 219893 402867 219959 402870
rect 219566 399876 219572 399940
rect 219636 399938 219642 399940
rect 220077 399938 220143 399941
rect 219636 399936 220143 399938
rect 219636 399880 220082 399936
rect 220138 399880 220143 399936
rect 219636 399878 220143 399880
rect 219636 399876 219642 399878
rect 220077 399875 220143 399878
rect 96040 399604 96046 399668
rect 96110 399666 96116 399668
rect 96470 399666 96476 399668
rect 96110 399606 96476 399666
rect 96110 399604 96116 399606
rect 96470 399604 96476 399606
rect 96540 399604 96546 399668
rect 218237 399530 218303 399533
rect 223614 399530 223620 399532
rect 218237 399528 223620 399530
rect 218237 399472 218242 399528
rect 218298 399472 223620 399528
rect 218237 399470 223620 399472
rect 218237 399467 218303 399470
rect 223614 399468 223620 399470
rect 223684 399468 223690 399532
rect 218462 398244 218468 398308
rect 218532 398306 218538 398308
rect 218605 398306 218671 398309
rect 226374 398306 226380 398308
rect 218532 398304 218671 398306
rect 218532 398248 218610 398304
rect 218666 398248 218671 398304
rect 218532 398246 218671 398248
rect 218532 398244 218538 398246
rect 218605 398243 218671 398246
rect 219390 398246 226380 398306
rect 85389 398172 85455 398173
rect 113633 398172 113699 398173
rect 85389 398168 85436 398172
rect 85500 398170 85506 398172
rect 113582 398170 113588 398172
rect 85389 398112 85394 398168
rect 85389 398108 85436 398112
rect 85500 398110 85546 398170
rect 113542 398110 113588 398170
rect 113652 398168 113699 398172
rect 113694 398112 113699 398168
rect 85500 398108 85506 398110
rect 113582 398108 113588 398110
rect 113652 398108 113699 398112
rect 85389 398107 85455 398108
rect 113633 398107 113699 398108
rect 217869 398170 217935 398173
rect 219390 398170 219450 398246
rect 226374 398244 226380 398246
rect 226444 398244 226450 398308
rect 235993 398172 236059 398173
rect 217869 398168 219450 398170
rect 217869 398112 217874 398168
rect 217930 398112 219450 398168
rect 217869 398110 219450 398112
rect 217869 398107 217935 398110
rect 219934 398108 219940 398172
rect 220004 398170 220010 398172
rect 227846 398170 227852 398172
rect 220004 398110 227852 398170
rect 220004 398108 220010 398110
rect 227846 398108 227852 398110
rect 227916 398108 227922 398172
rect 235942 398170 235948 398172
rect 235902 398110 235948 398170
rect 236012 398168 236059 398172
rect 236054 398112 236059 398168
rect 235942 398108 235948 398110
rect 236012 398108 236059 398112
rect 235993 398107 236059 398108
rect 265157 398172 265223 398173
rect 300853 398172 300919 398173
rect 315757 398172 315823 398173
rect 265157 398168 265204 398172
rect 265268 398170 265274 398172
rect 265157 398112 265162 398168
rect 265157 398108 265204 398112
rect 265268 398110 265314 398170
rect 300853 398168 300900 398172
rect 300964 398170 300970 398172
rect 300853 398112 300858 398168
rect 265268 398108 265274 398110
rect 300853 398108 300900 398112
rect 300964 398110 301010 398170
rect 315757 398168 315804 398172
rect 315868 398170 315874 398172
rect 325693 398170 325759 398173
rect 325918 398170 325924 398172
rect 315757 398112 315762 398168
rect 300964 398108 300970 398110
rect 315757 398108 315804 398112
rect 315868 398110 315914 398170
rect 325693 398168 325924 398170
rect 325693 398112 325698 398168
rect 325754 398112 325924 398168
rect 325693 398110 325924 398112
rect 315868 398108 315874 398110
rect 265157 398107 265223 398108
rect 300853 398107 300919 398108
rect 315757 398107 315823 398108
rect 325693 398107 325759 398110
rect 325918 398108 325924 398110
rect 325988 398108 325994 398172
rect 218053 398034 218119 398037
rect 218053 398032 219450 398034
rect 218053 397976 218058 398032
rect 218114 397976 219450 398032
rect 218053 397974 219450 397976
rect 218053 397971 218119 397974
rect 219390 397898 219450 397974
rect 219750 397972 219756 398036
rect 219820 398034 219826 398036
rect 227713 398034 227779 398037
rect 219820 398032 227779 398034
rect 219820 397976 227718 398032
rect 227774 397976 227779 398032
rect 219820 397974 227779 397976
rect 219820 397972 219826 397974
rect 227713 397971 227779 397974
rect 227662 397898 227668 397900
rect 219390 397838 227668 397898
rect 227662 397836 227668 397838
rect 227732 397836 227738 397900
rect -960 397490 480 397580
rect 3417 397490 3483 397493
rect -960 397488 3483 397490
rect -960 397432 3422 397488
rect 3478 397432 3483 397488
rect -960 397430 3483 397432
rect -960 397340 480 397430
rect 3417 397427 3483 397430
rect 78305 397356 78371 397357
rect 78254 397354 78260 397356
rect 78214 397294 78260 397354
rect 78324 397352 78371 397356
rect 78366 397296 78371 397352
rect 78254 397292 78260 397294
rect 78324 397292 78371 397296
rect 79542 397292 79548 397356
rect 79612 397354 79618 397356
rect 79961 397354 80027 397357
rect 79612 397352 80027 397354
rect 79612 397296 79966 397352
rect 80022 397296 80027 397352
rect 79612 397294 80027 397296
rect 79612 397292 79618 397294
rect 78305 397291 78371 397292
rect 79961 397291 80027 397294
rect 80421 397356 80487 397357
rect 83273 397356 83339 397357
rect 80421 397352 80468 397356
rect 80532 397354 80538 397356
rect 83222 397354 83228 397356
rect 80421 397296 80426 397352
rect 80421 397292 80468 397296
rect 80532 397294 80578 397354
rect 83182 397294 83228 397354
rect 83292 397352 83339 397356
rect 83334 397296 83339 397352
rect 80532 397292 80538 397294
rect 83222 397292 83228 397294
rect 83292 397292 83339 397296
rect 80421 397291 80487 397292
rect 83273 397291 83339 397292
rect 86493 397356 86559 397357
rect 87689 397356 87755 397357
rect 86493 397352 86540 397356
rect 86604 397354 86610 397356
rect 87638 397354 87644 397356
rect 86493 397296 86498 397352
rect 86493 397292 86540 397296
rect 86604 397294 86650 397354
rect 87598 397294 87644 397354
rect 87708 397352 87755 397356
rect 87750 397296 87755 397352
rect 86604 397292 86610 397294
rect 87638 397292 87644 397294
rect 87708 397292 87755 397296
rect 86493 397291 86559 397292
rect 87689 397291 87755 397292
rect 88701 397356 88767 397357
rect 88701 397352 88748 397356
rect 88812 397354 88818 397356
rect 88701 397296 88706 397352
rect 88701 397292 88748 397296
rect 88812 397294 88858 397354
rect 88812 397292 88818 397294
rect 91318 397292 91324 397356
rect 91388 397354 91394 397356
rect 92289 397354 92355 397357
rect 91388 397352 92355 397354
rect 91388 397296 92294 397352
rect 92350 397296 92355 397352
rect 91388 397294 92355 397296
rect 91388 397292 91394 397294
rect 88701 397291 88767 397292
rect 92289 397291 92355 397294
rect 93342 397292 93348 397356
rect 93412 397354 93418 397356
rect 93485 397354 93551 397357
rect 93412 397352 93551 397354
rect 93412 397296 93490 397352
rect 93546 397296 93551 397352
rect 93412 397294 93551 397296
rect 93412 397292 93418 397294
rect 93485 397291 93551 397294
rect 96286 397292 96292 397356
rect 96356 397354 96362 397356
rect 96521 397354 96587 397357
rect 96356 397352 96587 397354
rect 96356 397296 96526 397352
rect 96582 397296 96587 397352
rect 96356 397294 96587 397296
rect 96356 397292 96362 397294
rect 96521 397291 96587 397294
rect 98126 397292 98132 397356
rect 98196 397354 98202 397356
rect 98913 397354 98979 397357
rect 98196 397352 98979 397354
rect 98196 397296 98918 397352
rect 98974 397296 98979 397352
rect 98196 397294 98979 397296
rect 98196 397292 98202 397294
rect 98913 397291 98979 397294
rect 99966 397292 99972 397356
rect 100036 397354 100042 397356
rect 100109 397354 100175 397357
rect 100036 397352 100175 397354
rect 100036 397296 100114 397352
rect 100170 397296 100175 397352
rect 100036 397294 100175 397296
rect 100036 397292 100042 397294
rect 100109 397291 100175 397294
rect 100702 397292 100708 397356
rect 100772 397354 100778 397356
rect 101581 397354 101647 397357
rect 101857 397356 101923 397357
rect 101806 397354 101812 397356
rect 100772 397352 101647 397354
rect 100772 397296 101586 397352
rect 101642 397296 101647 397352
rect 100772 397294 101647 397296
rect 101766 397294 101812 397354
rect 101876 397352 101923 397356
rect 101918 397296 101923 397352
rect 100772 397292 100778 397294
rect 101581 397291 101647 397294
rect 101806 397292 101812 397294
rect 101876 397292 101923 397296
rect 102726 397292 102732 397356
rect 102796 397354 102802 397356
rect 102869 397354 102935 397357
rect 102796 397352 102935 397354
rect 102796 397296 102874 397352
rect 102930 397296 102935 397352
rect 102796 397294 102935 397296
rect 102796 397292 102802 397294
rect 101857 397291 101923 397292
rect 102869 397291 102935 397294
rect 103697 397354 103763 397357
rect 103830 397354 103836 397356
rect 103697 397352 103836 397354
rect 103697 397296 103702 397352
rect 103758 397296 103836 397352
rect 103697 397294 103836 397296
rect 103697 397291 103763 397294
rect 103830 397292 103836 397294
rect 103900 397292 103906 397356
rect 105302 397292 105308 397356
rect 105372 397354 105378 397356
rect 105905 397354 105971 397357
rect 105372 397352 105971 397354
rect 105372 397296 105910 397352
rect 105966 397296 105971 397352
rect 105372 397294 105971 397296
rect 105372 397292 105378 397294
rect 105905 397291 105971 397294
rect 106406 397292 106412 397356
rect 106476 397354 106482 397356
rect 107193 397354 107259 397357
rect 106476 397352 107259 397354
rect 106476 397296 107198 397352
rect 107254 397296 107259 397352
rect 106476 397294 107259 397296
rect 106476 397292 106482 397294
rect 107193 397291 107259 397294
rect 109534 397292 109540 397356
rect 109604 397354 109610 397356
rect 109769 397354 109835 397357
rect 109604 397352 109835 397354
rect 109604 397296 109774 397352
rect 109830 397296 109835 397352
rect 109604 397294 109835 397296
rect 109604 397292 109610 397294
rect 109769 397291 109835 397294
rect 111190 397292 111196 397356
rect 111260 397354 111266 397356
rect 111609 397354 111675 397357
rect 111260 397352 111675 397354
rect 111260 397296 111614 397352
rect 111670 397296 111675 397352
rect 111260 397294 111675 397296
rect 111260 397292 111266 397294
rect 111609 397291 111675 397294
rect 114461 397356 114527 397357
rect 115841 397356 115907 397357
rect 114461 397352 114508 397356
rect 114572 397354 114578 397356
rect 115790 397354 115796 397356
rect 114461 397296 114466 397352
rect 114461 397292 114508 397296
rect 114572 397294 114618 397354
rect 115750 397294 115796 397354
rect 115860 397352 115907 397356
rect 115902 397296 115907 397352
rect 114572 397292 114578 397294
rect 115790 397292 115796 397294
rect 115860 397292 115907 397296
rect 114461 397291 114527 397292
rect 115841 397291 115907 397292
rect 118141 397354 118207 397357
rect 118366 397354 118372 397356
rect 118141 397352 118372 397354
rect 118141 397296 118146 397352
rect 118202 397296 118372 397352
rect 118141 397294 118372 397296
rect 118141 397291 118207 397294
rect 118366 397292 118372 397294
rect 118436 397292 118442 397356
rect 136030 397292 136036 397356
rect 136100 397354 136106 397356
rect 136449 397354 136515 397357
rect 138473 397356 138539 397357
rect 138422 397354 138428 397356
rect 136100 397352 136515 397354
rect 136100 397296 136454 397352
rect 136510 397296 136515 397352
rect 136100 397294 136515 397296
rect 138382 397294 138428 397354
rect 138492 397352 138539 397356
rect 138534 397296 138539 397352
rect 136100 397292 136106 397294
rect 136449 397291 136515 397294
rect 138422 397292 138428 397294
rect 138492 397292 138539 397296
rect 138473 397291 138539 397292
rect 150709 397354 150775 397357
rect 183461 397356 183527 397357
rect 150934 397354 150940 397356
rect 150709 397352 150940 397354
rect 150709 397296 150714 397352
rect 150770 397296 150940 397352
rect 150709 397294 150940 397296
rect 150709 397291 150775 397294
rect 150934 397292 150940 397294
rect 151004 397292 151010 397356
rect 183461 397352 183508 397356
rect 183572 397354 183578 397356
rect 236177 397354 236243 397357
rect 239213 397356 239279 397357
rect 241605 397356 241671 397357
rect 242893 397356 242959 397357
rect 237046 397354 237052 397356
rect 183461 397296 183466 397352
rect 183461 397292 183508 397296
rect 183572 397294 183618 397354
rect 236177 397352 237052 397354
rect 236177 397296 236182 397352
rect 236238 397296 237052 397352
rect 236177 397294 237052 397296
rect 183572 397292 183578 397294
rect 183461 397291 183527 397292
rect 236177 397291 236243 397294
rect 237046 397292 237052 397294
rect 237116 397292 237122 397356
rect 239213 397352 239260 397356
rect 239324 397354 239330 397356
rect 239213 397296 239218 397352
rect 239213 397292 239260 397296
rect 239324 397294 239370 397354
rect 241605 397352 241652 397356
rect 241716 397354 241722 397356
rect 241605 397296 241610 397352
rect 239324 397292 239330 397294
rect 241605 397292 241652 397296
rect 241716 397294 241762 397354
rect 242893 397352 242940 397356
rect 243004 397354 243010 397356
rect 244457 397354 244523 397357
rect 248597 397356 248663 397357
rect 245326 397354 245332 397356
rect 242893 397296 242898 397352
rect 241716 397292 241722 397294
rect 242893 397292 242940 397296
rect 243004 397294 243050 397354
rect 244457 397352 245332 397354
rect 244457 397296 244462 397352
rect 244518 397296 245332 397352
rect 244457 397294 245332 397296
rect 243004 397292 243010 397294
rect 239213 397291 239279 397292
rect 241605 397291 241671 397292
rect 242893 397291 242959 397292
rect 244457 397291 244523 397294
rect 245326 397292 245332 397294
rect 245396 397292 245402 397356
rect 248597 397352 248644 397356
rect 248708 397354 248714 397356
rect 250069 397354 250135 397357
rect 250662 397354 250668 397356
rect 248597 397296 248602 397352
rect 248597 397292 248644 397296
rect 248708 397294 248754 397354
rect 250069 397352 250668 397354
rect 250069 397296 250074 397352
rect 250130 397296 250668 397352
rect 250069 397294 250668 397296
rect 248708 397292 248714 397294
rect 248597 397291 248663 397292
rect 250069 397291 250135 397294
rect 250662 397292 250668 397294
rect 250732 397292 250738 397356
rect 252645 397354 252711 397357
rect 253565 397356 253631 397357
rect 256141 397356 256207 397357
rect 260925 397356 260991 397357
rect 262029 397356 262095 397357
rect 263593 397356 263659 397357
rect 253422 397354 253428 397356
rect 252645 397352 253428 397354
rect 252645 397296 252650 397352
rect 252706 397296 253428 397352
rect 252645 397294 253428 397296
rect 252645 397291 252711 397294
rect 253422 397292 253428 397294
rect 253492 397292 253498 397356
rect 253565 397352 253612 397356
rect 253676 397354 253682 397356
rect 253565 397296 253570 397352
rect 253565 397292 253612 397296
rect 253676 397294 253722 397354
rect 256141 397352 256188 397356
rect 256252 397354 256258 397356
rect 256141 397296 256146 397352
rect 253676 397292 253682 397294
rect 256141 397292 256188 397296
rect 256252 397294 256298 397354
rect 260925 397352 260972 397356
rect 261036 397354 261042 397356
rect 260925 397296 260930 397352
rect 256252 397292 256258 397294
rect 260925 397292 260972 397296
rect 261036 397294 261082 397354
rect 262029 397352 262076 397356
rect 262140 397354 262146 397356
rect 263542 397354 263548 397356
rect 262029 397296 262034 397352
rect 261036 397292 261042 397294
rect 262029 397292 262076 397296
rect 262140 397294 262186 397354
rect 263502 397294 263548 397354
rect 263612 397352 263659 397356
rect 263654 397296 263659 397352
rect 262140 397292 262146 397294
rect 263542 397292 263548 397294
rect 263612 397292 263659 397296
rect 253565 397291 253631 397292
rect 256141 397291 256207 397292
rect 260925 397291 260991 397292
rect 262029 397291 262095 397292
rect 263593 397291 263659 397292
rect 271137 397354 271203 397357
rect 273253 397356 273319 397357
rect 271270 397354 271276 397356
rect 271137 397352 271276 397354
rect 271137 397296 271142 397352
rect 271198 397296 271276 397352
rect 271137 397294 271276 397296
rect 271137 397291 271203 397294
rect 271270 397292 271276 397294
rect 271340 397292 271346 397356
rect 273253 397352 273300 397356
rect 273364 397354 273370 397356
rect 273621 397354 273687 397357
rect 274398 397354 274404 397356
rect 273253 397296 273258 397352
rect 273253 397292 273300 397296
rect 273364 397294 273410 397354
rect 273621 397352 274404 397354
rect 273621 397296 273626 397352
rect 273682 397296 274404 397352
rect 273621 397294 274404 397296
rect 273364 397292 273370 397294
rect 273253 397291 273319 397292
rect 273621 397291 273687 397294
rect 274398 397292 274404 397294
rect 274468 397292 274474 397356
rect 274725 397354 274791 397357
rect 275318 397354 275324 397356
rect 274725 397352 275324 397354
rect 274725 397296 274730 397352
rect 274786 397296 275324 397352
rect 274725 397294 275324 397296
rect 274725 397291 274791 397294
rect 275318 397292 275324 397294
rect 275388 397292 275394 397356
rect 276381 397354 276447 397357
rect 278037 397356 278103 397357
rect 276974 397354 276980 397356
rect 276381 397352 276980 397354
rect 276381 397296 276386 397352
rect 276442 397296 276980 397352
rect 276381 397294 276980 397296
rect 276381 397291 276447 397294
rect 276974 397292 276980 397294
rect 277044 397292 277050 397356
rect 278037 397352 278084 397356
rect 278148 397354 278154 397356
rect 290181 397354 290247 397357
rect 293309 397356 293375 397357
rect 298461 397356 298527 397357
rect 308581 397356 308647 397357
rect 310973 397356 311039 397357
rect 313365 397356 313431 397357
rect 290958 397354 290964 397356
rect 278037 397296 278042 397352
rect 278037 397292 278084 397296
rect 278148 397294 278194 397354
rect 290181 397352 290964 397354
rect 290181 397296 290186 397352
rect 290242 397296 290964 397352
rect 290181 397294 290964 397296
rect 278148 397292 278154 397294
rect 278037 397291 278103 397292
rect 290181 397291 290247 397294
rect 290958 397292 290964 397294
rect 291028 397292 291034 397356
rect 293309 397352 293356 397356
rect 293420 397354 293426 397356
rect 293309 397296 293314 397352
rect 293309 397292 293356 397296
rect 293420 397294 293466 397354
rect 298461 397352 298508 397356
rect 298572 397354 298578 397356
rect 298461 397296 298466 397352
rect 293420 397292 293426 397294
rect 298461 397292 298508 397296
rect 298572 397294 298618 397354
rect 308581 397352 308628 397356
rect 308692 397354 308698 397356
rect 308581 397296 308586 397352
rect 298572 397292 298578 397294
rect 308581 397292 308628 397296
rect 308692 397294 308738 397354
rect 310973 397352 311020 397356
rect 311084 397354 311090 397356
rect 310973 397296 310978 397352
rect 308692 397292 308698 397294
rect 310973 397292 311020 397296
rect 311084 397294 311130 397354
rect 313365 397352 313412 397356
rect 313476 397354 313482 397356
rect 342253 397354 342319 397357
rect 343214 397354 343220 397356
rect 313365 397296 313370 397352
rect 311084 397292 311090 397294
rect 313365 397292 313412 397296
rect 313476 397294 313522 397354
rect 342253 397352 343220 397354
rect 342253 397296 342258 397352
rect 342314 397296 343220 397352
rect 342253 397294 343220 397296
rect 313476 397292 313482 397294
rect 293309 397291 293375 397292
rect 298461 397291 298527 397292
rect 308581 397291 308647 397292
rect 310973 397291 311039 397292
rect 313365 397291 313431 397292
rect 342253 397291 342319 397294
rect 343214 397292 343220 397294
rect 343284 397292 343290 397356
rect 96429 397220 96495 397221
rect 98453 397220 98519 397221
rect 96429 397216 96476 397220
rect 96540 397218 96546 397220
rect 96429 397160 96434 397216
rect 96429 397156 96476 397160
rect 96540 397158 96586 397218
rect 98453 397216 98500 397220
rect 98564 397218 98570 397220
rect 98453 397160 98458 397216
rect 96540 397156 96546 397158
rect 98453 397156 98500 397160
rect 98564 397158 98610 397218
rect 98564 397156 98570 397158
rect 103830 397156 103836 397220
rect 103900 397218 103906 397220
rect 104801 397218 104867 397221
rect 103900 397216 104867 397218
rect 103900 397160 104806 397216
rect 104862 397160 104867 397216
rect 103900 397158 104867 397160
rect 103900 397156 103906 397158
rect 96429 397155 96495 397156
rect 98453 397155 98519 397156
rect 104801 397155 104867 397158
rect 113173 397220 113239 397221
rect 263869 397220 263935 397221
rect 273437 397220 273503 397221
rect 113173 397216 113220 397220
rect 113284 397218 113290 397220
rect 113173 397160 113178 397216
rect 113173 397156 113220 397160
rect 113284 397158 113330 397218
rect 263869 397216 263916 397220
rect 263980 397218 263986 397220
rect 263869 397160 263874 397216
rect 113284 397156 113290 397158
rect 263869 397156 263916 397160
rect 263980 397158 264026 397218
rect 273437 397216 273484 397220
rect 273548 397218 273554 397220
rect 273437 397160 273442 397216
rect 263980 397156 263986 397158
rect 273437 397156 273484 397160
rect 273548 397158 273594 397218
rect 273548 397156 273554 397158
rect 113173 397155 113239 397156
rect 263869 397155 263935 397156
rect 273437 397155 273503 397156
rect 258073 396946 258139 396949
rect 258390 396946 258396 396948
rect 258073 396944 258396 396946
rect 258073 396888 258078 396944
rect 258134 396888 258396 396944
rect 258073 396886 258396 396888
rect 258073 396883 258139 396886
rect 258390 396884 258396 396886
rect 258460 396884 258466 396948
rect 76046 396748 76052 396812
rect 76116 396810 76122 396812
rect 77201 396810 77267 396813
rect 76116 396808 77267 396810
rect 76116 396752 77206 396808
rect 77262 396752 77267 396808
rect 76116 396750 77267 396752
rect 76116 396748 76122 396750
rect 77201 396747 77267 396750
rect 81934 396748 81940 396812
rect 82004 396810 82010 396812
rect 82721 396810 82787 396813
rect 82004 396808 82787 396810
rect 82004 396752 82726 396808
rect 82782 396752 82787 396808
rect 82004 396750 82787 396752
rect 82004 396748 82010 396750
rect 82721 396747 82787 396750
rect 84326 396748 84332 396812
rect 84396 396810 84402 396812
rect 85481 396810 85547 396813
rect 84396 396808 85547 396810
rect 84396 396752 85486 396808
rect 85542 396752 85547 396808
rect 84396 396750 85547 396752
rect 84396 396748 84402 396750
rect 85481 396747 85547 396750
rect 88374 396748 88380 396812
rect 88444 396810 88450 396812
rect 89621 396810 89687 396813
rect 88444 396808 89687 396810
rect 88444 396752 89626 396808
rect 89682 396752 89687 396808
rect 88444 396750 89687 396752
rect 88444 396748 88450 396750
rect 89621 396747 89687 396750
rect 90030 396748 90036 396812
rect 90100 396810 90106 396812
rect 91001 396810 91067 396813
rect 93761 396812 93827 396813
rect 93710 396810 93716 396812
rect 90100 396808 91067 396810
rect 90100 396752 91006 396808
rect 91062 396752 91067 396808
rect 90100 396750 91067 396752
rect 93670 396750 93716 396810
rect 93780 396808 93827 396812
rect 93822 396752 93827 396808
rect 90100 396748 90106 396750
rect 91001 396747 91067 396750
rect 93710 396748 93716 396750
rect 93780 396748 93827 396752
rect 94630 396748 94636 396812
rect 94700 396810 94706 396812
rect 95141 396810 95207 396813
rect 94700 396808 95207 396810
rect 94700 396752 95146 396808
rect 95202 396752 95207 396808
rect 94700 396750 95207 396752
rect 94700 396748 94706 396750
rect 93761 396747 93827 396748
rect 95141 396747 95207 396750
rect 97022 396748 97028 396812
rect 97092 396810 97098 396812
rect 97901 396810 97967 396813
rect 97092 396808 97967 396810
rect 97092 396752 97906 396808
rect 97962 396752 97967 396808
rect 97092 396750 97967 396752
rect 97092 396748 97098 396750
rect 97901 396747 97967 396750
rect 101070 396748 101076 396812
rect 101140 396810 101146 396812
rect 101949 396810 102015 396813
rect 101140 396808 102015 396810
rect 101140 396752 101954 396808
rect 102010 396752 102015 396808
rect 101140 396750 102015 396752
rect 101140 396748 101146 396750
rect 101949 396747 102015 396750
rect 105997 396812 106063 396813
rect 105997 396808 106044 396812
rect 106108 396810 106114 396812
rect 107377 396810 107443 396813
rect 108849 396812 108915 396813
rect 107510 396810 107516 396812
rect 105997 396752 106002 396808
rect 105997 396748 106044 396752
rect 106108 396750 106154 396810
rect 107377 396808 107516 396810
rect 107377 396752 107382 396808
rect 107438 396752 107516 396808
rect 107377 396750 107516 396752
rect 106108 396748 106114 396750
rect 105997 396747 106063 396748
rect 107377 396747 107443 396750
rect 107510 396748 107516 396750
rect 107580 396748 107586 396812
rect 108798 396810 108804 396812
rect 108758 396750 108804 396810
rect 108868 396808 108915 396812
rect 108910 396752 108915 396808
rect 108798 396748 108804 396750
rect 108868 396748 108915 396752
rect 111006 396748 111012 396812
rect 111076 396810 111082 396812
rect 111517 396810 111583 396813
rect 111076 396808 111583 396810
rect 111076 396752 111522 396808
rect 111578 396752 111583 396808
rect 111076 396750 111583 396752
rect 111076 396748 111082 396750
rect 108849 396747 108915 396748
rect 111517 396747 111583 396750
rect 112294 396748 112300 396812
rect 112364 396810 112370 396812
rect 113081 396810 113147 396813
rect 112364 396808 113147 396810
rect 112364 396752 113086 396808
rect 113142 396752 113147 396808
rect 112364 396750 113147 396752
rect 112364 396748 112370 396750
rect 113081 396747 113147 396750
rect 117078 396748 117084 396812
rect 117148 396810 117154 396812
rect 117221 396810 117287 396813
rect 117148 396808 117287 396810
rect 117148 396752 117226 396808
rect 117282 396752 117287 396808
rect 117148 396750 117287 396752
rect 117148 396748 117154 396750
rect 117221 396747 117287 396750
rect 118182 396748 118188 396812
rect 118252 396810 118258 396812
rect 118601 396810 118667 396813
rect 118252 396808 118667 396810
rect 118252 396752 118606 396808
rect 118662 396752 118667 396808
rect 118252 396750 118667 396752
rect 118252 396748 118258 396750
rect 118601 396747 118667 396750
rect 119102 396748 119108 396812
rect 119172 396810 119178 396812
rect 119889 396810 119955 396813
rect 119172 396808 119955 396810
rect 119172 396752 119894 396808
rect 119950 396752 119955 396808
rect 119172 396750 119955 396752
rect 119172 396748 119178 396750
rect 119889 396747 119955 396750
rect 120758 396748 120764 396812
rect 120828 396810 120834 396812
rect 121361 396810 121427 396813
rect 120828 396808 121427 396810
rect 120828 396752 121366 396808
rect 121422 396752 121427 396808
rect 120828 396750 121427 396752
rect 120828 396748 120834 396750
rect 121361 396747 121427 396750
rect 123518 396748 123524 396812
rect 123588 396810 123594 396812
rect 124121 396810 124187 396813
rect 123588 396808 124187 396810
rect 123588 396752 124126 396808
rect 124182 396752 124187 396808
rect 123588 396750 124187 396752
rect 123588 396748 123594 396750
rect 124121 396747 124187 396750
rect 125910 396748 125916 396812
rect 125980 396810 125986 396812
rect 126881 396810 126947 396813
rect 125980 396808 126947 396810
rect 125980 396752 126886 396808
rect 126942 396752 126947 396808
rect 125980 396750 126947 396752
rect 125980 396748 125986 396750
rect 126881 396747 126947 396750
rect 128670 396748 128676 396812
rect 128740 396810 128746 396812
rect 129641 396810 129707 396813
rect 128740 396808 129707 396810
rect 128740 396752 129646 396808
rect 129702 396752 129707 396808
rect 128740 396750 129707 396752
rect 128740 396748 128746 396750
rect 129641 396747 129707 396750
rect 131021 396812 131087 396813
rect 131021 396808 131068 396812
rect 131132 396810 131138 396812
rect 131021 396752 131026 396808
rect 131021 396748 131068 396752
rect 131132 396750 131178 396810
rect 131132 396748 131138 396750
rect 133454 396748 133460 396812
rect 133524 396810 133530 396812
rect 133781 396810 133847 396813
rect 133524 396808 133847 396810
rect 133524 396752 133786 396808
rect 133842 396752 133847 396808
rect 133524 396750 133847 396752
rect 133524 396748 133530 396750
rect 131021 396747 131087 396748
rect 133781 396747 133847 396750
rect 140773 396812 140839 396813
rect 140773 396808 140820 396812
rect 140884 396810 140890 396812
rect 140773 396752 140778 396808
rect 140773 396748 140820 396752
rect 140884 396750 140930 396810
rect 140884 396748 140890 396750
rect 143574 396748 143580 396812
rect 143644 396810 143650 396812
rect 144821 396810 144887 396813
rect 143644 396808 144887 396810
rect 143644 396752 144826 396808
rect 144882 396752 144887 396808
rect 143644 396750 144887 396752
rect 143644 396748 143650 396750
rect 140773 396747 140839 396748
rect 144821 396747 144887 396750
rect 145598 396748 145604 396812
rect 145668 396810 145674 396812
rect 146201 396810 146267 396813
rect 145668 396808 146267 396810
rect 145668 396752 146206 396808
rect 146262 396752 146267 396808
rect 145668 396750 146267 396752
rect 145668 396748 145674 396750
rect 146201 396747 146267 396750
rect 147673 396810 147739 396813
rect 148542 396810 148548 396812
rect 147673 396808 148548 396810
rect 147673 396752 147678 396808
rect 147734 396752 148548 396808
rect 147673 396750 148548 396752
rect 147673 396747 147739 396750
rect 148542 396748 148548 396750
rect 148612 396748 148618 396812
rect 154062 396748 154068 396812
rect 154132 396810 154138 396812
rect 154481 396810 154547 396813
rect 155953 396812 156019 396813
rect 155902 396810 155908 396812
rect 154132 396808 154547 396810
rect 154132 396752 154486 396808
rect 154542 396752 154547 396808
rect 154132 396750 154547 396752
rect 155862 396750 155908 396810
rect 155972 396808 156019 396812
rect 156014 396752 156019 396808
rect 154132 396748 154138 396750
rect 154481 396747 154547 396750
rect 155902 396748 155908 396750
rect 155972 396748 156019 396752
rect 158478 396748 158484 396812
rect 158548 396810 158554 396812
rect 158621 396810 158687 396813
rect 158548 396808 158687 396810
rect 158548 396752 158626 396808
rect 158682 396752 158687 396808
rect 158548 396750 158687 396752
rect 158548 396748 158554 396750
rect 155953 396747 156019 396748
rect 158621 396747 158687 396750
rect 160870 396748 160876 396812
rect 160940 396810 160946 396812
rect 161381 396810 161447 396813
rect 160940 396808 161447 396810
rect 160940 396752 161386 396808
rect 161442 396752 161447 396808
rect 160940 396750 161447 396752
rect 160940 396748 160946 396750
rect 161381 396747 161447 396750
rect 163446 396748 163452 396812
rect 163516 396810 163522 396812
rect 164141 396810 164207 396813
rect 163516 396808 164207 396810
rect 163516 396752 164146 396808
rect 164202 396752 164207 396808
rect 163516 396750 164207 396752
rect 163516 396748 163522 396750
rect 164141 396747 164207 396750
rect 166022 396748 166028 396812
rect 166092 396810 166098 396812
rect 166901 396810 166967 396813
rect 183185 396812 183251 396813
rect 183134 396810 183140 396812
rect 166092 396808 166967 396810
rect 166092 396752 166906 396808
rect 166962 396752 166967 396808
rect 166092 396750 166967 396752
rect 183094 396750 183140 396810
rect 183204 396808 183251 396812
rect 183246 396752 183251 396808
rect 166092 396748 166098 396750
rect 166901 396747 166967 396750
rect 183134 396748 183140 396750
rect 183204 396748 183251 396752
rect 183185 396747 183251 396748
rect 237373 396810 237439 396813
rect 238150 396810 238156 396812
rect 237373 396808 238156 396810
rect 237373 396752 237378 396808
rect 237434 396752 238156 396808
rect 237373 396750 238156 396752
rect 237373 396747 237439 396750
rect 238150 396748 238156 396750
rect 238220 396748 238226 396812
rect 240133 396810 240199 396813
rect 240542 396810 240548 396812
rect 240133 396808 240548 396810
rect 240133 396752 240138 396808
rect 240194 396752 240548 396808
rect 240133 396750 240548 396752
rect 240133 396747 240199 396750
rect 240542 396748 240548 396750
rect 240612 396748 240618 396812
rect 244222 396748 244228 396812
rect 244292 396810 244298 396812
rect 244365 396810 244431 396813
rect 244292 396808 244431 396810
rect 244292 396752 244370 396808
rect 244426 396752 244431 396808
rect 244292 396750 244431 396752
rect 244292 396748 244298 396750
rect 244365 396747 244431 396750
rect 245653 396810 245719 396813
rect 246430 396810 246436 396812
rect 245653 396808 246436 396810
rect 245653 396752 245658 396808
rect 245714 396752 246436 396808
rect 245653 396750 246436 396752
rect 245653 396747 245719 396750
rect 246430 396748 246436 396750
rect 246500 396748 246506 396812
rect 247125 396810 247191 396813
rect 248270 396810 248276 396812
rect 247125 396808 248276 396810
rect 247125 396752 247130 396808
rect 247186 396752 248276 396808
rect 247125 396750 248276 396752
rect 247125 396747 247191 396750
rect 248270 396748 248276 396750
rect 248340 396748 248346 396812
rect 249885 396810 249951 396813
rect 251265 396812 251331 396813
rect 250110 396810 250116 396812
rect 249885 396808 250116 396810
rect 249885 396752 249890 396808
rect 249946 396752 250116 396808
rect 249885 396750 250116 396752
rect 249885 396747 249951 396750
rect 250110 396748 250116 396750
rect 250180 396748 250186 396812
rect 251214 396810 251220 396812
rect 251174 396750 251220 396810
rect 251284 396808 251331 396812
rect 251326 396752 251331 396808
rect 251214 396748 251220 396750
rect 251284 396748 251331 396752
rect 251265 396747 251331 396748
rect 254485 396812 254551 396813
rect 254485 396808 254532 396812
rect 254596 396810 254602 396812
rect 255313 396810 255379 396813
rect 255814 396810 255820 396812
rect 254485 396752 254490 396808
rect 254485 396748 254532 396752
rect 254596 396750 254642 396810
rect 255313 396808 255820 396810
rect 255313 396752 255318 396808
rect 255374 396752 255820 396808
rect 255313 396750 255820 396752
rect 254596 396748 254602 396750
rect 254485 396747 254551 396748
rect 255313 396747 255379 396750
rect 255814 396748 255820 396750
rect 255884 396748 255890 396812
rect 256693 396810 256759 396813
rect 256918 396810 256924 396812
rect 256693 396808 256924 396810
rect 256693 396752 256698 396808
rect 256754 396752 256924 396808
rect 256693 396750 256924 396752
rect 256693 396747 256759 396750
rect 256918 396748 256924 396750
rect 256988 396748 256994 396812
rect 258165 396810 258231 396813
rect 259453 396812 259519 396813
rect 258390 396810 258396 396812
rect 258165 396808 258396 396810
rect 258165 396752 258170 396808
rect 258226 396752 258396 396808
rect 258165 396750 258396 396752
rect 258165 396747 258231 396750
rect 258390 396748 258396 396750
rect 258460 396748 258466 396812
rect 259453 396808 259500 396812
rect 259564 396810 259570 396812
rect 262213 396810 262279 396813
rect 262806 396810 262812 396812
rect 259453 396752 259458 396808
rect 259453 396748 259500 396752
rect 259564 396750 259610 396810
rect 262213 396808 262812 396810
rect 262213 396752 262218 396808
rect 262274 396752 262812 396808
rect 262213 396750 262812 396752
rect 259564 396748 259570 396750
rect 259453 396747 259519 396748
rect 262213 396747 262279 396750
rect 262806 396748 262812 396750
rect 262876 396748 262882 396812
rect 265249 396810 265315 396813
rect 265934 396810 265940 396812
rect 265249 396808 265940 396810
rect 265249 396752 265254 396808
rect 265310 396752 265940 396808
rect 265249 396750 265940 396752
rect 265249 396747 265315 396750
rect 265934 396748 265940 396750
rect 266004 396748 266010 396812
rect 266302 396748 266308 396812
rect 266372 396810 266378 396812
rect 266445 396810 266511 396813
rect 266372 396808 266511 396810
rect 266372 396752 266450 396808
rect 266506 396752 266511 396808
rect 266372 396750 266511 396752
rect 266372 396748 266378 396750
rect 266445 396747 266511 396750
rect 267825 396810 267891 396813
rect 268326 396810 268332 396812
rect 267825 396808 268332 396810
rect 267825 396752 267830 396808
rect 267886 396752 268332 396808
rect 267825 396750 268332 396752
rect 267825 396747 267891 396750
rect 268326 396748 268332 396750
rect 268396 396748 268402 396812
rect 269113 396810 269179 396813
rect 269798 396810 269804 396812
rect 269113 396808 269804 396810
rect 269113 396752 269118 396808
rect 269174 396752 269804 396808
rect 269113 396750 269804 396752
rect 269113 396747 269179 396750
rect 269798 396748 269804 396750
rect 269868 396748 269874 396812
rect 270585 396810 270651 396813
rect 272517 396812 272583 396813
rect 270902 396810 270908 396812
rect 270585 396808 270908 396810
rect 270585 396752 270590 396808
rect 270646 396752 270908 396808
rect 270585 396750 270908 396752
rect 270585 396747 270651 396750
rect 270902 396748 270908 396750
rect 270972 396748 270978 396812
rect 272517 396808 272564 396812
rect 272628 396810 272634 396812
rect 276105 396810 276171 396813
rect 276238 396810 276244 396812
rect 272517 396752 272522 396808
rect 272517 396748 272564 396752
rect 272628 396750 272674 396810
rect 276105 396808 276244 396810
rect 276105 396752 276110 396808
rect 276166 396752 276244 396808
rect 276105 396750 276244 396752
rect 272628 396748 272634 396750
rect 272517 396747 272583 396748
rect 276105 396747 276171 396750
rect 276238 396748 276244 396750
rect 276308 396748 276314 396812
rect 277485 396810 277551 396813
rect 278446 396810 278452 396812
rect 277485 396808 278452 396810
rect 277485 396752 277490 396808
rect 277546 396752 278452 396808
rect 277485 396750 278452 396752
rect 277485 396747 277551 396750
rect 278446 396748 278452 396750
rect 278516 396748 278522 396812
rect 278773 396810 278839 396813
rect 278998 396810 279004 396812
rect 278773 396808 279004 396810
rect 278773 396752 278778 396808
rect 278834 396752 279004 396808
rect 278773 396750 279004 396752
rect 278773 396747 278839 396750
rect 278998 396748 279004 396750
rect 279068 396748 279074 396812
rect 280153 396810 280219 396813
rect 280838 396810 280844 396812
rect 280153 396808 280844 396810
rect 280153 396752 280158 396808
rect 280214 396752 280844 396808
rect 280153 396750 280844 396752
rect 280153 396747 280219 396750
rect 280838 396748 280844 396750
rect 280908 396748 280914 396812
rect 283557 396810 283623 396813
rect 285949 396812 286015 396813
rect 283782 396810 283788 396812
rect 283557 396808 283788 396810
rect 283557 396752 283562 396808
rect 283618 396752 283788 396808
rect 283557 396750 283788 396752
rect 283557 396747 283623 396750
rect 283782 396748 283788 396750
rect 283852 396748 283858 396812
rect 285949 396808 285996 396812
rect 286060 396810 286066 396812
rect 287053 396810 287119 396813
rect 288198 396810 288204 396812
rect 285949 396752 285954 396808
rect 285949 396748 285996 396752
rect 286060 396750 286106 396810
rect 287053 396808 288204 396810
rect 287053 396752 287058 396808
rect 287114 396752 288204 396808
rect 287053 396750 288204 396752
rect 286060 396748 286066 396750
rect 285949 396747 286015 396748
rect 287053 396747 287119 396750
rect 288198 396748 288204 396750
rect 288268 396748 288274 396812
rect 295333 396810 295399 396813
rect 295926 396810 295932 396812
rect 295333 396808 295932 396810
rect 295333 396752 295338 396808
rect 295394 396752 295932 396808
rect 295333 396750 295932 396752
rect 295333 396747 295399 396750
rect 295926 396748 295932 396750
rect 295996 396748 296002 396812
rect 302233 396810 302299 396813
rect 303470 396810 303476 396812
rect 302233 396808 303476 396810
rect 302233 396752 302238 396808
rect 302294 396752 303476 396808
rect 302233 396750 303476 396752
rect 302233 396747 302299 396750
rect 303470 396748 303476 396750
rect 303540 396748 303546 396812
rect 304993 396810 305059 396813
rect 305862 396810 305868 396812
rect 304993 396808 305868 396810
rect 304993 396752 304998 396808
rect 305054 396752 305868 396808
rect 304993 396750 305868 396752
rect 304993 396747 305059 396750
rect 305862 396748 305868 396750
rect 305932 396748 305938 396812
rect 317413 396810 317479 396813
rect 318374 396810 318380 396812
rect 317413 396808 318380 396810
rect 317413 396752 317418 396808
rect 317474 396752 318380 396808
rect 317413 396750 318380 396752
rect 317413 396747 317479 396750
rect 318374 396748 318380 396750
rect 318444 396748 318450 396812
rect 320173 396810 320239 396813
rect 320950 396810 320956 396812
rect 320173 396808 320956 396810
rect 320173 396752 320178 396808
rect 320234 396752 320956 396808
rect 320173 396750 320956 396752
rect 320173 396747 320239 396750
rect 320950 396748 320956 396750
rect 321020 396748 321026 396812
rect 322933 396810 322999 396813
rect 323342 396810 323348 396812
rect 322933 396808 323348 396810
rect 322933 396752 322938 396808
rect 322994 396752 323348 396808
rect 322933 396750 323348 396752
rect 322933 396747 322999 396750
rect 323342 396748 323348 396750
rect 323412 396748 323418 396812
rect 342345 396810 342411 396813
rect 343398 396810 343404 396812
rect 342345 396808 343404 396810
rect 342345 396752 342350 396808
rect 342406 396752 343404 396808
rect 342345 396750 343404 396752
rect 342345 396747 342411 396750
rect 343398 396748 343404 396750
rect 343468 396748 343474 396812
rect 75913 396674 75979 396677
rect 77150 396674 77156 396676
rect 75913 396672 77156 396674
rect 75913 396616 75918 396672
rect 75974 396616 77156 396672
rect 75913 396614 77156 396616
rect 75913 396611 75979 396614
rect 77150 396612 77156 396614
rect 77220 396612 77226 396676
rect 89713 396674 89779 396677
rect 90766 396674 90772 396676
rect 89713 396672 90772 396674
rect 89713 396616 89718 396672
rect 89774 396616 90772 396672
rect 89713 396614 90772 396616
rect 89713 396611 89779 396614
rect 90766 396612 90772 396614
rect 90836 396612 90842 396676
rect 91093 396674 91159 396677
rect 91502 396674 91508 396676
rect 91093 396672 91508 396674
rect 91093 396616 91098 396672
rect 91154 396616 91508 396672
rect 91093 396614 91508 396616
rect 91093 396611 91159 396614
rect 91502 396612 91508 396614
rect 91572 396612 91578 396676
rect 108246 396612 108252 396676
rect 108316 396674 108322 396676
rect 108941 396674 109007 396677
rect 108316 396672 109007 396674
rect 108316 396616 108946 396672
rect 109002 396616 109007 396672
rect 108316 396614 109007 396616
rect 108316 396612 108322 396614
rect 108941 396611 109007 396614
rect 115974 396612 115980 396676
rect 116044 396674 116050 396676
rect 117129 396674 117195 396677
rect 116044 396672 117195 396674
rect 116044 396616 117134 396672
rect 117190 396616 117195 396672
rect 116044 396614 117195 396616
rect 116044 396612 116050 396614
rect 117129 396611 117195 396614
rect 247677 396676 247743 396677
rect 247677 396672 247724 396676
rect 247788 396674 247794 396676
rect 251173 396674 251239 396677
rect 252318 396674 252324 396676
rect 247677 396616 247682 396672
rect 247677 396612 247724 396616
rect 247788 396614 247834 396674
rect 251173 396672 252324 396674
rect 251173 396616 251178 396672
rect 251234 396616 252324 396672
rect 251173 396614 252324 396616
rect 247788 396612 247794 396614
rect 247677 396611 247743 396612
rect 251173 396611 251239 396614
rect 252318 396612 252324 396614
rect 252388 396612 252394 396676
rect 259545 396674 259611 396677
rect 260598 396674 260604 396676
rect 259545 396672 260604 396674
rect 259545 396616 259550 396672
rect 259606 396616 260604 396672
rect 259545 396614 260604 396616
rect 259545 396611 259611 396614
rect 260598 396612 260604 396614
rect 260668 396612 260674 396676
rect 266353 396674 266419 396677
rect 267590 396674 267596 396676
rect 266353 396672 267596 396674
rect 266353 396616 266358 396672
rect 266414 396616 267596 396672
rect 266353 396614 267596 396616
rect 266353 396611 266419 396614
rect 267590 396612 267596 396614
rect 267660 396612 267666 396676
rect 267733 396674 267799 396677
rect 268694 396674 268700 396676
rect 267733 396672 268700 396674
rect 267733 396616 267738 396672
rect 267794 396616 268700 396672
rect 267733 396614 268700 396616
rect 267733 396611 267799 396614
rect 268694 396612 268700 396614
rect 268764 396612 268770 396676
rect 218605 393410 218671 393413
rect 219382 393410 219388 393412
rect 218605 393408 219388 393410
rect 218605 393352 218610 393408
rect 218666 393352 219388 393408
rect 218605 393350 219388 393352
rect 218605 393347 218671 393350
rect 219382 393348 219388 393350
rect 219452 393348 219458 393412
rect 219198 392804 219204 392868
rect 219268 392866 219274 392868
rect 219341 392866 219407 392869
rect 219268 392864 219407 392866
rect 219268 392808 219346 392864
rect 219402 392808 219407 392864
rect 219268 392806 219407 392808
rect 219268 392804 219274 392806
rect 219341 392803 219407 392806
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 219341 383890 219407 383893
rect 219206 383888 219407 383890
rect 219206 383832 219346 383888
rect 219402 383832 219407 383888
rect 219206 383830 219407 383832
rect 219206 383756 219266 383830
rect 219341 383827 219407 383830
rect 219198 383692 219204 383756
rect 219268 383692 219274 383756
rect 219065 383618 219131 383621
rect 219382 383618 219388 383620
rect 219065 383616 219388 383618
rect 219065 383560 219070 383616
rect 219126 383560 219388 383616
rect 219065 383558 219388 383560
rect 219065 383555 219131 383558
rect 219382 383556 219388 383558
rect 219452 383556 219458 383620
rect 580165 378450 580231 378453
rect 583520 378450 584960 378540
rect 580165 378448 584960 378450
rect 580165 378392 580170 378448
rect 580226 378392 584960 378448
rect 580165 378390 584960 378392
rect 580165 378387 580231 378390
rect 583520 378300 584960 378390
rect 219065 374234 219131 374237
rect 219382 374234 219388 374236
rect 219065 374232 219388 374234
rect 219065 374176 219070 374232
rect 219126 374176 219388 374232
rect 219065 374174 219388 374176
rect 219065 374171 219131 374174
rect 219382 374172 219388 374174
rect 219452 374172 219458 374236
rect 218973 373962 219039 373965
rect 219382 373962 219388 373964
rect 218973 373960 219388 373962
rect 218973 373904 218978 373960
rect 219034 373904 219388 373960
rect 218973 373902 219388 373904
rect 218973 373899 219039 373902
rect 219382 373900 219388 373902
rect 219452 373900 219458 373964
rect -960 371378 480 371468
rect 3417 371378 3483 371381
rect -960 371376 3483 371378
rect -960 371320 3422 371376
rect 3478 371320 3483 371376
rect -960 371318 3483 371320
rect -960 371228 480 371318
rect 3417 371315 3483 371318
rect 579613 365122 579679 365125
rect 583520 365122 584960 365212
rect 579613 365120 584960 365122
rect 579613 365064 579618 365120
rect 579674 365064 584960 365120
rect 579613 365062 584960 365064
rect 579613 365059 579679 365062
rect 583520 364972 584960 365062
rect 218973 364442 219039 364445
rect 219382 364442 219388 364444
rect 218973 364440 219388 364442
rect 218973 364384 218978 364440
rect 219034 364384 219388 364440
rect 218973 364382 219388 364384
rect 218973 364379 219039 364382
rect 219382 364380 219388 364382
rect 219452 364380 219458 364444
rect 218973 364306 219039 364309
rect 219382 364306 219388 364308
rect 218973 364304 219388 364306
rect 218973 364248 218978 364304
rect 219034 364248 219388 364304
rect 218973 364246 219388 364248
rect 218973 364243 219039 364246
rect 219382 364244 219388 364246
rect 219452 364244 219458 364308
rect -960 358458 480 358548
rect 3141 358458 3207 358461
rect -960 358456 3207 358458
rect -960 358400 3146 358456
rect 3202 358400 3207 358456
rect -960 358398 3207 358400
rect -960 358308 480 358398
rect 3141 358395 3207 358398
rect 218973 354786 219039 354789
rect 219382 354786 219388 354788
rect 218973 354784 219388 354786
rect 218973 354728 218978 354784
rect 219034 354728 219388 354784
rect 218973 354726 219388 354728
rect 218973 354723 219039 354726
rect 219382 354724 219388 354726
rect 219452 354724 219458 354788
rect 218973 354650 219039 354653
rect 219382 354650 219388 354652
rect 218973 354648 219388 354650
rect 218973 354592 218978 354648
rect 219034 354592 219388 354648
rect 218973 354590 219388 354592
rect 218973 354587 219039 354590
rect 219382 354588 219388 354590
rect 219452 354588 219458 354652
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 3325 345402 3391 345405
rect -960 345400 3391 345402
rect -960 345344 3330 345400
rect 3386 345344 3391 345400
rect -960 345342 3391 345344
rect -960 345252 480 345342
rect 3325 345339 3391 345342
rect 218973 345130 219039 345133
rect 219382 345130 219388 345132
rect 218973 345128 219388 345130
rect 218973 345072 218978 345128
rect 219034 345072 219388 345128
rect 218973 345070 219388 345072
rect 218973 345067 219039 345070
rect 219382 345068 219388 345070
rect 219452 345068 219458 345132
rect 219065 344586 219131 344589
rect 219198 344586 219204 344588
rect 219065 344584 219204 344586
rect 219065 344528 219070 344584
rect 219126 344528 219204 344584
rect 219065 344526 219204 344528
rect 219065 344523 219131 344526
rect 219198 344524 219204 344526
rect 219268 344524 219274 344588
rect 583520 338452 584960 338692
rect 219065 335474 219131 335477
rect 219198 335474 219204 335476
rect 219065 335472 219204 335474
rect 219065 335416 219070 335472
rect 219126 335416 219204 335472
rect 219065 335414 219204 335416
rect 219065 335411 219131 335414
rect 219198 335412 219204 335414
rect 219268 335412 219274 335476
rect 219198 335004 219204 335068
rect 219268 335066 219274 335068
rect 219341 335066 219407 335069
rect 219268 335064 219407 335066
rect 219268 335008 219346 335064
rect 219402 335008 219407 335064
rect 219268 335006 219407 335008
rect 219268 335004 219274 335006
rect 219341 335003 219407 335006
rect -960 332196 480 332436
rect 219198 325892 219204 325956
rect 219268 325954 219274 325956
rect 219341 325954 219407 325957
rect 219268 325952 219407 325954
rect 219268 325896 219346 325952
rect 219402 325896 219407 325952
rect 219268 325894 219407 325896
rect 219268 325892 219274 325894
rect 219341 325891 219407 325894
rect 219065 325682 219131 325685
rect 219382 325682 219388 325684
rect 219065 325680 219388 325682
rect 219065 325624 219070 325680
rect 219126 325624 219388 325680
rect 219065 325622 219388 325624
rect 219065 325619 219131 325622
rect 219382 325620 219388 325622
rect 219452 325620 219458 325684
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 3417 319290 3483 319293
rect -960 319288 3483 319290
rect -960 319232 3422 319288
rect 3478 319232 3483 319288
rect -960 319230 3483 319232
rect -960 319140 480 319230
rect 3417 319227 3483 319230
rect 219065 316298 219131 316301
rect 219382 316298 219388 316300
rect 219065 316296 219388 316298
rect 219065 316240 219070 316296
rect 219126 316240 219388 316296
rect 219065 316238 219388 316240
rect 219065 316235 219131 316238
rect 219382 316236 219388 316238
rect 219452 316236 219458 316300
rect 218973 316026 219039 316029
rect 219382 316026 219388 316028
rect 218973 316024 219388 316026
rect 218973 315968 218978 316024
rect 219034 315968 219388 316024
rect 218973 315966 219388 315968
rect 218973 315963 219039 315966
rect 219382 315964 219388 315966
rect 219452 315964 219458 316028
rect 579981 312082 580047 312085
rect 583520 312082 584960 312172
rect 579981 312080 584960 312082
rect 579981 312024 579986 312080
rect 580042 312024 584960 312080
rect 579981 312022 584960 312024
rect 579981 312019 580047 312022
rect 583520 311932 584960 312022
rect 218973 306506 219039 306509
rect 219382 306506 219388 306508
rect 218973 306504 219388 306506
rect 218973 306448 218978 306504
rect 219034 306448 219388 306504
rect 218973 306446 219388 306448
rect 218973 306443 219039 306446
rect 219382 306444 219388 306446
rect 219452 306444 219458 306508
rect 218973 306370 219039 306373
rect 219382 306370 219388 306372
rect 218973 306368 219388 306370
rect -960 306234 480 306324
rect 218973 306312 218978 306368
rect 219034 306312 219388 306368
rect 218973 306310 219388 306312
rect 218973 306307 219039 306310
rect 219382 306308 219388 306310
rect 219452 306308 219458 306372
rect 3233 306234 3299 306237
rect -960 306232 3299 306234
rect -960 306176 3238 306232
rect 3294 306176 3299 306232
rect -960 306174 3299 306176
rect -960 306084 480 306174
rect 3233 306171 3299 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect 218973 296850 219039 296853
rect 219382 296850 219388 296852
rect 218973 296848 219388 296850
rect 218973 296792 218978 296848
rect 219034 296792 219388 296848
rect 218973 296790 219388 296792
rect 218973 296787 219039 296790
rect 219382 296788 219388 296790
rect 219452 296788 219458 296852
rect 218973 296714 219039 296717
rect 219382 296714 219388 296716
rect 218973 296712 219388 296714
rect 218973 296656 218978 296712
rect 219034 296656 219388 296712
rect 218973 296654 219388 296656
rect 218973 296651 219039 296654
rect 219382 296652 219388 296654
rect 219452 296652 219458 296716
rect -960 293178 480 293268
rect 3417 293178 3483 293181
rect -960 293176 3483 293178
rect -960 293120 3422 293176
rect 3478 293120 3483 293176
rect -960 293118 3483 293120
rect -960 293028 480 293118
rect 3417 293115 3483 293118
rect 218973 287194 219039 287197
rect 219382 287194 219388 287196
rect 218973 287192 219388 287194
rect 218973 287136 218978 287192
rect 219034 287136 219388 287192
rect 218973 287134 219388 287136
rect 218973 287131 219039 287134
rect 219382 287132 219388 287134
rect 219452 287132 219458 287196
rect 218973 287058 219039 287061
rect 219382 287058 219388 287060
rect 218973 287056 219388 287058
rect 218973 287000 218978 287056
rect 219034 287000 219388 287056
rect 218973 286998 219388 287000
rect 218973 286995 219039 286998
rect 219382 286996 219388 286998
rect 219452 286996 219458 287060
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 218973 277538 219039 277541
rect 219382 277538 219388 277540
rect 218973 277536 219388 277538
rect 218973 277480 218978 277536
rect 219034 277480 219388 277536
rect 218973 277478 219388 277480
rect 218973 277475 219039 277478
rect 219382 277476 219388 277478
rect 219452 277476 219458 277540
rect 218973 277402 219039 277405
rect 219382 277402 219388 277404
rect 218973 277400 219388 277402
rect 218973 277344 218978 277400
rect 219034 277344 219388 277400
rect 218973 277342 219388 277344
rect 218973 277339 219039 277342
rect 219382 277340 219388 277342
rect 219452 277340 219458 277404
rect 580165 272234 580231 272237
rect 583520 272234 584960 272324
rect 580165 272232 584960 272234
rect 580165 272176 580170 272232
rect 580226 272176 584960 272232
rect 580165 272174 584960 272176
rect 580165 272171 580231 272174
rect 583520 272084 584960 272174
rect 218973 267882 219039 267885
rect 219382 267882 219388 267884
rect 218973 267880 219388 267882
rect 218973 267824 218978 267880
rect 219034 267824 219388 267880
rect 218973 267822 219388 267824
rect 218973 267819 219039 267822
rect 219382 267820 219388 267822
rect 219452 267820 219458 267884
rect 218421 267746 218487 267749
rect 219382 267746 219388 267748
rect 218421 267744 219388 267746
rect 218421 267688 218426 267744
rect 218482 267688 219388 267744
rect 218421 267686 219388 267688
rect 218421 267683 218487 267686
rect 219382 267684 219388 267686
rect 219452 267684 219458 267748
rect -960 267202 480 267292
rect 3049 267202 3115 267205
rect -960 267200 3115 267202
rect -960 267144 3054 267200
rect 3110 267144 3115 267200
rect -960 267142 3115 267144
rect -960 267052 480 267142
rect 3049 267139 3115 267142
rect 583520 258906 584960 258996
rect 583342 258846 584960 258906
rect 583342 258770 583402 258846
rect 583520 258770 584960 258846
rect 583342 258756 584960 258770
rect 583342 258710 583586 258756
rect 218421 258362 218487 258365
rect 219382 258362 219388 258364
rect 218421 258360 219388 258362
rect 218421 258304 218426 258360
rect 218482 258304 219388 258360
rect 218421 258302 219388 258304
rect 218421 258299 218487 258302
rect 219382 258300 219388 258302
rect 219452 258300 219458 258364
rect 218286 258166 219634 258226
rect 86217 257954 86283 257957
rect 218286 257954 218346 258166
rect 86217 257952 218346 257954
rect 86217 257896 86222 257952
rect 86278 257896 218346 257952
rect 86217 257894 218346 257896
rect 218421 257954 218487 257957
rect 219382 257954 219388 257956
rect 218421 257952 219388 257954
rect 218421 257896 218426 257952
rect 218482 257896 219388 257952
rect 218421 257894 219388 257896
rect 86217 257891 86283 257894
rect 218421 257891 218487 257894
rect 219382 257892 219388 257894
rect 219452 257892 219458 257956
rect 219574 257954 219634 258166
rect 583526 257954 583586 258710
rect 219574 257894 583586 257954
rect 141417 255914 141483 255917
rect 146937 255914 147003 255917
rect 141417 255912 147003 255914
rect 141417 255856 141422 255912
rect 141478 255856 146942 255912
rect 146998 255856 147003 255912
rect 141417 255854 147003 255856
rect 141417 255851 141483 255854
rect 146937 255851 147003 255854
rect -960 254146 480 254236
rect 3417 254146 3483 254149
rect -960 254144 3483 254146
rect -960 254088 3422 254144
rect 3478 254088 3483 254144
rect -960 254086 3483 254088
rect -960 253996 480 254086
rect 3417 254083 3483 254086
rect 124121 250474 124187 250477
rect 226241 250474 226307 250477
rect 124121 250472 226307 250474
rect 124121 250416 124126 250472
rect 124182 250416 226246 250472
rect 226302 250416 226307 250472
rect 124121 250414 226307 250416
rect 124121 250411 124187 250414
rect 226241 250411 226307 250414
rect 118601 249250 118667 249253
rect 230933 249250 230999 249253
rect 118601 249248 230999 249250
rect 118601 249192 118606 249248
rect 118662 249192 230938 249248
rect 230994 249192 230999 249248
rect 118601 249190 230999 249192
rect 118601 249187 118667 249190
rect 230933 249187 230999 249190
rect 3417 249114 3483 249117
rect 155953 249114 156019 249117
rect 3417 249112 156019 249114
rect 3417 249056 3422 249112
rect 3478 249056 155958 249112
rect 156014 249056 156019 249112
rect 3417 249054 156019 249056
rect 3417 249051 3483 249054
rect 155953 249051 156019 249054
rect 218421 248434 218487 248437
rect 219382 248434 219388 248436
rect 218421 248432 219388 248434
rect 218421 248376 218426 248432
rect 218482 248376 219388 248432
rect 218421 248374 219388 248376
rect 218421 248371 218487 248374
rect 219382 248372 219388 248374
rect 219452 248372 219458 248436
rect 218421 248026 218487 248029
rect 219198 248026 219204 248028
rect 218421 248024 219204 248026
rect 218421 247968 218426 248024
rect 218482 247968 219204 248024
rect 218421 247966 219204 247968
rect 218421 247963 218487 247966
rect 219198 247964 219204 247966
rect 219268 247964 219274 248028
rect 78581 247074 78647 247077
rect 281993 247074 282059 247077
rect 78581 247072 282059 247074
rect 78581 247016 78586 247072
rect 78642 247016 281998 247072
rect 282054 247016 282059 247072
rect 78581 247014 282059 247016
rect 78581 247011 78647 247014
rect 281993 247011 282059 247014
rect 138197 245714 138263 245717
rect 141417 245714 141483 245717
rect 138197 245712 141483 245714
rect 138197 245656 138202 245712
rect 138258 245656 141422 245712
rect 141478 245656 141483 245712
rect 138197 245654 141483 245656
rect 138197 245651 138263 245654
rect 141417 245651 141483 245654
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect 108941 244898 109007 244901
rect 225321 244898 225387 244901
rect 108941 244896 225387 244898
rect 108941 244840 108946 244896
rect 109002 244840 225326 244896
rect 225382 244840 225387 244896
rect 108941 244838 225387 244840
rect 108941 244835 109007 244838
rect 225321 244835 225387 244838
rect 113081 243538 113147 243541
rect 229553 243538 229619 243541
rect 113081 243536 229619 243538
rect 113081 243480 113086 243536
rect 113142 243480 229558 243536
rect 229614 243480 229619 243536
rect 113081 243478 229619 243480
rect 113081 243475 113147 243478
rect 229553 243475 229619 243478
rect 117221 242314 117287 242317
rect 229001 242314 229067 242317
rect 117221 242312 229067 242314
rect 117221 242256 117226 242312
rect 117282 242256 229006 242312
rect 229062 242256 229067 242312
rect 117221 242254 229067 242256
rect 117221 242251 117287 242254
rect 229001 242251 229067 242254
rect 58341 242178 58407 242181
rect 198825 242178 198891 242181
rect 58341 242176 198891 242178
rect 58341 242120 58346 242176
rect 58402 242120 198830 242176
rect 198886 242120 198891 242176
rect 58341 242118 198891 242120
rect 58341 242115 58407 242118
rect 198825 242115 198891 242118
rect -960 241090 480 241180
rect 4061 241090 4127 241093
rect -960 241088 4127 241090
rect -960 241032 4066 241088
rect 4122 241032 4127 241088
rect -960 241030 4127 241032
rect -960 240940 480 241030
rect 4061 241027 4127 241030
rect 124121 240818 124187 240821
rect 138197 240818 138263 240821
rect 124121 240816 138263 240818
rect 124121 240760 124126 240816
rect 124182 240760 138202 240816
rect 138258 240760 138263 240816
rect 124121 240758 138263 240760
rect 124121 240755 124187 240758
rect 138197 240755 138263 240758
rect 158621 240818 158687 240821
rect 225413 240818 225479 240821
rect 158621 240816 225479 240818
rect 158621 240760 158626 240816
rect 158682 240760 225418 240816
rect 225474 240760 225479 240816
rect 158621 240758 225479 240760
rect 158621 240755 158687 240758
rect 225413 240755 225479 240758
rect 57329 239458 57395 239461
rect 197353 239458 197419 239461
rect 57329 239456 197419 239458
rect 57329 239400 57334 239456
rect 57390 239400 197358 239456
rect 197414 239400 197419 239456
rect 57329 239398 197419 239400
rect 57329 239395 57395 239398
rect 197353 239395 197419 239398
rect 197905 239458 197971 239461
rect 226977 239458 227043 239461
rect 197905 239456 227043 239458
rect 197905 239400 197910 239456
rect 197966 239400 226982 239456
rect 227038 239400 227043 239456
rect 197905 239398 227043 239400
rect 197905 239395 197971 239398
rect 226977 239395 227043 239398
rect 218421 238914 218487 238917
rect 219382 238914 219388 238916
rect 218421 238912 219388 238914
rect 218421 238856 218426 238912
rect 218482 238856 219388 238912
rect 218421 238854 219388 238856
rect 218421 238851 218487 238854
rect 219382 238852 219388 238854
rect 219452 238852 219458 238916
rect 218513 238506 218579 238509
rect 218646 238506 218652 238508
rect 218513 238504 218652 238506
rect 218513 238448 218518 238504
rect 218574 238448 218652 238504
rect 218513 238446 218652 238448
rect 218513 238443 218579 238446
rect 218646 238444 218652 238446
rect 218716 238444 218722 238508
rect 218830 238172 218836 238236
rect 218900 238234 218906 238236
rect 219382 238234 219388 238236
rect 218900 238174 219388 238234
rect 218900 238172 218906 238174
rect 219382 238172 219388 238174
rect 219452 238172 219458 238236
rect 104801 238098 104867 238101
rect 225505 238098 225571 238101
rect 104801 238096 225571 238098
rect 104801 238040 104806 238096
rect 104862 238040 225510 238096
rect 225566 238040 225571 238096
rect 104801 238038 225571 238040
rect 104801 238035 104867 238038
rect 225505 238035 225571 238038
rect 57053 237962 57119 237965
rect 357433 237962 357499 237965
rect 57053 237960 357499 237962
rect 57053 237904 57058 237960
rect 57114 237904 357438 237960
rect 357494 237904 357499 237960
rect 57053 237902 357499 237904
rect 57053 237899 57119 237902
rect 357433 237899 357499 237902
rect 198457 236874 198523 236877
rect 226742 236874 226748 236876
rect 198457 236872 226748 236874
rect 198457 236816 198462 236872
rect 198518 236816 226748 236872
rect 198457 236814 226748 236816
rect 198457 236811 198523 236814
rect 226742 236812 226748 236814
rect 226812 236812 226818 236876
rect 122649 236738 122715 236741
rect 196525 236738 196591 236741
rect 122649 236736 196591 236738
rect 122649 236680 122654 236736
rect 122710 236680 196530 236736
rect 196586 236680 196591 236736
rect 122649 236678 196591 236680
rect 122649 236675 122715 236678
rect 196525 236675 196591 236678
rect 198641 236738 198707 236741
rect 227069 236738 227135 236741
rect 198641 236736 227135 236738
rect 198641 236680 198646 236736
rect 198702 236680 227074 236736
rect 227130 236680 227135 236736
rect 198641 236678 227135 236680
rect 198641 236675 198707 236678
rect 227069 236675 227135 236678
rect 58249 236602 58315 236605
rect 198733 236602 198799 236605
rect 58249 236600 198799 236602
rect 58249 236544 58254 236600
rect 58310 236544 198738 236600
rect 198794 236544 198799 236600
rect 58249 236542 198799 236544
rect 58249 236539 58315 236542
rect 198733 236539 198799 236542
rect 80605 236330 80671 236333
rect 86217 236330 86283 236333
rect 80605 236328 86283 236330
rect 80605 236272 80610 236328
rect 80666 236272 86222 236328
rect 86278 236272 86283 236328
rect 80605 236270 86283 236272
rect 80605 236267 80671 236270
rect 86217 236267 86283 236270
rect 217685 235922 217751 235925
rect 220077 235922 220143 235925
rect 217685 235920 220143 235922
rect 217685 235864 217690 235920
rect 217746 235864 220082 235920
rect 220138 235864 220143 235920
rect 217685 235862 220143 235864
rect 217685 235859 217751 235862
rect 220077 235859 220143 235862
rect 219198 235316 219204 235380
rect 219268 235378 219274 235380
rect 226558 235378 226564 235380
rect 219268 235318 226564 235378
rect 219268 235316 219274 235318
rect 226558 235316 226564 235318
rect 226628 235316 226634 235380
rect 4153 235242 4219 235245
rect 156045 235242 156111 235245
rect 4153 235240 156111 235242
rect 4153 235184 4158 235240
rect 4214 235184 156050 235240
rect 156106 235184 156111 235240
rect 4153 235182 156111 235184
rect 4153 235179 4219 235182
rect 156045 235179 156111 235182
rect 203517 235242 203583 235245
rect 226609 235242 226675 235245
rect 203517 235240 226675 235242
rect 203517 235184 203522 235240
rect 203578 235184 226614 235240
rect 226670 235184 226675 235240
rect 203517 235182 226675 235184
rect 203517 235179 203583 235182
rect 226609 235179 226675 235182
rect 218513 235106 218579 235109
rect 219198 235106 219204 235108
rect 218513 235104 219204 235106
rect 218513 235048 218518 235104
rect 218574 235048 219204 235104
rect 218513 235046 219204 235048
rect 218513 235043 218579 235046
rect 219198 235044 219204 235046
rect 219268 235044 219274 235108
rect 76557 234834 76623 234837
rect 205633 234834 205699 234837
rect 76557 234832 205699 234834
rect 76557 234776 76562 234832
rect 76618 234776 205638 234832
rect 205694 234776 205699 234832
rect 76557 234774 205699 234776
rect 76557 234771 76623 234774
rect 205633 234771 205699 234774
rect 73613 234698 73679 234701
rect 229737 234698 229803 234701
rect 73613 234696 229803 234698
rect 73613 234640 73618 234696
rect 73674 234640 229742 234696
rect 229798 234640 229803 234696
rect 73613 234638 229803 234640
rect 73613 234635 73679 234638
rect 229737 234635 229803 234638
rect 218646 234228 218652 234292
rect 218716 234290 218722 234292
rect 226190 234290 226196 234292
rect 218716 234230 226196 234290
rect 218716 234228 218722 234230
rect 226190 234228 226196 234230
rect 226260 234228 226266 234292
rect 218830 234092 218836 234156
rect 218900 234154 218906 234156
rect 226006 234154 226012 234156
rect 218900 234094 226012 234154
rect 218900 234092 218906 234094
rect 226006 234092 226012 234094
rect 226076 234092 226082 234156
rect 219801 234018 219867 234021
rect 227161 234018 227227 234021
rect 219801 234016 227227 234018
rect 219801 233960 219806 234016
rect 219862 233960 227166 234016
rect 227222 233960 227227 234016
rect 219801 233958 227227 233960
rect 219801 233955 219867 233958
rect 227161 233955 227227 233958
rect 101121 233882 101187 233885
rect 102041 233882 102107 233885
rect 101121 233880 102107 233882
rect 101121 233824 101126 233880
rect 101182 233824 102046 233880
rect 102102 233824 102107 233880
rect 101121 233822 102107 233824
rect 101121 233819 101187 233822
rect 102041 233819 102107 233822
rect 104065 233882 104131 233885
rect 104709 233882 104775 233885
rect 104065 233880 104775 233882
rect 104065 233824 104070 233880
rect 104126 233824 104714 233880
rect 104770 233824 104775 233880
rect 104065 233822 104775 233824
rect 104065 233819 104131 233822
rect 104709 233819 104775 233822
rect 114921 233882 114987 233885
rect 115841 233882 115907 233885
rect 114921 233880 115907 233882
rect 114921 233824 114926 233880
rect 114982 233824 115846 233880
rect 115902 233824 115907 233880
rect 114921 233822 115907 233824
rect 114921 233819 114987 233822
rect 115841 233819 115907 233822
rect 174169 233882 174235 233885
rect 175181 233882 175247 233885
rect 174169 233880 175247 233882
rect 174169 233824 174174 233880
rect 174230 233824 175186 233880
rect 175242 233824 175247 233880
rect 174169 233822 175247 233824
rect 174169 233819 174235 233822
rect 175181 233819 175247 233822
rect 187969 233882 188035 233885
rect 188981 233882 189047 233885
rect 187969 233880 189047 233882
rect 187969 233824 187974 233880
rect 188030 233824 188986 233880
rect 189042 233824 189047 233880
rect 187969 233822 189047 233824
rect 187969 233819 188035 233822
rect 188981 233819 189047 233822
rect 190913 233882 190979 233885
rect 191741 233882 191807 233885
rect 190913 233880 191807 233882
rect 190913 233824 190918 233880
rect 190974 233824 191746 233880
rect 191802 233824 191807 233880
rect 190913 233822 191807 233824
rect 190913 233819 190979 233822
rect 191741 233819 191807 233822
rect 201769 233882 201835 233885
rect 202781 233882 202847 233885
rect 201769 233880 202847 233882
rect 201769 233824 201774 233880
rect 201830 233824 202786 233880
rect 202842 233824 202847 233880
rect 201769 233822 202847 233824
rect 201769 233819 201835 233822
rect 202781 233819 202847 233822
rect 215569 233882 215635 233885
rect 216581 233882 216647 233885
rect 215569 233880 216647 233882
rect 215569 233824 215574 233880
rect 215630 233824 216586 233880
rect 216642 233824 216647 233880
rect 215569 233822 216647 233824
rect 215569 233819 215635 233822
rect 216581 233819 216647 233822
rect 217133 233882 217199 233885
rect 229461 233882 229527 233885
rect 217133 233880 229527 233882
rect 217133 233824 217138 233880
rect 217194 233824 229466 233880
rect 229522 233824 229527 233880
rect 217133 233822 229527 233824
rect 217133 233819 217199 233822
rect 229461 233819 229527 233822
rect 21357 233746 21423 233749
rect 164601 233746 164667 233749
rect 21357 233744 164667 233746
rect 21357 233688 21362 233744
rect 21418 233688 164606 233744
rect 164662 233688 164667 233744
rect 21357 233686 164667 233688
rect 21357 233683 21423 233686
rect 164601 233683 164667 233686
rect 18597 233610 18663 233613
rect 161657 233610 161723 233613
rect 18597 233608 161723 233610
rect 18597 233552 18602 233608
rect 18658 233552 161662 233608
rect 161718 233552 161723 233608
rect 18597 233550 161723 233552
rect 18597 233547 18663 233550
rect 161657 233547 161723 233550
rect 67541 233474 67607 233477
rect 228214 233474 228220 233476
rect 67541 233472 228220 233474
rect 67541 233416 67546 233472
rect 67602 233416 228220 233472
rect 67541 233414 228220 233416
rect 67541 233411 67607 233414
rect 228214 233412 228220 233414
rect 228284 233412 228290 233476
rect 64781 233338 64847 233341
rect 242433 233338 242499 233341
rect 64781 233336 242499 233338
rect 64781 233280 64786 233336
rect 64842 233280 242438 233336
rect 242494 233280 242499 233336
rect 64781 233278 242499 233280
rect 64781 233275 64847 233278
rect 242433 233275 242499 233278
rect 58617 232794 58683 232797
rect 125133 232794 125199 232797
rect 58617 232792 125199 232794
rect 58617 232736 58622 232792
rect 58678 232736 125138 232792
rect 125194 232736 125199 232792
rect 58617 232734 125199 232736
rect 58617 232731 58683 232734
rect 125133 232731 125199 232734
rect 146201 232794 146267 232797
rect 225781 232794 225847 232797
rect 146201 232792 225847 232794
rect 146201 232736 146206 232792
rect 146262 232736 225786 232792
rect 225842 232736 225847 232792
rect 146201 232734 225847 232736
rect 146201 232731 146267 232734
rect 225781 232731 225847 232734
rect 58157 232658 58223 232661
rect 91093 232658 91159 232661
rect 58157 232656 91159 232658
rect 58157 232600 58162 232656
rect 58218 232600 91098 232656
rect 91154 232600 91159 232656
rect 58157 232598 91159 232600
rect 58157 232595 58223 232598
rect 91093 232595 91159 232598
rect 105997 232658 106063 232661
rect 225689 232658 225755 232661
rect 105997 232656 225755 232658
rect 105997 232600 106002 232656
rect 106058 232600 225694 232656
rect 225750 232600 225755 232656
rect 105997 232598 225755 232600
rect 105997 232595 106063 232598
rect 225689 232595 225755 232598
rect 85481 232522 85547 232525
rect 225597 232522 225663 232525
rect 85481 232520 225663 232522
rect 85481 232464 85486 232520
rect 85542 232464 225602 232520
rect 225658 232464 225663 232520
rect 85481 232462 225663 232464
rect 85481 232459 85547 232462
rect 225597 232459 225663 232462
rect 583520 232386 584960 232476
rect 583342 232326 584960 232386
rect 583342 232250 583402 232326
rect 583520 232250 584960 232326
rect 583342 232236 584960 232250
rect 583342 232190 583586 232236
rect 72693 232114 72759 232117
rect 235533 232114 235599 232117
rect 72693 232112 235599 232114
rect 72693 232056 72698 232112
rect 72754 232056 235538 232112
rect 235594 232056 235599 232112
rect 72693 232054 235599 232056
rect 72693 232051 72759 232054
rect 235533 232051 235599 232054
rect 14457 231978 14523 231981
rect 166993 231978 167059 231981
rect 14457 231976 167059 231978
rect 14457 231920 14462 231976
rect 14518 231920 166998 231976
rect 167054 231920 167059 231976
rect 14457 231918 167059 231920
rect 14457 231915 14523 231918
rect 166993 231915 167059 231918
rect 205633 231978 205699 231981
rect 583526 231978 583586 232190
rect 205633 231976 583586 231978
rect 205633 231920 205638 231976
rect 205694 231920 583586 231976
rect 205633 231918 583586 231920
rect 205633 231915 205699 231918
rect 218881 231842 218947 231845
rect 224902 231842 224908 231844
rect 218881 231840 224908 231842
rect 218881 231784 218886 231840
rect 218942 231784 224908 231840
rect 218881 231782 224908 231784
rect 218881 231779 218947 231782
rect 224902 231780 224908 231782
rect 224972 231780 224978 231844
rect 218145 231706 218211 231709
rect 224718 231706 224724 231708
rect 218145 231704 224724 231706
rect 218145 231648 218150 231704
rect 218206 231648 224724 231704
rect 218145 231646 224724 231648
rect 218145 231643 218211 231646
rect 224718 231644 224724 231646
rect 224788 231644 224794 231708
rect 219249 231570 219315 231573
rect 226333 231570 226399 231573
rect 219249 231568 226399 231570
rect 219249 231512 219254 231568
rect 219310 231512 226338 231568
rect 226394 231512 226399 231568
rect 219249 231510 226399 231512
rect 219249 231507 219315 231510
rect 226333 231507 226399 231510
rect 218329 231434 218395 231437
rect 225873 231434 225939 231437
rect 218329 231432 225939 231434
rect 218329 231376 218334 231432
rect 218390 231376 225878 231432
rect 225934 231376 225939 231432
rect 218329 231374 225939 231376
rect 218329 231371 218395 231374
rect 225873 231371 225939 231374
rect 202137 231298 202203 231301
rect 226793 231298 226859 231301
rect 202137 231296 226859 231298
rect 202137 231240 202142 231296
rect 202198 231240 226798 231296
rect 226854 231240 226859 231296
rect 202137 231238 226859 231240
rect 202137 231235 202203 231238
rect 226793 231235 226859 231238
rect 11697 231162 11763 231165
rect 164049 231162 164115 231165
rect 11697 231160 164115 231162
rect 11697 231104 11702 231160
rect 11758 231104 164054 231160
rect 164110 231104 164115 231160
rect 11697 231102 164115 231104
rect 11697 231099 11763 231102
rect 164049 231099 164115 231102
rect 198273 231162 198339 231165
rect 226701 231162 226767 231165
rect 198273 231160 226767 231162
rect 198273 231104 198278 231160
rect 198334 231104 226706 231160
rect 226762 231104 226767 231160
rect 198273 231102 226767 231104
rect 198273 231099 198339 231102
rect 226701 231099 226767 231102
rect 7557 231026 7623 231029
rect 161013 231026 161079 231029
rect 7557 231024 161079 231026
rect 7557 230968 7562 231024
rect 7618 230968 161018 231024
rect 161074 230968 161079 231024
rect 7557 230966 161079 230968
rect 7557 230963 7623 230966
rect 161013 230963 161079 230966
rect 218421 231026 218487 231029
rect 223982 231026 223988 231028
rect 218421 231024 223988 231026
rect 218421 230968 218426 231024
rect 218482 230968 223988 231024
rect 218421 230966 223988 230968
rect 218421 230963 218487 230966
rect 223982 230964 223988 230966
rect 224052 230964 224058 231028
rect 4797 230890 4863 230893
rect 158069 230890 158135 230893
rect 4797 230888 158135 230890
rect 4797 230832 4802 230888
rect 4858 230832 158074 230888
rect 158130 230832 158135 230888
rect 4797 230830 158135 230832
rect 4797 230827 4863 230830
rect 158069 230827 158135 230830
rect 219198 230828 219204 230892
rect 219268 230890 219274 230892
rect 223798 230890 223804 230892
rect 219268 230830 223804 230890
rect 219268 230828 219274 230830
rect 223798 230828 223804 230830
rect 223868 230828 223874 230892
rect 15837 230754 15903 230757
rect 169937 230754 170003 230757
rect 15837 230752 170003 230754
rect 15837 230696 15842 230752
rect 15898 230696 169942 230752
rect 169998 230696 170003 230752
rect 15837 230694 170003 230696
rect 15837 230691 15903 230694
rect 169937 230691 170003 230694
rect 69289 230618 69355 230621
rect 260097 230618 260163 230621
rect 69289 230616 260163 230618
rect 69289 230560 69294 230616
rect 69350 230560 260102 230616
rect 260158 230560 260163 230616
rect 69289 230558 260163 230560
rect 69289 230555 69355 230558
rect 260097 230555 260163 230558
rect 128353 230482 128419 230485
rect 129181 230482 129247 230485
rect 128353 230480 129247 230482
rect 128353 230424 128358 230480
rect 128414 230424 129186 230480
rect 129242 230424 129247 230480
rect 128353 230422 129247 230424
rect 128353 230419 128419 230422
rect 129181 230419 129247 230422
rect 131113 230482 131179 230485
rect 132125 230482 132191 230485
rect 131113 230480 132191 230482
rect 131113 230424 131118 230480
rect 131174 230424 132130 230480
rect 132186 230424 132191 230480
rect 131113 230422 132191 230424
rect 131113 230419 131179 230422
rect 132125 230419 132191 230422
rect 135253 230482 135319 230485
rect 135989 230482 136055 230485
rect 135253 230480 136055 230482
rect 135253 230424 135258 230480
rect 135314 230424 135994 230480
rect 136050 230424 136055 230480
rect 135253 230422 136055 230424
rect 135253 230419 135319 230422
rect 135989 230419 136055 230422
rect 138013 230482 138079 230485
rect 138933 230482 138999 230485
rect 138013 230480 138999 230482
rect 138013 230424 138018 230480
rect 138074 230424 138938 230480
rect 138994 230424 138999 230480
rect 138013 230422 138999 230424
rect 138013 230419 138079 230422
rect 138933 230419 138999 230422
rect 142153 230482 142219 230485
rect 142981 230482 143047 230485
rect 142153 230480 143047 230482
rect 142153 230424 142158 230480
rect 142214 230424 142986 230480
rect 143042 230424 143047 230480
rect 142153 230422 143047 230424
rect 142153 230419 142219 230422
rect 142981 230419 143047 230422
rect 146293 230482 146359 230485
rect 146845 230482 146911 230485
rect 146293 230480 146911 230482
rect 146293 230424 146298 230480
rect 146354 230424 146850 230480
rect 146906 230424 146911 230480
rect 146293 230422 146911 230424
rect 146293 230419 146359 230422
rect 146845 230419 146911 230422
rect 153193 230482 153259 230485
rect 153837 230482 153903 230485
rect 153193 230480 153903 230482
rect 153193 230424 153198 230480
rect 153254 230424 153842 230480
rect 153898 230424 153903 230480
rect 153193 230422 153903 230424
rect 153193 230419 153259 230422
rect 153837 230419 153903 230422
rect 211337 230482 211403 230485
rect 213177 230482 213243 230485
rect 211337 230480 213243 230482
rect 211337 230424 211342 230480
rect 211398 230424 213182 230480
rect 213238 230424 213243 230480
rect 211337 230422 213243 230424
rect 211337 230419 211403 230422
rect 213177 230419 213243 230422
rect 63401 230346 63467 230349
rect 242341 230346 242407 230349
rect 63401 230344 242407 230346
rect 63401 230288 63406 230344
rect 63462 230288 242346 230344
rect 242402 230288 242407 230344
rect 63401 230286 242407 230288
rect 63401 230283 63467 230286
rect 242341 230283 242407 230286
rect 183737 230210 183803 230213
rect 196709 230210 196775 230213
rect 183737 230208 196775 230210
rect 183737 230152 183742 230208
rect 183798 230152 196714 230208
rect 196770 230152 196775 230208
rect 183737 230150 196775 230152
rect 183737 230147 183803 230150
rect 196709 230147 196775 230150
rect 184749 230074 184815 230077
rect 198365 230074 198431 230077
rect 184749 230072 198431 230074
rect 184749 230016 184754 230072
rect 184810 230016 198370 230072
rect 198426 230016 198431 230072
rect 184749 230014 198431 230016
rect 184749 230011 184815 230014
rect 198365 230011 198431 230014
rect 219065 230074 219131 230077
rect 223205 230074 223271 230077
rect 219065 230072 223271 230074
rect 219065 230016 219070 230072
rect 219126 230016 223210 230072
rect 223266 230016 223271 230072
rect 219065 230014 223271 230016
rect 219065 230011 219131 230014
rect 223205 230011 223271 230014
rect 59997 229938 60063 229941
rect 127525 229938 127591 229941
rect 163037 229938 163103 229941
rect 59997 229936 127591 229938
rect 59997 229880 60002 229936
rect 60058 229880 127530 229936
rect 127586 229880 127591 229936
rect 59997 229878 127591 229880
rect 59997 229875 60063 229878
rect 127525 229875 127591 229878
rect 137970 229936 163103 229938
rect 137970 229880 163042 229936
rect 163098 229880 163103 229936
rect 137970 229878 163103 229880
rect 74533 229802 74599 229805
rect 137970 229802 138030 229878
rect 163037 229875 163103 229878
rect 182725 229938 182791 229941
rect 198549 229938 198615 229941
rect 182725 229936 198615 229938
rect 182725 229880 182730 229936
rect 182786 229880 198554 229936
rect 198610 229880 198615 229936
rect 182725 229878 198615 229880
rect 182725 229875 182791 229878
rect 198549 229875 198615 229878
rect 217961 229938 218027 229941
rect 230749 229938 230815 229941
rect 217961 229936 230815 229938
rect 217961 229880 217966 229936
rect 218022 229880 230754 229936
rect 230810 229880 230815 229936
rect 217961 229878 230815 229880
rect 217961 229875 218027 229878
rect 230749 229875 230815 229878
rect 160185 229802 160251 229805
rect 74533 229800 138030 229802
rect 74533 229744 74538 229800
rect 74594 229744 138030 229800
rect 74533 229742 138030 229744
rect 147630 229800 160251 229802
rect 147630 229744 160190 229800
rect 160246 229744 160251 229800
rect 147630 229742 160251 229744
rect 74533 229739 74599 229742
rect 70301 229666 70367 229669
rect 147630 229666 147690 229742
rect 160185 229739 160251 229742
rect 179781 229802 179847 229805
rect 196801 229802 196867 229805
rect 179781 229800 196867 229802
rect 179781 229744 179786 229800
rect 179842 229744 196806 229800
rect 196862 229744 196867 229800
rect 179781 229742 196867 229744
rect 179781 229739 179847 229742
rect 196801 229739 196867 229742
rect 198089 229802 198155 229805
rect 227437 229802 227503 229805
rect 198089 229800 227503 229802
rect 198089 229744 198094 229800
rect 198150 229744 227442 229800
rect 227498 229744 227503 229800
rect 198089 229742 227503 229744
rect 198089 229739 198155 229742
rect 227437 229739 227503 229742
rect 70301 229664 147690 229666
rect 70301 229608 70306 229664
rect 70362 229608 147690 229664
rect 70301 229606 147690 229608
rect 160093 229666 160159 229669
rect 167913 229666 167979 229669
rect 160093 229664 167979 229666
rect 160093 229608 160098 229664
rect 160154 229608 167918 229664
rect 167974 229608 167979 229664
rect 160093 229606 167979 229608
rect 70301 229603 70367 229606
rect 160093 229603 160159 229606
rect 167913 229603 167979 229606
rect 25497 229530 25563 229533
rect 165981 229530 166047 229533
rect 25497 229528 166047 229530
rect 25497 229472 25502 229528
rect 25558 229472 165986 229528
rect 166042 229472 166047 229528
rect 25497 229470 166047 229472
rect 25497 229467 25563 229470
rect 165981 229467 166047 229470
rect 29637 229394 29703 229397
rect 171869 229394 171935 229397
rect 29637 229392 171935 229394
rect 29637 229336 29642 229392
rect 29698 229336 171874 229392
rect 171930 229336 171935 229392
rect 29637 229334 171935 229336
rect 29637 229331 29703 229334
rect 171869 229331 171935 229334
rect 66345 229258 66411 229261
rect 224585 229258 224651 229261
rect 66345 229256 224651 229258
rect 66345 229200 66350 229256
rect 66406 229200 224590 229256
rect 224646 229200 224651 229256
rect 66345 229198 224651 229200
rect 66345 229195 66411 229198
rect 224585 229195 224651 229198
rect 219014 228788 219020 228852
rect 219084 228850 219090 228852
rect 224166 228850 224172 228852
rect 219084 228790 224172 228850
rect 219084 228788 219090 228790
rect 224166 228788 224172 228790
rect 224236 228788 224242 228852
rect 218789 228714 218855 228717
rect 224350 228714 224356 228716
rect 218789 228712 224356 228714
rect 218789 228656 218794 228712
rect 218850 228656 224356 228712
rect 218789 228654 224356 228656
rect 218789 228651 218855 228654
rect 224350 228652 224356 228654
rect 224420 228652 224426 228716
rect 3601 228578 3667 228581
rect 70301 228578 70367 228581
rect 3601 228576 70367 228578
rect 3601 228520 3606 228576
rect 3662 228520 70306 228576
rect 70362 228520 70367 228576
rect 3601 228518 70367 228520
rect 3601 228515 3667 228518
rect 70301 228515 70367 228518
rect 219157 228578 219223 228581
rect 225270 228578 225276 228580
rect 219157 228576 225276 228578
rect 219157 228520 219162 228576
rect 219218 228520 225276 228576
rect 219157 228518 225276 228520
rect 219157 228515 219223 228518
rect 225270 228516 225276 228518
rect 225340 228516 225346 228580
rect 22737 228442 22803 228445
rect 170949 228442 171015 228445
rect 22737 228440 171015 228442
rect 22737 228384 22742 228440
rect 22798 228384 170954 228440
rect 171010 228384 171015 228440
rect 22737 228382 171015 228384
rect 22737 228379 22803 228382
rect 170949 228379 171015 228382
rect 219893 228442 219959 228445
rect 227529 228442 227595 228445
rect 219893 228440 227595 228442
rect 219893 228384 219898 228440
rect 219954 228384 227534 228440
rect 227590 228384 227595 228440
rect 219893 228382 227595 228384
rect 219893 228379 219959 228382
rect 227529 228379 227595 228382
rect 3417 228306 3483 228309
rect 160093 228306 160159 228309
rect 3417 228304 160159 228306
rect 3417 228248 3422 228304
rect 3478 228248 160098 228304
rect 160154 228248 160159 228304
rect 3417 228246 160159 228248
rect 3417 228243 3483 228246
rect 160093 228243 160159 228246
rect 199377 228306 199443 228309
rect 225965 228306 226031 228309
rect 199377 228304 226031 228306
rect 199377 228248 199382 228304
rect 199438 228248 225970 228304
rect 226026 228248 226031 228304
rect 199377 228246 226031 228248
rect 199377 228243 199443 228246
rect 225965 228243 226031 228246
rect 74257 228170 74323 228173
rect 239397 228170 239463 228173
rect 74257 228168 239463 228170
rect -960 227884 480 228124
rect 74257 228112 74262 228168
rect 74318 228112 239402 228168
rect 239458 228112 239463 228168
rect 74257 228110 239463 228112
rect 74257 228107 74323 228110
rect 239397 228107 239463 228110
rect 71221 228034 71287 228037
rect 236637 228034 236703 228037
rect 71221 228032 236703 228034
rect 71221 227976 71226 228032
rect 71282 227976 236642 228032
rect 236698 227976 236703 228032
rect 71221 227974 236703 227976
rect 71221 227971 71287 227974
rect 236637 227971 236703 227974
rect 65333 227898 65399 227901
rect 240777 227898 240843 227901
rect 65333 227896 240843 227898
rect 65333 227840 65338 227896
rect 65394 227840 240782 227896
rect 240838 227840 240843 227896
rect 65333 227838 240843 227840
rect 65333 227835 65399 227838
rect 240777 227835 240843 227838
rect 57789 227762 57855 227765
rect 62757 227762 62823 227765
rect 57789 227760 62823 227762
rect 57789 227704 57794 227760
rect 57850 227704 62762 227760
rect 62818 227704 62823 227760
rect 57789 227702 62823 227704
rect 57789 227699 57855 227702
rect 62757 227699 62823 227702
rect 70301 227762 70367 227765
rect 396717 227762 396783 227765
rect 70301 227760 396783 227762
rect 70301 227704 70306 227760
rect 70362 227704 396722 227760
rect 396778 227704 396783 227760
rect 70301 227702 396783 227704
rect 70301 227699 70367 227702
rect 396717 227699 396783 227702
rect 58617 227354 58683 227357
rect 75913 227354 75979 227357
rect 58617 227352 75979 227354
rect 58617 227296 58622 227352
rect 58678 227296 75918 227352
rect 75974 227296 75979 227352
rect 58617 227294 75979 227296
rect 58617 227291 58683 227294
rect 75913 227291 75979 227294
rect 3693 227218 3759 227221
rect 74533 227218 74599 227221
rect 3693 227216 74599 227218
rect 3693 227160 3698 227216
rect 3754 227160 74538 227216
rect 74594 227160 74599 227216
rect 3693 227158 74599 227160
rect 3693 227155 3759 227158
rect 74533 227155 74599 227158
rect 219341 227218 219407 227221
rect 227621 227218 227687 227221
rect 219341 227216 227687 227218
rect 219341 227160 219346 227216
rect 219402 227160 227626 227216
rect 227682 227160 227687 227216
rect 219341 227158 227687 227160
rect 219341 227155 219407 227158
rect 227621 227155 227687 227158
rect 3509 227082 3575 227085
rect 168557 227082 168623 227085
rect 3509 227080 168623 227082
rect 3509 227024 3514 227080
rect 3570 227024 168562 227080
rect 168618 227024 168623 227080
rect 3509 227022 168623 227024
rect 3509 227019 3575 227022
rect 168557 227019 168623 227022
rect 217409 227082 217475 227085
rect 227253 227082 227319 227085
rect 217409 227080 227319 227082
rect 217409 227024 217414 227080
rect 217470 227024 227258 227080
rect 227314 227024 227319 227080
rect 217409 227022 227319 227024
rect 217409 227019 217475 227022
rect 227253 227019 227319 227022
rect 61285 226946 61351 226949
rect 580257 226946 580323 226949
rect 61285 226944 580323 226946
rect 61285 226888 61290 226944
rect 61346 226888 580262 226944
rect 580318 226888 580323 226944
rect 61285 226886 580323 226888
rect 61285 226883 61351 226886
rect 580257 226883 580323 226886
rect 17217 226810 17283 226813
rect 158805 226810 158871 226813
rect 17217 226808 158871 226810
rect 17217 226752 17222 226808
rect 17278 226752 158810 226808
rect 158866 226752 158871 226808
rect 17217 226750 158871 226752
rect 17217 226747 17283 226750
rect 158805 226747 158871 226750
rect 181161 226810 181227 226813
rect 182081 226810 182147 226813
rect 181161 226808 182147 226810
rect 181161 226752 181166 226808
rect 181222 226752 182086 226808
rect 182142 226752 182147 226808
rect 181161 226750 182147 226752
rect 181161 226747 181227 226750
rect 182081 226747 182147 226750
rect 60590 226612 60596 226676
rect 60660 226674 60666 226676
rect 61101 226674 61167 226677
rect 60660 226672 61167 226674
rect 60660 226616 61106 226672
rect 61162 226616 61167 226672
rect 60660 226614 61167 226616
rect 60660 226612 60666 226614
rect 61101 226611 61167 226614
rect 77385 226674 77451 226677
rect 235625 226674 235691 226677
rect 77385 226672 235691 226674
rect 77385 226616 77390 226672
rect 77446 226616 235630 226672
rect 235686 226616 235691 226672
rect 77385 226614 235691 226616
rect 77385 226611 77451 226614
rect 235625 226611 235691 226614
rect 55673 226538 55739 226541
rect 62113 226538 62179 226541
rect 55673 226536 62179 226538
rect 55673 226480 55678 226536
rect 55734 226480 62118 226536
rect 62174 226480 62179 226536
rect 55673 226478 62179 226480
rect 55673 226475 55739 226478
rect 62113 226475 62179 226478
rect 75545 226538 75611 226541
rect 236729 226538 236795 226541
rect 75545 226536 236795 226538
rect 75545 226480 75550 226536
rect 75606 226480 236734 226536
rect 236790 226480 236795 226536
rect 75545 226478 236795 226480
rect 75545 226475 75611 226478
rect 236729 226475 236795 226478
rect 55765 226402 55831 226405
rect 60181 226402 60247 226405
rect 61745 226402 61811 226405
rect 55765 226400 60247 226402
rect 55765 226344 55770 226400
rect 55826 226344 60186 226400
rect 60242 226344 60247 226400
rect 55765 226342 60247 226344
rect 55765 226339 55831 226342
rect 60181 226339 60247 226342
rect 60598 226400 61811 226402
rect 60598 226344 61750 226400
rect 61806 226344 61811 226400
rect 60598 226342 61811 226344
rect 57697 226266 57763 226269
rect 60598 226266 60658 226342
rect 61745 226339 61811 226342
rect 68553 226402 68619 226405
rect 235441 226402 235507 226405
rect 68553 226400 235507 226402
rect 68553 226344 68558 226400
rect 68614 226344 235446 226400
rect 235502 226344 235507 226400
rect 68553 226342 235507 226344
rect 68553 226339 68619 226342
rect 235441 226339 235507 226342
rect 57697 226264 60658 226266
rect 57697 226208 57702 226264
rect 57758 226208 60658 226264
rect 57697 226206 60658 226208
rect 57697 226203 57763 226206
rect 60774 226204 60780 226268
rect 60844 226266 60850 226268
rect 61101 226266 61167 226269
rect 61929 226266 61995 226269
rect 60844 226264 61167 226266
rect 60844 226208 61106 226264
rect 61162 226208 61167 226264
rect 60844 226206 61167 226208
rect 60844 226204 60850 226206
rect 61101 226203 61167 226206
rect 61702 226264 61995 226266
rect 61702 226208 61934 226264
rect 61990 226208 61995 226264
rect 61702 226206 61995 226208
rect 57881 226130 57947 226133
rect 61702 226130 61762 226206
rect 61929 226203 61995 226206
rect 218697 226266 218763 226269
rect 220537 226266 220603 226269
rect 218697 226264 219450 226266
rect 218697 226208 218702 226264
rect 218758 226208 219450 226264
rect 218697 226206 219450 226208
rect 218697 226203 218763 226206
rect 57881 226128 61762 226130
rect 57881 226072 57886 226128
rect 57942 226072 61762 226128
rect 57881 226070 61762 226072
rect 57881 226067 57947 226070
rect 56777 225994 56843 225997
rect 60590 225994 60596 225996
rect 56777 225992 60596 225994
rect 56777 225936 56782 225992
rect 56838 225936 60596 225992
rect 56777 225934 60596 225936
rect 56777 225931 56843 225934
rect 60590 225932 60596 225934
rect 60660 225932 60666 225996
rect 60774 225858 60780 225860
rect 60598 225798 60780 225858
rect 60598 225284 60658 225798
rect 60774 225796 60780 225798
rect 60844 225796 60850 225860
rect 219390 225858 219450 226206
rect 220537 226264 220922 226266
rect 220537 226208 220542 226264
rect 220598 226208 220922 226264
rect 220537 226206 220922 226208
rect 220537 226203 220603 226206
rect 220862 226130 220922 226206
rect 223430 226204 223436 226268
rect 223500 226266 223506 226268
rect 223573 226266 223639 226269
rect 224585 226266 224651 226269
rect 223500 226264 223639 226266
rect 223500 226208 223578 226264
rect 223634 226208 223639 226264
rect 223500 226206 223639 226208
rect 223500 226204 223506 226206
rect 223573 226203 223639 226206
rect 223806 226206 224418 226266
rect 223806 226130 223866 226206
rect 220862 226070 223866 226130
rect 224358 226130 224418 226206
rect 224585 226264 229110 226266
rect 224585 226208 224590 226264
rect 224646 226208 229110 226264
rect 224585 226206 229110 226208
rect 224585 226203 224651 226206
rect 226885 226130 226951 226133
rect 224358 226128 226951 226130
rect 224358 226072 226890 226128
rect 226946 226072 226951 226128
rect 224358 226070 226951 226072
rect 226885 226067 226951 226070
rect 219390 225798 224234 225858
rect 223430 225660 223436 225724
rect 223500 225722 223506 225724
rect 224174 225722 224234 225798
rect 226926 225722 226932 225724
rect 223500 225662 224050 225722
rect 224174 225662 226932 225722
rect 223500 225660 223506 225662
rect 223990 225420 224050 225662
rect 226926 225660 226932 225662
rect 226996 225660 227002 225724
rect 229050 225722 229110 226206
rect 580349 225722 580415 225725
rect 229050 225720 580415 225722
rect 229050 225664 580354 225720
rect 580410 225664 580415 225720
rect 229050 225662 580415 225664
rect 580349 225659 580415 225662
rect 226333 222730 226399 222733
rect 224572 222728 226399 222730
rect 224572 222672 226338 222728
rect 226394 222672 226399 222728
rect 224572 222670 226399 222672
rect 226333 222667 226399 222670
rect 56225 222322 56291 222325
rect 56225 222320 60076 222322
rect 56225 222264 56230 222320
rect 56286 222264 60076 222320
rect 56225 222262 60076 222264
rect 56225 222259 56291 222262
rect 228909 220010 228975 220013
rect 224572 220008 228975 220010
rect 224572 219952 228914 220008
rect 228970 219952 228975 220008
rect 224572 219950 228975 219952
rect 228909 219947 228975 219950
rect 57789 219330 57855 219333
rect 57789 219328 60076 219330
rect 57789 219272 57794 219328
rect 57850 219272 60076 219328
rect 57789 219270 60076 219272
rect 57789 219267 57855 219270
rect 583520 219058 584960 219148
rect 583342 218998 584960 219058
rect 583342 218922 583402 218998
rect 583520 218922 584960 218998
rect 583342 218908 584960 218922
rect 583342 218862 583586 218908
rect 235625 218106 235691 218109
rect 583526 218106 583586 218862
rect 235625 218104 583586 218106
rect 235625 218048 235630 218104
rect 235686 218048 583586 218104
rect 235625 218046 583586 218048
rect 235625 218043 235691 218046
rect 230933 217290 230999 217293
rect 224572 217288 230999 217290
rect 224572 217232 230938 217288
rect 230994 217232 230999 217288
rect 224572 217230 230999 217232
rect 230933 217227 230999 217230
rect 56409 216338 56475 216341
rect 56409 216336 60076 216338
rect 56409 216280 56414 216336
rect 56470 216280 60076 216336
rect 56409 216278 60076 216280
rect 56409 216275 56475 216278
rect -960 214978 480 215068
rect 2773 214978 2839 214981
rect -960 214976 2839 214978
rect -960 214920 2778 214976
rect 2834 214920 2839 214976
rect -960 214918 2839 214920
rect -960 214828 480 214918
rect 2773 214915 2839 214918
rect 227529 214570 227595 214573
rect 224572 214568 227595 214570
rect 224572 214512 227534 214568
rect 227590 214512 227595 214568
rect 224572 214510 227595 214512
rect 227529 214507 227595 214510
rect 59445 213346 59511 213349
rect 59445 213344 60076 213346
rect 59445 213288 59450 213344
rect 59506 213288 60076 213344
rect 59445 213286 60076 213288
rect 59445 213283 59511 213286
rect 229001 211850 229067 211853
rect 224572 211848 229067 211850
rect 224572 211792 229006 211848
rect 229062 211792 229067 211848
rect 224572 211790 229067 211792
rect 229001 211787 229067 211790
rect 57513 210354 57579 210357
rect 57513 210352 60076 210354
rect 57513 210296 57518 210352
rect 57574 210296 60076 210352
rect 57513 210294 60076 210296
rect 57513 210291 57579 210294
rect 228817 209130 228883 209133
rect 224572 209128 228883 209130
rect 224572 209072 228822 209128
rect 228878 209072 228883 209128
rect 224572 209070 228883 209072
rect 228817 209067 228883 209070
rect 55857 207362 55923 207365
rect 55857 207360 60076 207362
rect 55857 207304 55862 207360
rect 55918 207304 60076 207360
rect 55857 207302 60076 207304
rect 55857 207299 55923 207302
rect 231301 206410 231367 206413
rect 224572 206408 231367 206410
rect 224572 206352 231306 206408
rect 231362 206352 231367 206408
rect 224572 206350 231367 206352
rect 231301 206347 231367 206350
rect 236729 205730 236795 205733
rect 583520 205730 584960 205820
rect 236729 205728 584960 205730
rect 236729 205672 236734 205728
rect 236790 205672 584960 205728
rect 236729 205670 584960 205672
rect 236729 205667 236795 205670
rect 583520 205580 584960 205670
rect 58709 204370 58775 204373
rect 58709 204368 60076 204370
rect 58709 204312 58714 204368
rect 58770 204312 60076 204368
rect 58709 204310 60076 204312
rect 58709 204307 58775 204310
rect 226333 204234 226399 204237
rect 242249 204234 242315 204237
rect 226333 204232 242315 204234
rect 226333 204176 226338 204232
rect 226394 204176 242254 204232
rect 242310 204176 242315 204232
rect 226333 204174 242315 204176
rect 226333 204171 226399 204174
rect 242249 204171 242315 204174
rect 226333 203554 226399 203557
rect 224572 203552 226399 203554
rect 224572 203496 226338 203552
rect 226394 203496 226399 203552
rect 224572 203494 226399 203496
rect 226333 203491 226399 203494
rect -960 201922 480 202012
rect 3601 201922 3667 201925
rect -960 201920 3667 201922
rect -960 201864 3606 201920
rect 3662 201864 3667 201920
rect -960 201862 3667 201864
rect -960 201772 480 201862
rect 3601 201859 3667 201862
rect 58433 201378 58499 201381
rect 58433 201376 60076 201378
rect 58433 201320 58438 201376
rect 58494 201320 60076 201376
rect 58433 201318 60076 201320
rect 58433 201315 58499 201318
rect 227437 200834 227503 200837
rect 224572 200832 227503 200834
rect 224572 200776 227442 200832
rect 227498 200776 227503 200832
rect 224572 200774 227503 200776
rect 227437 200771 227503 200774
rect 57881 198386 57947 198389
rect 57881 198384 60076 198386
rect 57881 198328 57886 198384
rect 57942 198328 60076 198384
rect 57881 198326 60076 198328
rect 57881 198323 57947 198326
rect 227621 198114 227687 198117
rect 224572 198112 227687 198114
rect 224572 198056 227626 198112
rect 227682 198056 227687 198112
rect 224572 198054 227687 198056
rect 227621 198051 227687 198054
rect 57513 195394 57579 195397
rect 238109 195394 238175 195397
rect 57513 195392 60076 195394
rect 57513 195336 57518 195392
rect 57574 195336 60076 195392
rect 57513 195334 60076 195336
rect 224572 195392 238175 195394
rect 224572 195336 238114 195392
rect 238170 195336 238175 195392
rect 224572 195334 238175 195336
rect 57513 195331 57579 195334
rect 238109 195331 238175 195334
rect 227161 192674 227227 192677
rect 224572 192672 227227 192674
rect 224572 192616 227166 192672
rect 227222 192616 227227 192672
rect 224572 192614 227227 192616
rect 227161 192611 227227 192614
rect 57513 192538 57579 192541
rect 583520 192538 584960 192628
rect 57513 192536 60076 192538
rect 57513 192480 57518 192536
rect 57574 192480 60076 192536
rect 57513 192478 60076 192480
rect 583342 192478 584960 192538
rect 57513 192475 57579 192478
rect 583342 192402 583402 192478
rect 583520 192402 584960 192478
rect 583342 192388 584960 192402
rect 583342 192342 583586 192388
rect 229737 191858 229803 191861
rect 583526 191858 583586 192342
rect 229737 191856 583586 191858
rect 229737 191800 229742 191856
rect 229798 191800 583586 191856
rect 229737 191798 583586 191800
rect 229737 191795 229803 191798
rect 229553 189954 229619 189957
rect 224572 189952 229619 189954
rect 224572 189896 229558 189952
rect 229614 189896 229619 189952
rect 224572 189894 229619 189896
rect 229553 189891 229619 189894
rect 55949 189546 56015 189549
rect 55949 189544 60076 189546
rect 55949 189488 55954 189544
rect 56010 189488 60076 189544
rect 55949 189486 60076 189488
rect 55949 189483 56015 189486
rect -960 188866 480 188956
rect 3141 188866 3207 188869
rect -960 188864 3207 188866
rect -960 188808 3146 188864
rect 3202 188808 3207 188864
rect -960 188806 3207 188808
rect -960 188716 480 188806
rect 3141 188803 3207 188806
rect 227253 187234 227319 187237
rect 224572 187232 227319 187234
rect 224572 187176 227258 187232
rect 227314 187176 227319 187232
rect 224572 187174 227319 187176
rect 227253 187171 227319 187174
rect 57237 186554 57303 186557
rect 57237 186552 60076 186554
rect 57237 186496 57242 186552
rect 57298 186496 60076 186552
rect 57237 186494 60076 186496
rect 57237 186491 57303 186494
rect 233969 184514 234035 184517
rect 224572 184512 234035 184514
rect 224572 184456 233974 184512
rect 234030 184456 234035 184512
rect 224572 184454 234035 184456
rect 233969 184451 234035 184454
rect 57513 183562 57579 183565
rect 57513 183560 60076 183562
rect 57513 183504 57518 183560
rect 57574 183504 60076 183560
rect 57513 183502 60076 183504
rect 57513 183499 57579 183502
rect 226517 181794 226583 181797
rect 224572 181792 226583 181794
rect 224572 181736 226522 181792
rect 226578 181736 226583 181792
rect 224572 181734 226583 181736
rect 226517 181731 226583 181734
rect 58893 180570 58959 180573
rect 58893 180568 60076 180570
rect 58893 180512 58898 180568
rect 58954 180512 60076 180568
rect 58893 180510 60076 180512
rect 58893 180507 58959 180510
rect 583520 179210 584960 179300
rect 583342 179150 584960 179210
rect 583342 179074 583402 179150
rect 583520 179074 584960 179150
rect 583342 179060 584960 179074
rect 583342 179014 583586 179060
rect 230841 178938 230907 178941
rect 224572 178936 230907 178938
rect 224572 178880 230846 178936
rect 230902 178880 230907 178936
rect 224572 178878 230907 178880
rect 230841 178875 230907 178878
rect 239397 178122 239463 178125
rect 583526 178122 583586 179014
rect 239397 178120 583586 178122
rect 239397 178064 239402 178120
rect 239458 178064 583586 178120
rect 239397 178062 583586 178064
rect 239397 178059 239463 178062
rect 56041 177578 56107 177581
rect 56041 177576 60076 177578
rect 56041 177520 56046 177576
rect 56102 177520 60076 177576
rect 56041 177518 60076 177520
rect 56041 177515 56107 177518
rect 227069 176218 227135 176221
rect 224572 176216 227135 176218
rect 224572 176160 227074 176216
rect 227130 176160 227135 176216
rect 224572 176158 227135 176160
rect 227069 176155 227135 176158
rect -960 175796 480 176036
rect 58985 174586 59051 174589
rect 58985 174584 60076 174586
rect 58985 174528 58990 174584
rect 59046 174528 60076 174584
rect 58985 174526 60076 174528
rect 58985 174523 59051 174526
rect 232405 173498 232471 173501
rect 224572 173496 232471 173498
rect 224572 173440 232410 173496
rect 232466 173440 232471 173496
rect 224572 173438 232471 173440
rect 232405 173435 232471 173438
rect 56777 171594 56843 171597
rect 56777 171592 60076 171594
rect 56777 171536 56782 171592
rect 56838 171536 60076 171592
rect 56777 171534 60076 171536
rect 56777 171531 56843 171534
rect 240869 171050 240935 171053
rect 229050 171048 240935 171050
rect 229050 170992 240874 171048
rect 240930 170992 240935 171048
rect 229050 170990 240935 170992
rect 229050 170778 229110 170990
rect 240869 170987 240935 170990
rect 224572 170718 229110 170778
rect 57789 168602 57855 168605
rect 57789 168600 60076 168602
rect 57789 168544 57794 168600
rect 57850 168544 60076 168600
rect 57789 168542 60076 168544
rect 57789 168539 57855 168542
rect 226977 168058 227043 168061
rect 224572 168056 227043 168058
rect 224572 168000 226982 168056
rect 227038 168000 227043 168056
rect 224572 167998 227043 168000
rect 226977 167995 227043 167998
rect 583520 165882 584960 165972
rect 567150 165822 584960 165882
rect 235533 165746 235599 165749
rect 567150 165746 567210 165822
rect 235533 165744 567210 165746
rect 235533 165688 235538 165744
rect 235594 165688 567210 165744
rect 583520 165732 584960 165822
rect 235533 165686 567210 165688
rect 235533 165683 235599 165686
rect 58525 165610 58591 165613
rect 58525 165608 60076 165610
rect 58525 165552 58530 165608
rect 58586 165552 60076 165608
rect 58525 165550 60076 165552
rect 58525 165547 58591 165550
rect 228541 165338 228607 165341
rect 224572 165336 228607 165338
rect 224572 165280 228546 165336
rect 228602 165280 228607 165336
rect 224572 165278 228607 165280
rect 228541 165275 228607 165278
rect -960 162890 480 162980
rect 3325 162890 3391 162893
rect -960 162888 3391 162890
rect -960 162832 3330 162888
rect 3386 162832 3391 162888
rect -960 162830 3391 162832
rect -960 162740 480 162830
rect 3325 162827 3391 162830
rect 57421 162618 57487 162621
rect 228449 162618 228515 162621
rect 57421 162616 60076 162618
rect 57421 162560 57426 162616
rect 57482 162560 60076 162616
rect 57421 162558 60076 162560
rect 224572 162616 228515 162618
rect 224572 162560 228454 162616
rect 228510 162560 228515 162616
rect 224572 162558 228515 162560
rect 57421 162555 57487 162558
rect 228449 162555 228515 162558
rect 231209 159898 231275 159901
rect 224572 159896 231275 159898
rect 224572 159840 231214 159896
rect 231270 159840 231275 159896
rect 224572 159838 231275 159840
rect 231209 159835 231275 159838
rect 57789 159762 57855 159765
rect 57789 159760 60076 159762
rect 57789 159704 57794 159760
rect 57850 159704 60076 159760
rect 57789 159702 60076 159704
rect 57789 159699 57855 159702
rect 228725 157178 228791 157181
rect 224572 157176 228791 157178
rect 224572 157120 228730 157176
rect 228786 157120 228791 157176
rect 224572 157118 228791 157120
rect 228725 157115 228791 157118
rect 57421 156770 57487 156773
rect 57421 156768 60076 156770
rect 57421 156712 57426 156768
rect 57482 156712 60076 156768
rect 57421 156710 60076 156712
rect 57421 156707 57487 156710
rect 226885 154322 226951 154325
rect 224572 154320 226951 154322
rect 224572 154264 226890 154320
rect 226946 154264 226951 154320
rect 224572 154262 226951 154264
rect 226885 154259 226951 154262
rect 57421 153778 57487 153781
rect 57421 153776 60076 153778
rect 57421 153720 57426 153776
rect 57482 153720 60076 153776
rect 57421 153718 60076 153720
rect 57421 153715 57487 153718
rect 579613 152690 579679 152693
rect 583520 152690 584960 152780
rect 579613 152688 584960 152690
rect 579613 152632 579618 152688
rect 579674 152632 584960 152688
rect 579613 152630 584960 152632
rect 579613 152627 579679 152630
rect 583520 152540 584960 152630
rect 226793 151602 226859 151605
rect 224572 151600 226859 151602
rect 224572 151544 226798 151600
rect 226854 151544 226859 151600
rect 224572 151542 226859 151544
rect 226793 151539 226859 151542
rect 57421 150786 57487 150789
rect 57421 150784 60076 150786
rect 57421 150728 57426 150784
rect 57482 150728 60076 150784
rect 57421 150726 60076 150728
rect 57421 150723 57487 150726
rect -960 149834 480 149924
rect 3693 149834 3759 149837
rect -960 149832 3759 149834
rect -960 149776 3698 149832
rect 3754 149776 3759 149832
rect -960 149774 3759 149776
rect -960 149684 480 149774
rect 3693 149771 3759 149774
rect 226241 148882 226307 148885
rect 224572 148880 226307 148882
rect 224572 148824 226246 148880
rect 226302 148824 226307 148880
rect 224572 148822 226307 148824
rect 226241 148819 226307 148822
rect 56317 147794 56383 147797
rect 56317 147792 60076 147794
rect 56317 147736 56322 147792
rect 56378 147736 60076 147792
rect 56317 147734 60076 147736
rect 56317 147731 56383 147734
rect 226006 147732 226012 147796
rect 226076 147794 226082 147796
rect 226241 147794 226307 147797
rect 226076 147792 226307 147794
rect 226076 147736 226246 147792
rect 226302 147736 226307 147792
rect 226076 147734 226307 147736
rect 226076 147732 226082 147734
rect 226241 147731 226307 147734
rect 226425 146162 226491 146165
rect 224572 146160 226491 146162
rect 224572 146104 226430 146160
rect 226486 146104 226491 146160
rect 224572 146102 226491 146104
rect 226425 146099 226491 146102
rect 57421 144802 57487 144805
rect 57421 144800 60076 144802
rect 57421 144744 57426 144800
rect 57482 144744 60076 144800
rect 57421 144742 60076 144744
rect 57421 144739 57487 144742
rect 226149 143578 226215 143581
rect 225830 143576 226215 143578
rect 225830 143520 226154 143576
rect 226210 143520 226215 143576
rect 225830 143518 226215 143520
rect 225830 143442 225890 143518
rect 226149 143515 226215 143518
rect 226149 143444 226215 143445
rect 226149 143442 226196 143444
rect 224572 143382 225890 143442
rect 226104 143440 226196 143442
rect 226104 143384 226154 143440
rect 226104 143382 226196 143384
rect 226149 143380 226196 143382
rect 226260 143380 226266 143444
rect 226149 143379 226215 143380
rect 57789 141810 57855 141813
rect 57789 141808 60076 141810
rect 57789 141752 57794 141808
rect 57850 141752 60076 141808
rect 57789 141750 60076 141752
rect 57789 141747 57855 141750
rect 234061 140722 234127 140725
rect 224572 140720 234127 140722
rect 224572 140664 234066 140720
rect 234122 140664 234127 140720
rect 224572 140662 234127 140664
rect 234061 140659 234127 140662
rect 583520 139362 584960 139452
rect 583342 139302 584960 139362
rect 583342 139226 583402 139302
rect 583520 139226 584960 139302
rect 583342 139212 584960 139226
rect 583342 139166 583586 139212
rect 59537 138818 59603 138821
rect 59537 138816 60076 138818
rect 59537 138760 59542 138816
rect 59598 138760 60076 138816
rect 59537 138758 60076 138760
rect 59537 138755 59603 138758
rect 236637 138138 236703 138141
rect 583526 138138 583586 139166
rect 236637 138136 583586 138138
rect 236637 138080 236642 138136
rect 236698 138080 583586 138136
rect 236637 138078 583586 138080
rect 236637 138075 236703 138078
rect 226609 138002 226675 138005
rect 224572 138000 226675 138002
rect 224572 137944 226614 138000
rect 226670 137944 226675 138000
rect 224572 137942 226675 137944
rect 226609 137939 226675 137942
rect -960 136778 480 136868
rect 3325 136778 3391 136781
rect -960 136776 3391 136778
rect -960 136720 3330 136776
rect 3386 136720 3391 136776
rect -960 136718 3391 136720
rect -960 136628 480 136718
rect 3325 136715 3391 136718
rect 57605 135826 57671 135829
rect 57605 135824 60076 135826
rect 57605 135768 57610 135824
rect 57666 135768 60076 135824
rect 57605 135766 60076 135768
rect 57605 135763 57671 135766
rect 226701 135282 226767 135285
rect 224572 135280 226767 135282
rect 224572 135224 226706 135280
rect 226762 135224 226767 135280
rect 224572 135222 226767 135224
rect 226701 135219 226767 135222
rect 57789 132834 57855 132837
rect 57789 132832 60076 132834
rect 57789 132776 57794 132832
rect 57850 132776 60076 132832
rect 57789 132774 60076 132776
rect 57789 132771 57855 132774
rect 226057 132426 226123 132429
rect 224572 132424 226123 132426
rect 224572 132368 226062 132424
rect 226118 132368 226123 132424
rect 224572 132366 226123 132368
rect 226057 132363 226123 132366
rect 58157 129842 58223 129845
rect 58157 129840 60076 129842
rect 58157 129784 58162 129840
rect 58218 129784 60076 129840
rect 58157 129782 60076 129784
rect 58157 129779 58223 129782
rect 230657 129706 230723 129709
rect 224572 129704 230723 129706
rect 224572 129648 230662 129704
rect 230718 129648 230723 129704
rect 224572 129646 230723 129648
rect 230657 129643 230723 129646
rect 57605 126986 57671 126989
rect 226926 126986 226932 126988
rect 57605 126984 60076 126986
rect 57605 126928 57610 126984
rect 57666 126928 60076 126984
rect 57605 126926 60076 126928
rect 224572 126926 226932 126986
rect 57605 126923 57671 126926
rect 226926 126924 226932 126926
rect 226996 126924 227002 126988
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect 226517 125490 226583 125493
rect 235257 125490 235323 125493
rect 226517 125488 235323 125490
rect 226517 125432 226522 125488
rect 226578 125432 235262 125488
rect 235318 125432 235323 125488
rect 226517 125430 235323 125432
rect 226517 125427 226583 125430
rect 235257 125427 235323 125430
rect 226517 124266 226583 124269
rect 224572 124264 226583 124266
rect 224572 124208 226522 124264
rect 226578 124208 226583 124264
rect 224572 124206 226583 124208
rect 226517 124203 226583 124206
rect 59077 123994 59143 123997
rect 59077 123992 60076 123994
rect 59077 123936 59082 123992
rect 59138 123936 60076 123992
rect 59077 123934 60076 123936
rect 59077 123931 59143 123934
rect -960 123572 480 123812
rect 226517 122770 226583 122773
rect 238201 122770 238267 122773
rect 226517 122768 238267 122770
rect 226517 122712 226522 122768
rect 226578 122712 238206 122768
rect 238262 122712 238267 122768
rect 226517 122710 238267 122712
rect 226517 122707 226583 122710
rect 238201 122707 238267 122710
rect 226517 121546 226583 121549
rect 224572 121544 226583 121546
rect 224572 121488 226522 121544
rect 226578 121488 226583 121544
rect 224572 121486 226583 121488
rect 226517 121483 226583 121486
rect 57605 121002 57671 121005
rect 57605 121000 60076 121002
rect 57605 120944 57610 121000
rect 57666 120944 60076 121000
rect 57605 120942 60076 120944
rect 57605 120939 57671 120942
rect 230749 118826 230815 118829
rect 224572 118824 230815 118826
rect 224572 118768 230754 118824
rect 230810 118768 230815 118824
rect 224572 118766 230815 118768
rect 230749 118763 230815 118766
rect 57145 118010 57211 118013
rect 57145 118008 60076 118010
rect 57145 117952 57150 118008
rect 57206 117952 60076 118008
rect 57145 117950 60076 117952
rect 57145 117947 57211 117950
rect 226517 117194 226583 117197
rect 251265 117194 251331 117197
rect 226517 117192 251331 117194
rect 226517 117136 226522 117192
rect 226578 117136 251270 117192
rect 251326 117136 251331 117192
rect 226517 117134 251331 117136
rect 226517 117131 226583 117134
rect 251265 117131 251331 117134
rect 226517 116106 226583 116109
rect 224572 116104 226583 116106
rect 224572 116048 226522 116104
rect 226578 116048 226583 116104
rect 224572 116046 226583 116048
rect 226517 116043 226583 116046
rect 57697 115018 57763 115021
rect 57697 115016 60076 115018
rect 57697 114960 57702 115016
rect 57758 114960 60076 115016
rect 57697 114958 60076 114960
rect 57697 114955 57763 114958
rect 226742 113386 226748 113388
rect 224572 113326 226748 113386
rect 226742 113324 226748 113326
rect 226812 113324 226818 113388
rect 583520 112842 584960 112932
rect 583342 112782 584960 112842
rect 583342 112706 583402 112782
rect 583520 112706 584960 112782
rect 583342 112692 584960 112706
rect 583342 112646 583586 112692
rect 57605 112026 57671 112029
rect 57605 112024 60076 112026
rect 57605 111968 57610 112024
rect 57666 111968 60076 112024
rect 57605 111966 60076 111968
rect 57605 111963 57671 111966
rect 228214 111828 228220 111892
rect 228284 111890 228290 111892
rect 583526 111890 583586 112646
rect 228284 111830 583586 111890
rect 228284 111828 228290 111830
rect -960 110666 480 110756
rect 3141 110666 3207 110669
rect 233417 110666 233483 110669
rect -960 110664 3207 110666
rect -960 110608 3146 110664
rect 3202 110608 3207 110664
rect -960 110606 3207 110608
rect 224572 110664 233483 110666
rect 224572 110608 233422 110664
rect 233478 110608 233483 110664
rect 224572 110606 233483 110608
rect -960 110516 480 110606
rect 3141 110603 3207 110606
rect 233417 110603 233483 110606
rect 57053 109034 57119 109037
rect 57053 109032 60076 109034
rect 57053 108976 57058 109032
rect 57114 108976 60076 109032
rect 57053 108974 60076 108976
rect 57053 108971 57119 108974
rect 232313 107810 232379 107813
rect 224572 107808 232379 107810
rect 224572 107752 232318 107808
rect 232374 107752 232379 107808
rect 224572 107750 232379 107752
rect 232313 107747 232379 107750
rect 57605 106042 57671 106045
rect 57605 106040 60076 106042
rect 57605 105984 57610 106040
rect 57666 105984 60076 106040
rect 57605 105982 60076 105984
rect 57605 105979 57671 105982
rect 231117 105090 231183 105093
rect 224572 105088 231183 105090
rect 224572 105032 231122 105088
rect 231178 105032 231183 105088
rect 224572 105030 231183 105032
rect 231117 105027 231183 105030
rect 57605 103050 57671 103053
rect 57605 103048 60076 103050
rect 57605 102992 57610 103048
rect 57666 102992 60076 103048
rect 57605 102990 60076 102992
rect 57605 102987 57671 102990
rect 233325 102370 233391 102373
rect 224572 102368 233391 102370
rect 224572 102312 233330 102368
rect 233386 102312 233391 102368
rect 224572 102310 233391 102312
rect 233325 102307 233391 102310
rect 57605 100058 57671 100061
rect 57605 100056 60076 100058
rect 57605 100000 57610 100056
rect 57666 100000 60076 100056
rect 57605 99998 60076 100000
rect 57605 99995 57671 99998
rect 233233 99650 233299 99653
rect 224572 99648 233299 99650
rect 224572 99592 233238 99648
rect 233294 99592 233299 99648
rect 224572 99590 233299 99592
rect 233233 99587 233299 99590
rect 235441 99514 235507 99517
rect 583520 99514 584960 99604
rect 235441 99512 584960 99514
rect 235441 99456 235446 99512
rect 235502 99456 584960 99512
rect 235441 99454 584960 99456
rect 235441 99451 235507 99454
rect 583520 99364 584960 99454
rect 226517 97882 226583 97885
rect 246297 97882 246363 97885
rect 226517 97880 246363 97882
rect 226517 97824 226522 97880
rect 226578 97824 246302 97880
rect 246358 97824 246363 97880
rect 226517 97822 246363 97824
rect 226517 97819 226583 97822
rect 246297 97819 246363 97822
rect -960 97610 480 97700
rect 3233 97610 3299 97613
rect -960 97608 3299 97610
rect -960 97552 3238 97608
rect 3294 97552 3299 97608
rect -960 97550 3299 97552
rect -960 97460 480 97550
rect 3233 97547 3299 97550
rect 58801 97066 58867 97069
rect 58801 97064 60076 97066
rect 58801 97008 58806 97064
rect 58862 97008 60076 97064
rect 58801 97006 60076 97008
rect 58801 97003 58867 97006
rect 226517 96930 226583 96933
rect 224572 96928 226583 96930
rect 224572 96872 226522 96928
rect 226578 96872 226583 96928
rect 224572 96870 226583 96872
rect 226517 96867 226583 96870
rect 58249 94210 58315 94213
rect 233509 94210 233575 94213
rect 58249 94208 60076 94210
rect 58249 94152 58254 94208
rect 58310 94152 60076 94208
rect 58249 94150 60076 94152
rect 224572 94208 233575 94210
rect 224572 94152 233514 94208
rect 233570 94152 233575 94208
rect 224572 94150 233575 94152
rect 58249 94147 58315 94150
rect 233509 94147 233575 94150
rect 226517 92442 226583 92445
rect 249149 92442 249215 92445
rect 226517 92440 249215 92442
rect 226517 92384 226522 92440
rect 226578 92384 249154 92440
rect 249210 92384 249215 92440
rect 226517 92382 249215 92384
rect 226517 92379 226583 92382
rect 249149 92379 249215 92382
rect 226517 91490 226583 91493
rect 224572 91488 226583 91490
rect 224572 91432 226522 91488
rect 226578 91432 226583 91488
rect 224572 91430 226583 91432
rect 226517 91427 226583 91430
rect 57513 91218 57579 91221
rect 57513 91216 60076 91218
rect 57513 91160 57518 91216
rect 57574 91160 60076 91216
rect 57513 91158 60076 91160
rect 57513 91155 57579 91158
rect 229277 88770 229343 88773
rect 224572 88768 229343 88770
rect 224572 88712 229282 88768
rect 229338 88712 229343 88768
rect 224572 88710 229343 88712
rect 229277 88707 229343 88710
rect 57605 88226 57671 88229
rect 57605 88224 60076 88226
rect 57605 88168 57610 88224
rect 57666 88168 60076 88224
rect 57605 88166 60076 88168
rect 57605 88163 57671 88166
rect 226517 86866 226583 86869
rect 233877 86866 233943 86869
rect 226517 86864 233943 86866
rect 226517 86808 226522 86864
rect 226578 86808 233882 86864
rect 233938 86808 233943 86864
rect 226517 86806 233943 86808
rect 226517 86803 226583 86806
rect 233877 86803 233943 86806
rect 580349 86186 580415 86189
rect 583520 86186 584960 86276
rect 580349 86184 584960 86186
rect 580349 86128 580354 86184
rect 580410 86128 584960 86184
rect 580349 86126 584960 86128
rect 580349 86123 580415 86126
rect 226517 86050 226583 86053
rect 224572 86048 226583 86050
rect 224572 85992 226522 86048
rect 226578 85992 226583 86048
rect 583520 86036 584960 86126
rect 224572 85990 226583 85992
rect 226517 85987 226583 85990
rect 58341 85234 58407 85237
rect 58341 85232 60076 85234
rect 58341 85176 58346 85232
rect 58402 85176 60076 85232
rect 58341 85174 60076 85176
rect 58341 85171 58407 85174
rect -960 84690 480 84780
rect 3325 84690 3391 84693
rect -960 84688 3391 84690
rect -960 84632 3330 84688
rect 3386 84632 3391 84688
rect -960 84630 3391 84632
rect -960 84540 480 84630
rect 3325 84627 3391 84630
rect 232037 83194 232103 83197
rect 224572 83192 232103 83194
rect 224572 83136 232042 83192
rect 232098 83136 232103 83192
rect 224572 83134 232103 83136
rect 232037 83131 232103 83134
rect 57237 82242 57303 82245
rect 57237 82240 60076 82242
rect 57237 82184 57242 82240
rect 57298 82184 60076 82240
rect 57237 82182 60076 82184
rect 57237 82179 57303 82182
rect 232129 80474 232195 80477
rect 224572 80472 232195 80474
rect 224572 80416 232134 80472
rect 232190 80416 232195 80472
rect 224572 80414 232195 80416
rect 232129 80411 232195 80414
rect 57145 79250 57211 79253
rect 57145 79248 60076 79250
rect 57145 79192 57150 79248
rect 57206 79192 60076 79248
rect 57145 79190 60076 79192
rect 57145 79187 57211 79190
rect 228633 77754 228699 77757
rect 224572 77752 228699 77754
rect 224572 77696 228638 77752
rect 228694 77696 228699 77752
rect 224572 77694 228699 77696
rect 228633 77691 228699 77694
rect 59169 76258 59235 76261
rect 59169 76256 60076 76258
rect 59169 76200 59174 76256
rect 59230 76200 60076 76256
rect 59169 76198 60076 76200
rect 59169 76195 59235 76198
rect 226558 75034 226564 75036
rect 224572 74974 226564 75034
rect 226558 74972 226564 74974
rect 226628 74972 226634 75036
rect 56133 73266 56199 73269
rect 56133 73264 60076 73266
rect 56133 73208 56138 73264
rect 56194 73208 60076 73264
rect 56133 73206 60076 73208
rect 56133 73203 56199 73206
rect 226517 73130 226583 73133
rect 232497 73130 232563 73133
rect 226517 73128 232563 73130
rect 226517 73072 226522 73128
rect 226578 73072 232502 73128
rect 232558 73072 232563 73128
rect 226517 73070 232563 73072
rect 226517 73067 226583 73070
rect 232497 73067 232563 73070
rect 583520 72994 584960 73084
rect 583342 72934 584960 72994
rect 583342 72858 583402 72934
rect 583520 72858 584960 72934
rect 583342 72844 584960 72858
rect 583342 72798 583586 72844
rect 226517 72314 226583 72317
rect 224572 72312 226583 72314
rect 224572 72256 226522 72312
rect 226578 72256 226583 72312
rect 224572 72254 226583 72256
rect 226517 72251 226583 72254
rect 242433 71906 242499 71909
rect 583526 71906 583586 72798
rect 242433 71904 583586 71906
rect 242433 71848 242438 71904
rect 242494 71848 583586 71904
rect 242433 71846 583586 71848
rect 242433 71843 242499 71846
rect -960 71634 480 71724
rect 3325 71634 3391 71637
rect -960 71632 3391 71634
rect -960 71576 3330 71632
rect 3386 71576 3391 71632
rect -960 71574 3391 71576
rect -960 71484 480 71574
rect 3325 71571 3391 71574
rect 57605 70274 57671 70277
rect 57605 70272 60076 70274
rect 57605 70216 57610 70272
rect 57666 70216 60076 70272
rect 57605 70214 60076 70216
rect 57605 70211 57671 70214
rect 224902 70212 224908 70276
rect 224972 70274 224978 70276
rect 225454 70274 225460 70276
rect 224972 70214 225460 70274
rect 224972 70212 224978 70214
rect 225454 70212 225460 70214
rect 225524 70212 225530 70276
rect 232221 69594 232287 69597
rect 224572 69592 232287 69594
rect 224572 69536 232226 69592
rect 232282 69536 232287 69592
rect 224572 69534 232287 69536
rect 232221 69531 232287 69534
rect 59261 67282 59327 67285
rect 59261 67280 60076 67282
rect 59261 67224 59266 67280
rect 59322 67224 60076 67280
rect 59261 67222 60076 67224
rect 59261 67219 59327 67222
rect 227345 66874 227411 66877
rect 224572 66872 227411 66874
rect 224572 66816 227350 66872
rect 227406 66816 227411 66872
rect 224572 66814 227411 66816
rect 227345 66811 227411 66814
rect 225781 65650 225847 65653
rect 225646 65648 225847 65650
rect 225646 65592 225786 65648
rect 225842 65592 225847 65648
rect 225646 65590 225847 65592
rect 225646 65242 225706 65590
rect 225781 65587 225847 65590
rect 225965 65650 226031 65653
rect 225965 65648 226258 65650
rect 225965 65592 225970 65648
rect 226026 65592 226258 65648
rect 225965 65590 226258 65592
rect 225965 65587 226031 65590
rect 225873 65514 225939 65517
rect 226057 65514 226123 65517
rect 225873 65512 226123 65514
rect 225873 65456 225878 65512
rect 225934 65456 226062 65512
rect 226118 65456 226123 65512
rect 225873 65454 226123 65456
rect 225873 65451 225939 65454
rect 226057 65451 226123 65454
rect 225965 65378 226031 65381
rect 226198 65378 226258 65590
rect 225965 65376 226258 65378
rect 225965 65320 225970 65376
rect 226026 65320 226258 65376
rect 225965 65318 226258 65320
rect 225965 65315 226031 65318
rect 225781 65242 225847 65245
rect 225646 65240 225847 65242
rect 225646 65184 225786 65240
rect 225842 65184 225847 65240
rect 225646 65182 225847 65184
rect 225781 65179 225847 65182
rect 56869 64290 56935 64293
rect 56869 64288 60076 64290
rect 56869 64232 56874 64288
rect 56930 64232 60076 64288
rect 56869 64230 60076 64232
rect 56869 64227 56935 64230
rect 225229 64154 225295 64157
rect 224572 64152 225295 64154
rect 224572 64096 225234 64152
rect 225290 64096 225295 64152
rect 224572 64094 225295 64096
rect 225229 64091 225295 64094
rect 225689 62794 225755 62797
rect 225873 62794 225939 62797
rect 225689 62792 225939 62794
rect 225689 62736 225694 62792
rect 225750 62736 225878 62792
rect 225934 62736 225939 62792
rect 225689 62734 225939 62736
rect 225689 62731 225755 62734
rect 225873 62731 225939 62734
rect 227621 62114 227687 62117
rect 235349 62114 235415 62117
rect 227621 62112 235415 62114
rect 227621 62056 227626 62112
rect 227682 62056 235354 62112
rect 235410 62056 235415 62112
rect 227621 62054 235415 62056
rect 227621 62051 227687 62054
rect 235349 62051 235415 62054
rect 57329 61434 57395 61437
rect 227621 61434 227687 61437
rect 57329 61432 60076 61434
rect 57329 61376 57334 61432
rect 57390 61376 60076 61432
rect 57329 61374 60076 61376
rect 224572 61432 227687 61434
rect 224572 61376 227626 61432
rect 227682 61376 227687 61432
rect 224572 61374 227687 61376
rect 57329 61371 57395 61374
rect 227621 61371 227687 61374
rect 224902 60692 224908 60756
rect 224972 60754 224978 60756
rect 225454 60754 225460 60756
rect 224972 60694 225460 60754
rect 224972 60692 224978 60694
rect 225454 60692 225460 60694
rect 225524 60692 225530 60756
rect 225321 60482 225387 60485
rect 225689 60482 225755 60485
rect 225321 60480 225755 60482
rect 225321 60424 225326 60480
rect 225382 60424 225694 60480
rect 225750 60424 225755 60480
rect 225321 60422 225755 60424
rect 225321 60419 225387 60422
rect 225689 60419 225755 60422
rect 223614 60284 223620 60348
rect 223684 60346 223690 60348
rect 224401 60346 224467 60349
rect 223684 60344 224467 60346
rect 223684 60288 224406 60344
rect 224462 60288 224467 60344
rect 223684 60286 224467 60288
rect 223684 60284 223690 60286
rect 224401 60283 224467 60286
rect 225321 60346 225387 60349
rect 225321 60344 229110 60346
rect 225321 60288 225326 60344
rect 225382 60288 229110 60344
rect 225321 60286 229110 60288
rect 225321 60283 225387 60286
rect 222653 60210 222719 60213
rect 225086 60210 225092 60212
rect 222653 60208 225092 60210
rect 222653 60152 222658 60208
rect 222714 60152 225092 60208
rect 222653 60150 225092 60152
rect 222653 60147 222719 60150
rect 225086 60148 225092 60150
rect 225156 60148 225162 60212
rect 225229 60210 225295 60213
rect 229050 60210 229110 60286
rect 244365 60210 244431 60213
rect 225229 60208 226258 60210
rect 225229 60152 225234 60208
rect 225290 60152 226258 60208
rect 225229 60150 226258 60152
rect 229050 60208 244431 60210
rect 229050 60152 244370 60208
rect 244426 60152 244431 60208
rect 229050 60150 244431 60152
rect 225229 60147 225295 60150
rect 211889 60074 211955 60077
rect 223573 60074 223639 60077
rect 226057 60074 226123 60077
rect 211889 60072 219450 60074
rect 211889 60016 211894 60072
rect 211950 60016 219450 60072
rect 211889 60014 219450 60016
rect 211889 60011 211955 60014
rect 219390 59938 219450 60014
rect 223573 60072 226123 60074
rect 223573 60016 223578 60072
rect 223634 60016 226062 60072
rect 226118 60016 226123 60072
rect 223573 60014 226123 60016
rect 226198 60074 226258 60150
rect 244365 60147 244431 60150
rect 255313 60074 255379 60077
rect 226198 60072 255379 60074
rect 226198 60016 255318 60072
rect 255374 60016 255379 60072
rect 226198 60014 255379 60016
rect 223573 60011 223639 60014
rect 226057 60011 226123 60014
rect 255313 60011 255379 60014
rect 249885 59938 249951 59941
rect 219390 59936 249951 59938
rect 219390 59880 249890 59936
rect 249946 59880 249951 59936
rect 219390 59878 249951 59880
rect 249885 59875 249951 59878
rect 204713 59802 204779 59805
rect 224166 59802 224172 59804
rect 204713 59800 224172 59802
rect 204713 59744 204718 59800
rect 204774 59744 224172 59800
rect 204713 59742 224172 59744
rect 204713 59739 204779 59742
rect 224166 59740 224172 59742
rect 224236 59740 224242 59804
rect 224401 59802 224467 59805
rect 229369 59802 229435 59805
rect 224401 59800 229435 59802
rect 224401 59744 224406 59800
rect 224462 59744 229374 59800
rect 229430 59744 229435 59800
rect 224401 59742 229435 59744
rect 224401 59739 224467 59742
rect 229369 59739 229435 59742
rect 209037 59666 209103 59669
rect 242157 59666 242223 59669
rect 209037 59664 242223 59666
rect 209037 59608 209042 59664
rect 209098 59608 242162 59664
rect 242218 59608 242223 59664
rect 209037 59606 242223 59608
rect 209037 59603 209103 59606
rect 242157 59603 242223 59606
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 222745 59530 222811 59533
rect 269757 59530 269823 59533
rect 222745 59528 269823 59530
rect 222745 59472 222750 59528
rect 222806 59472 269762 59528
rect 269818 59472 269823 59528
rect 583520 59516 584960 59606
rect 222745 59470 269823 59472
rect 222745 59467 222811 59470
rect 269757 59467 269823 59470
rect 221641 59394 221707 59397
rect 269113 59394 269179 59397
rect 221641 59392 269179 59394
rect 221641 59336 221646 59392
rect 221702 59336 269118 59392
rect 269174 59336 269179 59392
rect 221641 59334 269179 59336
rect 221641 59331 221707 59334
rect 269113 59331 269179 59334
rect 218145 59258 218211 59261
rect 220169 59258 220235 59261
rect 227662 59258 227668 59260
rect 218145 59256 220002 59258
rect 218145 59200 218150 59256
rect 218206 59200 220002 59256
rect 218145 59198 220002 59200
rect 218145 59195 218211 59198
rect 219249 59122 219315 59125
rect 219249 59120 219818 59122
rect 219249 59064 219254 59120
rect 219310 59064 219818 59120
rect 219249 59062 219818 59064
rect 219249 59059 219315 59062
rect 218697 58986 218763 58989
rect 219617 58986 219683 58989
rect 218697 58984 219683 58986
rect 218697 58928 218702 58984
rect 218758 58928 219622 58984
rect 219678 58928 219683 58984
rect 218697 58926 219683 58928
rect 218697 58923 218763 58926
rect 219617 58923 219683 58926
rect 219758 58850 219818 59062
rect 219942 58986 220002 59198
rect 220169 59256 227668 59258
rect 220169 59200 220174 59256
rect 220230 59200 227668 59256
rect 220169 59198 227668 59200
rect 220169 59195 220235 59198
rect 227662 59196 227668 59198
rect 227732 59196 227738 59260
rect 223573 59122 223639 59125
rect 223941 59124 224007 59125
rect 224309 59124 224375 59125
rect 223798 59122 223804 59124
rect 223573 59120 223804 59122
rect 223573 59064 223578 59120
rect 223634 59064 223804 59120
rect 223573 59062 223804 59064
rect 223573 59059 223639 59062
rect 223798 59060 223804 59062
rect 223868 59060 223874 59124
rect 223941 59120 223988 59124
rect 224052 59122 224058 59124
rect 224309 59122 224356 59124
rect 223941 59064 223946 59120
rect 223941 59060 223988 59064
rect 224052 59062 224098 59122
rect 224264 59120 224356 59122
rect 224264 59064 224314 59120
rect 224264 59062 224356 59064
rect 224052 59060 224058 59062
rect 224309 59060 224356 59062
rect 224420 59060 224426 59124
rect 223941 59059 224007 59060
rect 224309 59059 224375 59060
rect 227805 58986 227871 58989
rect 219942 58984 227871 58986
rect 219942 58928 227810 58984
rect 227866 58928 227871 58984
rect 219942 58926 227871 58928
rect 227805 58923 227871 58926
rect 227846 58850 227852 58852
rect 219758 58790 227852 58850
rect 227846 58788 227852 58790
rect 227916 58788 227922 58852
rect 206185 58714 206251 58717
rect 356513 58714 356579 58717
rect 206185 58712 356579 58714
rect -960 58578 480 58668
rect 206185 58656 206190 58712
rect 206246 58656 356518 58712
rect 356574 58656 356579 58712
rect 206185 58654 356579 58656
rect 206185 58651 206251 58654
rect 356513 58651 356579 58654
rect 3509 58578 3575 58581
rect -960 58576 3575 58578
rect -960 58520 3514 58576
rect 3570 58520 3575 58576
rect -960 58518 3575 58520
rect -960 58428 480 58518
rect 3509 58515 3575 58518
rect 214649 58578 214715 58581
rect 219617 58578 219683 58581
rect 227713 58578 227779 58581
rect 214649 58576 219450 58578
rect 214649 58520 214654 58576
rect 214710 58520 219450 58576
rect 214649 58518 219450 58520
rect 214649 58515 214715 58518
rect 219390 58442 219450 58518
rect 219617 58576 227779 58578
rect 219617 58520 219622 58576
rect 219678 58520 227718 58576
rect 227774 58520 227779 58576
rect 219617 58518 227779 58520
rect 219617 58515 219683 58518
rect 227713 58515 227779 58518
rect 226374 58442 226380 58444
rect 219390 58382 226380 58442
rect 226374 58380 226380 58382
rect 226444 58380 226450 58444
rect 221825 58306 221891 58309
rect 224401 58306 224467 58309
rect 221825 58304 224467 58306
rect 221825 58248 221830 58304
rect 221886 58248 224406 58304
rect 224462 58248 224467 58304
rect 221825 58246 224467 58248
rect 221825 58243 221891 58246
rect 224401 58243 224467 58246
rect 58893 57898 58959 57901
rect 210509 57898 210575 57901
rect 58893 57896 210575 57898
rect 58893 57840 58898 57896
rect 58954 57840 210514 57896
rect 210570 57840 210575 57896
rect 58893 57838 210575 57840
rect 58893 57835 58959 57838
rect 210509 57835 210575 57838
rect 211429 57898 211495 57901
rect 220445 57898 220511 57901
rect 224902 57898 224908 57900
rect 211429 57896 219450 57898
rect 211429 57840 211434 57896
rect 211490 57840 219450 57896
rect 211429 57838 219450 57840
rect 211429 57835 211495 57838
rect 56501 57762 56567 57765
rect 62113 57762 62179 57765
rect 207013 57762 207079 57765
rect 56501 57760 62179 57762
rect 56501 57704 56506 57760
rect 56562 57704 62118 57760
rect 62174 57704 62179 57760
rect 56501 57702 62179 57704
rect 56501 57699 56567 57702
rect 62113 57699 62179 57702
rect 70350 57760 207079 57762
rect 70350 57704 207018 57760
rect 207074 57704 207079 57760
rect 70350 57702 207079 57704
rect 12341 57626 12407 57629
rect 62665 57626 62731 57629
rect 12341 57624 62731 57626
rect 12341 57568 12346 57624
rect 12402 57568 62670 57624
rect 62726 57568 62731 57624
rect 12341 57566 62731 57568
rect 12341 57563 12407 57566
rect 62665 57563 62731 57566
rect 10961 57490 11027 57493
rect 59997 57490 60063 57493
rect 62941 57490 63007 57493
rect 10961 57488 58818 57490
rect 10961 57432 10966 57488
rect 11022 57432 58818 57488
rect 10961 57430 58818 57432
rect 10961 57427 11027 57430
rect 9581 57354 9647 57357
rect 56501 57354 56567 57357
rect 9581 57352 56567 57354
rect 9581 57296 9586 57352
rect 9642 57296 56506 57352
rect 56562 57296 56567 57352
rect 9581 57294 56567 57296
rect 58758 57354 58818 57430
rect 59997 57488 63007 57490
rect 59997 57432 60002 57488
rect 60058 57432 62946 57488
rect 63002 57432 63007 57488
rect 59997 57430 63007 57432
rect 59997 57427 60063 57430
rect 62941 57427 63007 57430
rect 62389 57354 62455 57357
rect 58758 57352 62455 57354
rect 58758 57296 62394 57352
rect 62450 57296 62455 57352
rect 58758 57294 62455 57296
rect 9581 57291 9647 57294
rect 56501 57291 56567 57294
rect 62389 57291 62455 57294
rect 4061 57218 4127 57221
rect 60917 57218 60983 57221
rect 4061 57216 60983 57218
rect 4061 57160 4066 57216
rect 4122 57160 60922 57216
rect 60978 57160 60983 57216
rect 4061 57158 60983 57160
rect 4061 57155 4127 57158
rect 60917 57155 60983 57158
rect 61837 57218 61903 57221
rect 66897 57218 66963 57221
rect 61837 57216 66963 57218
rect 61837 57160 61842 57216
rect 61898 57160 66902 57216
rect 66958 57160 66963 57216
rect 61837 57158 66963 57160
rect 61837 57155 61903 57158
rect 66897 57155 66963 57158
rect 15101 57082 15167 57085
rect 58617 57082 58683 57085
rect 70350 57082 70410 57702
rect 207013 57699 207079 57702
rect 209957 57762 210023 57765
rect 219249 57762 219315 57765
rect 209957 57760 219315 57762
rect 209957 57704 209962 57760
rect 210018 57704 219254 57760
rect 219310 57704 219315 57760
rect 209957 57702 219315 57704
rect 219390 57762 219450 57838
rect 220445 57896 224908 57898
rect 220445 57840 220450 57896
rect 220506 57840 224908 57896
rect 220445 57838 224908 57840
rect 220445 57835 220511 57838
rect 224902 57836 224908 57838
rect 224972 57836 224978 57900
rect 223481 57762 223547 57765
rect 219390 57760 223547 57762
rect 219390 57704 223486 57760
rect 223542 57704 223547 57760
rect 219390 57702 223547 57704
rect 209957 57699 210023 57702
rect 219249 57699 219315 57702
rect 223481 57699 223547 57702
rect 143901 57626 143967 57629
rect 137326 57624 143967 57626
rect 137326 57568 143906 57624
rect 143962 57568 143967 57624
rect 137326 57566 143967 57568
rect 103053 57490 103119 57493
rect 103513 57490 103579 57493
rect 103053 57488 103579 57490
rect 103053 57432 103058 57488
rect 103114 57432 103518 57488
rect 103574 57432 103579 57488
rect 103053 57430 103579 57432
rect 103053 57427 103119 57430
rect 103513 57427 103579 57430
rect 131941 57490 132007 57493
rect 132861 57490 132927 57493
rect 131941 57488 132927 57490
rect 131941 57432 131946 57488
rect 132002 57432 132866 57488
rect 132922 57432 132927 57488
rect 131941 57430 132927 57432
rect 131941 57427 132007 57430
rect 132861 57427 132927 57430
rect 120993 57354 121059 57357
rect 137326 57354 137386 57566
rect 143901 57563 143967 57566
rect 171041 57626 171107 57629
rect 171593 57626 171659 57629
rect 171041 57624 171659 57626
rect 171041 57568 171046 57624
rect 171102 57568 171598 57624
rect 171654 57568 171659 57624
rect 171041 57566 171659 57568
rect 171041 57563 171107 57566
rect 171593 57563 171659 57566
rect 206737 57626 206803 57629
rect 225597 57626 225663 57629
rect 206737 57624 225663 57626
rect 206737 57568 206742 57624
rect 206798 57568 225602 57624
rect 225658 57568 225663 57624
rect 206737 57566 225663 57568
rect 206737 57563 206803 57566
rect 225597 57563 225663 57566
rect 140405 57490 140471 57493
rect 160461 57490 160527 57493
rect 140405 57488 160527 57490
rect 140405 57432 140410 57488
rect 140466 57432 160466 57488
rect 160522 57432 160527 57488
rect 140405 57430 160527 57432
rect 140405 57427 140471 57430
rect 160461 57427 160527 57430
rect 209681 57490 209747 57493
rect 225137 57490 225203 57493
rect 209681 57488 225203 57490
rect 209681 57432 209686 57488
rect 209742 57432 225142 57488
rect 225198 57432 225203 57488
rect 209681 57430 225203 57432
rect 209681 57427 209747 57430
rect 225137 57427 225203 57430
rect 120993 57352 137386 57354
rect 120993 57296 120998 57352
rect 121054 57296 137386 57352
rect 120993 57294 137386 57296
rect 146293 57354 146359 57357
rect 347037 57354 347103 57357
rect 146293 57352 347103 57354
rect 146293 57296 146298 57352
rect 146354 57296 347042 57352
rect 347098 57296 347103 57352
rect 146293 57294 347103 57296
rect 120993 57291 121059 57294
rect 146293 57291 146359 57294
rect 347037 57291 347103 57294
rect 118325 57218 118391 57221
rect 142061 57218 142127 57221
rect 142245 57218 142311 57221
rect 118325 57216 137386 57218
rect 118325 57160 118330 57216
rect 118386 57160 137386 57216
rect 118325 57158 137386 57160
rect 118325 57155 118391 57158
rect 15101 57080 58450 57082
rect 15101 57024 15106 57080
rect 15162 57024 58450 57080
rect 15101 57022 58450 57024
rect 15101 57019 15167 57022
rect 13721 56946 13787 56949
rect 58390 56946 58450 57022
rect 58617 57080 70410 57082
rect 58617 57024 58622 57080
rect 58678 57024 70410 57080
rect 58617 57022 70410 57024
rect 116853 57082 116919 57085
rect 118969 57082 119035 57085
rect 116853 57080 119035 57082
rect 116853 57024 116858 57080
rect 116914 57024 118974 57080
rect 119030 57024 119035 57080
rect 116853 57022 119035 57024
rect 58617 57019 58683 57022
rect 116853 57019 116919 57022
rect 118969 57019 119035 57022
rect 129181 57082 129247 57085
rect 133045 57082 133111 57085
rect 134793 57082 134859 57085
rect 129181 57080 132970 57082
rect 129181 57024 129186 57080
rect 129242 57024 132970 57080
rect 129181 57022 132970 57024
rect 129181 57019 129247 57022
rect 63585 56946 63651 56949
rect 13721 56944 58266 56946
rect 13721 56888 13726 56944
rect 13782 56888 58266 56944
rect 13721 56886 58266 56888
rect 58390 56944 63651 56946
rect 58390 56888 63590 56944
rect 63646 56888 63651 56944
rect 58390 56886 63651 56888
rect 13721 56883 13787 56886
rect 17861 56810 17927 56813
rect 58206 56810 58266 56886
rect 63585 56883 63651 56886
rect 63769 56946 63835 56949
rect 65517 56946 65583 56949
rect 63769 56944 65583 56946
rect 63769 56888 63774 56944
rect 63830 56888 65522 56944
rect 65578 56888 65583 56944
rect 63769 56886 65583 56888
rect 63769 56883 63835 56886
rect 65517 56883 65583 56886
rect 118601 56946 118667 56949
rect 126329 56946 126395 56949
rect 118601 56944 126395 56946
rect 118601 56888 118606 56944
rect 118662 56888 126334 56944
rect 126390 56888 126395 56944
rect 118601 56886 126395 56888
rect 118601 56883 118667 56886
rect 126329 56883 126395 56886
rect 129917 56946 129983 56949
rect 132493 56946 132559 56949
rect 129917 56944 132559 56946
rect 129917 56888 129922 56944
rect 129978 56888 132498 56944
rect 132554 56888 132559 56944
rect 129917 56886 132559 56888
rect 129917 56883 129983 56886
rect 132493 56883 132559 56886
rect 132677 56946 132743 56949
rect 132910 56946 132970 57022
rect 133045 57080 134859 57082
rect 133045 57024 133050 57080
rect 133106 57024 134798 57080
rect 134854 57024 134859 57080
rect 133045 57022 134859 57024
rect 137326 57082 137386 57158
rect 142061 57216 142311 57218
rect 142061 57160 142066 57216
rect 142122 57160 142250 57216
rect 142306 57160 142311 57216
rect 142061 57158 142311 57160
rect 142061 57155 142127 57158
rect 142245 57155 142311 57158
rect 203517 57218 203583 57221
rect 429837 57218 429903 57221
rect 203517 57216 429903 57218
rect 203517 57160 203522 57216
rect 203578 57160 429842 57216
rect 429898 57160 429903 57216
rect 203517 57158 429903 57160
rect 203517 57155 203583 57158
rect 429837 57155 429903 57158
rect 142889 57082 142955 57085
rect 137326 57080 142955 57082
rect 137326 57024 142894 57080
rect 142950 57024 142955 57080
rect 137326 57022 142955 57024
rect 133045 57019 133111 57022
rect 134793 57019 134859 57022
rect 142889 57019 142955 57022
rect 166349 57082 166415 57085
rect 168649 57082 168715 57085
rect 166349 57080 168715 57082
rect 166349 57024 166354 57080
rect 166410 57024 168654 57080
rect 168710 57024 168715 57080
rect 166349 57022 168715 57024
rect 166349 57019 166415 57022
rect 168649 57019 168715 57022
rect 218973 57082 219039 57085
rect 224902 57082 224908 57084
rect 218973 57080 224908 57082
rect 218973 57024 218978 57080
rect 219034 57024 224908 57080
rect 218973 57022 224908 57024
rect 218973 57019 219039 57022
rect 224902 57020 224908 57022
rect 224972 57020 224978 57084
rect 137921 56946 137987 56949
rect 132677 56944 132786 56946
rect 132677 56888 132682 56944
rect 132738 56888 132786 56944
rect 132677 56883 132786 56888
rect 132910 56944 137987 56946
rect 132910 56888 137926 56944
rect 137982 56888 137987 56944
rect 132910 56886 137987 56888
rect 137921 56883 137987 56886
rect 208761 56946 208827 56949
rect 258073 56946 258139 56949
rect 208761 56944 258139 56946
rect 208761 56888 208766 56944
rect 208822 56888 258078 56944
rect 258134 56888 258139 56944
rect 208761 56886 258139 56888
rect 208761 56883 208827 56886
rect 258073 56883 258139 56886
rect 63217 56810 63283 56813
rect 17861 56808 45570 56810
rect 17861 56752 17866 56808
rect 17922 56752 45570 56808
rect 17861 56750 45570 56752
rect 58206 56808 63283 56810
rect 58206 56752 63222 56808
rect 63278 56752 63283 56808
rect 58206 56750 63283 56752
rect 17861 56747 17927 56750
rect 45510 56674 45570 56750
rect 63217 56747 63283 56750
rect 63401 56810 63467 56813
rect 65609 56810 65675 56813
rect 63401 56808 65675 56810
rect 63401 56752 63406 56808
rect 63462 56752 65614 56808
rect 65670 56752 65675 56808
rect 63401 56750 65675 56752
rect 63401 56747 63467 56750
rect 65609 56747 65675 56750
rect 118601 56810 118667 56813
rect 118785 56810 118851 56813
rect 118601 56808 118851 56810
rect 118601 56752 118606 56808
rect 118662 56752 118790 56808
rect 118846 56752 118851 56808
rect 118601 56750 118851 56752
rect 132726 56810 132786 56883
rect 136817 56810 136883 56813
rect 132726 56808 136883 56810
rect 132726 56752 136822 56808
rect 136878 56752 136883 56808
rect 132726 56750 136883 56752
rect 118601 56747 118667 56750
rect 118785 56747 118851 56750
rect 136817 56747 136883 56750
rect 180701 56810 180767 56813
rect 204437 56810 204503 56813
rect 244917 56810 244983 56813
rect 180701 56808 180810 56810
rect 180701 56752 180706 56808
rect 180762 56752 180810 56808
rect 180701 56747 180810 56752
rect 204437 56808 244983 56810
rect 204437 56752 204442 56808
rect 204498 56752 244922 56808
rect 244978 56752 244983 56808
rect 204437 56750 244983 56752
rect 204437 56747 204503 56750
rect 244917 56747 244983 56750
rect 180750 56677 180810 56747
rect 64137 56674 64203 56677
rect 45510 56672 64203 56674
rect 45510 56616 64142 56672
rect 64198 56616 64203 56672
rect 45510 56614 64203 56616
rect 64137 56611 64203 56614
rect 117497 56674 117563 56677
rect 123477 56674 123543 56677
rect 117497 56672 123543 56674
rect 117497 56616 117502 56672
rect 117558 56616 123482 56672
rect 123538 56616 123543 56672
rect 117497 56614 123543 56616
rect 180750 56672 180859 56677
rect 180750 56616 180798 56672
rect 180854 56616 180859 56672
rect 180750 56614 180859 56616
rect 117497 56611 117563 56614
rect 123477 56611 123543 56614
rect 180793 56611 180859 56614
rect 211153 56674 211219 56677
rect 225413 56674 225479 56677
rect 211153 56672 225479 56674
rect 211153 56616 211158 56672
rect 211214 56616 225418 56672
rect 225474 56616 225479 56672
rect 211153 56614 225479 56616
rect 211153 56611 211219 56614
rect 225413 56611 225479 56614
rect 579981 46338 580047 46341
rect 583520 46338 584960 46428
rect 579981 46336 584960 46338
rect 579981 46280 579986 46336
rect 580042 46280 584960 46336
rect 579981 46278 584960 46280
rect 579981 46275 580047 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3417 45522 3483 45525
rect -960 45520 3483 45522
rect -960 45464 3422 45520
rect 3478 45464 3483 45520
rect -960 45462 3483 45464
rect -960 45372 480 45462
rect 3417 45459 3483 45462
rect 580257 33146 580323 33149
rect 583520 33146 584960 33236
rect 580257 33144 584960 33146
rect 580257 33088 580262 33144
rect 580318 33088 584960 33144
rect 580257 33086 584960 33088
rect 580257 33083 580323 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2865 32466 2931 32469
rect -960 32464 2931 32466
rect -960 32408 2870 32464
rect 2926 32408 2931 32464
rect -960 32406 2931 32408
rect -960 32316 480 32406
rect 2865 32403 2931 32406
rect 580073 19818 580139 19821
rect 583520 19818 584960 19908
rect 580073 19816 584960 19818
rect 580073 19760 580078 19816
rect 580134 19760 584960 19816
rect 580073 19758 584960 19760
rect 580073 19755 580139 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 158621 6898 158687 6901
rect 397729 6898 397795 6901
rect 158621 6896 397795 6898
rect 158621 6840 158626 6896
rect 158682 6840 397734 6896
rect 397790 6840 397795 6896
rect 158621 6838 397795 6840
rect 158621 6835 158687 6838
rect 397729 6835 397795 6838
rect 165245 6762 165311 6765
rect 426157 6762 426223 6765
rect 165245 6760 426223 6762
rect 165245 6704 165250 6760
rect 165306 6704 426162 6760
rect 426218 6704 426223 6760
rect 165245 6702 426223 6704
rect 165245 6699 165311 6702
rect 426157 6699 426223 6702
rect 210417 6626 210483 6629
rect 472249 6626 472315 6629
rect 210417 6624 472315 6626
rect -960 6490 480 6580
rect 210417 6568 210422 6624
rect 210478 6568 472254 6624
rect 472310 6568 472315 6624
rect 210417 6566 472315 6568
rect 210417 6563 210483 6566
rect 472249 6563 472315 6566
rect 580349 6626 580415 6629
rect 583520 6626 584960 6716
rect 580349 6624 584960 6626
rect 580349 6568 580354 6624
rect 580410 6568 584960 6624
rect 580349 6566 584960 6568
rect 580349 6563 580415 6566
rect 3417 6490 3483 6493
rect -960 6488 3483 6490
rect -960 6432 3422 6488
rect 3478 6432 3483 6488
rect -960 6430 3483 6432
rect -960 6340 480 6430
rect 3417 6427 3483 6430
rect 166625 6490 166691 6493
rect 433241 6490 433307 6493
rect 166625 6488 433307 6490
rect 166625 6432 166630 6488
rect 166686 6432 433246 6488
rect 433302 6432 433307 6488
rect 583520 6476 584960 6566
rect 166625 6430 433307 6432
rect 166625 6427 166691 6430
rect 433241 6427 433307 6430
rect 168005 6354 168071 6357
rect 436645 6354 436711 6357
rect 168005 6352 436711 6354
rect 168005 6296 168010 6352
rect 168066 6296 436650 6352
rect 436706 6296 436711 6352
rect 168005 6294 436711 6296
rect 168005 6291 168071 6294
rect 436645 6291 436711 6294
rect 204069 6218 204135 6221
rect 582189 6218 582255 6221
rect 204069 6216 582255 6218
rect 204069 6160 204074 6216
rect 204130 6160 582194 6216
rect 582250 6160 582255 6216
rect 204069 6158 582255 6160
rect 204069 6155 204135 6158
rect 582189 6155 582255 6158
rect 157241 6082 157307 6085
rect 394233 6082 394299 6085
rect 157241 6080 394299 6082
rect 157241 6024 157246 6080
rect 157302 6024 394238 6080
rect 394294 6024 394299 6080
rect 157241 6022 394299 6024
rect 157241 6019 157307 6022
rect 394233 6019 394299 6022
rect 155861 5946 155927 5949
rect 383561 5946 383627 5949
rect 155861 5944 383627 5946
rect 155861 5888 155866 5944
rect 155922 5888 383566 5944
rect 383622 5888 383627 5944
rect 155861 5886 383627 5888
rect 155861 5883 155927 5886
rect 383561 5883 383627 5886
rect 151721 5810 151787 5813
rect 368473 5810 368539 5813
rect 151721 5808 368539 5810
rect 151721 5752 151726 5808
rect 151782 5752 368478 5808
rect 368534 5752 368539 5808
rect 151721 5750 368539 5752
rect 151721 5747 151787 5750
rect 368473 5747 368539 5750
rect 199653 5130 199719 5133
rect 565629 5130 565695 5133
rect 199653 5128 565695 5130
rect 199653 5072 199658 5128
rect 199714 5072 565634 5128
rect 565690 5072 565695 5128
rect 199653 5070 565695 5072
rect 199653 5067 199719 5070
rect 565629 5067 565695 5070
rect 201401 4994 201467 4997
rect 572805 4994 572871 4997
rect 201401 4992 572871 4994
rect 201401 4936 201406 4992
rect 201462 4936 572810 4992
rect 572866 4936 572871 4992
rect 201401 4934 572871 4936
rect 201401 4931 201467 4934
rect 572805 4931 572871 4934
rect 202781 4858 202847 4861
rect 576301 4858 576367 4861
rect 202781 4856 576367 4858
rect 202781 4800 202786 4856
rect 202842 4800 576306 4856
rect 576362 4800 576367 4856
rect 202781 4798 576367 4800
rect 202781 4795 202847 4798
rect 576301 4795 576367 4798
rect 213177 4042 213243 4045
rect 429653 4042 429719 4045
rect 213177 4040 429719 4042
rect 213177 3984 213182 4040
rect 213238 3984 429658 4040
rect 429714 3984 429719 4040
rect 213177 3982 429719 3984
rect 213177 3979 213243 3982
rect 429653 3979 429719 3982
rect 161105 3906 161171 3909
rect 408401 3906 408467 3909
rect 161105 3904 408467 3906
rect 161105 3848 161110 3904
rect 161166 3848 408406 3904
rect 408462 3848 408467 3904
rect 161105 3846 408467 3848
rect 161105 3843 161171 3846
rect 408401 3843 408467 3846
rect 162577 3770 162643 3773
rect 415485 3770 415551 3773
rect 162577 3768 415551 3770
rect 162577 3712 162582 3768
rect 162638 3712 415490 3768
rect 415546 3712 415551 3768
rect 162577 3710 415551 3712
rect 162577 3707 162643 3710
rect 415485 3707 415551 3710
rect 55673 3634 55739 3637
rect 59721 3634 59787 3637
rect 55673 3632 59787 3634
rect 55673 3576 55678 3632
rect 55734 3576 59726 3632
rect 59782 3576 59787 3632
rect 55673 3574 59787 3576
rect 55673 3571 55739 3574
rect 59721 3571 59787 3574
rect 163865 3634 163931 3637
rect 422569 3634 422635 3637
rect 163865 3632 422635 3634
rect 163865 3576 163870 3632
rect 163926 3576 422574 3632
rect 422630 3576 422635 3632
rect 163865 3574 422635 3576
rect 163865 3571 163931 3574
rect 422569 3571 422635 3574
rect 169661 3498 169727 3501
rect 443821 3498 443887 3501
rect 169661 3496 443887 3498
rect 169661 3440 169666 3496
rect 169722 3440 443826 3496
rect 443882 3440 443887 3496
rect 169661 3438 443887 3440
rect 169661 3435 169727 3438
rect 443821 3435 443887 3438
rect 565 3362 631 3365
rect 59353 3362 59419 3365
rect 565 3360 59419 3362
rect 565 3304 570 3360
rect 626 3304 59358 3360
rect 59414 3304 59419 3360
rect 565 3302 59419 3304
rect 565 3299 631 3302
rect 59353 3299 59419 3302
rect 175181 3362 175247 3365
rect 465165 3362 465231 3365
rect 175181 3360 465231 3362
rect 175181 3304 175186 3360
rect 175242 3304 465170 3360
rect 465226 3304 465231 3360
rect 175181 3302 465231 3304
rect 175181 3299 175247 3302
rect 465165 3299 465231 3302
rect 213545 3226 213611 3229
rect 418981 3226 419047 3229
rect 213545 3224 419047 3226
rect 213545 3168 213550 3224
rect 213606 3168 418986 3224
rect 419042 3168 419047 3224
rect 213545 3166 419047 3168
rect 213545 3163 213611 3166
rect 418981 3163 419047 3166
rect 213453 3090 213519 3093
rect 411897 3090 411963 3093
rect 213453 3088 411963 3090
rect 213453 3032 213458 3088
rect 213514 3032 411902 3088
rect 411958 3032 411963 3088
rect 213453 3030 411963 3032
rect 213453 3027 213519 3030
rect 411897 3027 411963 3030
<< via3 >>
rect 218652 491404 218716 491468
rect 218836 491268 218900 491332
rect 219204 490180 219268 490244
rect 145604 487460 145668 487524
rect 271092 487460 271156 487524
rect 111196 487188 111260 487252
rect 90956 487052 91020 487116
rect 217548 487052 217612 487116
rect 138612 486916 138676 486980
rect 326660 486916 326724 486980
rect 150940 486780 151004 486844
rect 248644 486780 248708 486844
rect 266124 486840 266188 486844
rect 266124 486784 266138 486840
rect 266138 486784 266188 486840
rect 266124 486780 266188 486784
rect 126100 486644 126164 486708
rect 130884 486704 130948 486708
rect 130884 486648 130898 486704
rect 130898 486648 130948 486704
rect 130884 486644 130948 486648
rect 143580 486644 143644 486708
rect 283788 486644 283852 486708
rect 101076 486508 101140 486572
rect 103836 486508 103900 486572
rect 108620 486508 108684 486572
rect 123708 486508 123772 486572
rect 288572 486508 288636 486572
rect 116164 486372 116228 486436
rect 305868 486372 305932 486436
rect 339724 486372 339788 486436
rect 350764 486372 350828 486436
rect 118556 486236 118620 486300
rect 313596 486236 313660 486300
rect 106228 486100 106292 486164
rect 318380 486100 318444 486164
rect 93348 485964 93412 486028
rect 98500 485964 98564 486028
rect 114324 485964 114388 486028
rect 323348 485964 323412 486028
rect 88748 485828 88812 485892
rect 158484 485828 158548 485892
rect 253428 485828 253492 485892
rect 256188 485888 256252 485892
rect 256188 485832 256202 485888
rect 256202 485832 256252 485888
rect 256188 485828 256252 485832
rect 263548 485888 263612 485892
rect 263548 485832 263598 485888
rect 263598 485832 263612 485888
rect 263548 485828 263612 485832
rect 276244 485888 276308 485892
rect 276244 485832 276258 485888
rect 276258 485832 276308 485888
rect 276244 485828 276308 485832
rect 303476 485888 303540 485892
rect 303476 485832 303490 485888
rect 303490 485832 303540 485888
rect 303476 485828 303540 485832
rect 338436 485828 338500 485892
rect 166028 485692 166092 485756
rect 178356 485616 178420 485620
rect 178356 485560 178370 485616
rect 178370 485560 178420 485616
rect 178356 485556 178420 485560
rect 260972 485556 261036 485620
rect 219020 485420 219084 485484
rect 136036 485284 136100 485348
rect 128492 485148 128556 485212
rect 251036 485148 251100 485212
rect 308260 485148 308324 485212
rect 120948 485012 121012 485076
rect 219940 485012 220004 485076
rect 295932 485012 295996 485076
rect 301084 485072 301148 485076
rect 301084 485016 301098 485072
rect 301098 485016 301148 485072
rect 301084 485012 301148 485016
rect 268516 484876 268580 484940
rect 278452 484740 278516 484804
rect 311020 484604 311084 484668
rect 179644 484468 179708 484532
rect 190868 484468 190932 484532
rect 298508 484468 298572 484532
rect 155908 484196 155972 484260
rect 219572 484256 219636 484260
rect 219572 484200 219622 484256
rect 219622 484200 219636 484256
rect 219572 484196 219636 484200
rect 161060 484060 161124 484124
rect 273484 484060 273548 484124
rect 163268 483924 163332 483988
rect 258396 483924 258460 483988
rect 133644 483788 133708 483852
rect 280934 483788 280998 483852
rect 316172 483788 316236 483852
rect 96182 483380 96246 483444
rect 141062 483380 141126 483444
rect 153574 483652 153638 483716
rect 286102 483652 286166 483716
rect 148406 483516 148470 483580
rect 290998 483516 291062 483580
rect 219756 483380 219820 483444
rect 293582 483380 293646 483444
rect 321054 483380 321118 483444
rect 218100 480252 218164 480316
rect 219388 480252 219452 480316
rect 218468 479844 218532 479908
rect 219204 479844 219268 479908
rect 218468 470732 218532 470796
rect 219204 470732 219268 470796
rect 218468 470460 218532 470524
rect 219388 470460 219452 470524
rect 218468 460940 218532 461004
rect 219388 460940 219452 461004
rect 218468 460804 218532 460868
rect 219388 460804 219452 460868
rect 218468 451284 218532 451348
rect 219388 451284 219452 451348
rect 218468 451148 218532 451212
rect 219388 451148 219452 451212
rect 218468 441628 218532 441692
rect 219388 441628 219452 441692
rect 218468 441492 218532 441556
rect 219388 441492 219452 441556
rect 218468 431972 218532 432036
rect 219388 431972 219452 432036
rect 218468 431836 218532 431900
rect 219388 431836 219452 431900
rect 218468 422316 218532 422380
rect 219388 422316 219452 422380
rect 218468 422180 218532 422244
rect 219388 422180 219452 422244
rect 218468 412660 218532 412724
rect 219388 412660 219452 412724
rect 218468 412524 218532 412588
rect 219388 412524 219452 412588
rect 219572 403276 219636 403340
rect 219572 403140 219636 403204
rect 218468 403004 218532 403068
rect 219388 403004 219452 403068
rect 218468 402868 218532 402932
rect 219388 402868 219452 402932
rect 219572 399876 219636 399940
rect 96046 399604 96110 399668
rect 96476 399604 96540 399668
rect 223620 399468 223684 399532
rect 218468 398244 218532 398308
rect 85436 398168 85500 398172
rect 85436 398112 85450 398168
rect 85450 398112 85500 398168
rect 85436 398108 85500 398112
rect 113588 398168 113652 398172
rect 113588 398112 113638 398168
rect 113638 398112 113652 398168
rect 113588 398108 113652 398112
rect 226380 398244 226444 398308
rect 219940 398108 220004 398172
rect 227852 398108 227916 398172
rect 235948 398168 236012 398172
rect 235948 398112 235998 398168
rect 235998 398112 236012 398168
rect 235948 398108 236012 398112
rect 265204 398168 265268 398172
rect 265204 398112 265218 398168
rect 265218 398112 265268 398168
rect 265204 398108 265268 398112
rect 300900 398168 300964 398172
rect 300900 398112 300914 398168
rect 300914 398112 300964 398168
rect 300900 398108 300964 398112
rect 315804 398168 315868 398172
rect 315804 398112 315818 398168
rect 315818 398112 315868 398168
rect 315804 398108 315868 398112
rect 325924 398108 325988 398172
rect 219756 397972 219820 398036
rect 227668 397836 227732 397900
rect 78260 397352 78324 397356
rect 78260 397296 78310 397352
rect 78310 397296 78324 397352
rect 78260 397292 78324 397296
rect 79548 397292 79612 397356
rect 80468 397352 80532 397356
rect 80468 397296 80482 397352
rect 80482 397296 80532 397352
rect 80468 397292 80532 397296
rect 83228 397352 83292 397356
rect 83228 397296 83278 397352
rect 83278 397296 83292 397352
rect 83228 397292 83292 397296
rect 86540 397352 86604 397356
rect 86540 397296 86554 397352
rect 86554 397296 86604 397352
rect 86540 397292 86604 397296
rect 87644 397352 87708 397356
rect 87644 397296 87694 397352
rect 87694 397296 87708 397352
rect 87644 397292 87708 397296
rect 88748 397352 88812 397356
rect 88748 397296 88762 397352
rect 88762 397296 88812 397352
rect 88748 397292 88812 397296
rect 91324 397292 91388 397356
rect 93348 397292 93412 397356
rect 96292 397292 96356 397356
rect 98132 397292 98196 397356
rect 99972 397292 100036 397356
rect 100708 397292 100772 397356
rect 101812 397352 101876 397356
rect 101812 397296 101862 397352
rect 101862 397296 101876 397352
rect 101812 397292 101876 397296
rect 102732 397292 102796 397356
rect 103836 397292 103900 397356
rect 105308 397292 105372 397356
rect 106412 397292 106476 397356
rect 109540 397292 109604 397356
rect 111196 397292 111260 397356
rect 114508 397352 114572 397356
rect 114508 397296 114522 397352
rect 114522 397296 114572 397352
rect 114508 397292 114572 397296
rect 115796 397352 115860 397356
rect 115796 397296 115846 397352
rect 115846 397296 115860 397352
rect 115796 397292 115860 397296
rect 118372 397292 118436 397356
rect 136036 397292 136100 397356
rect 138428 397352 138492 397356
rect 138428 397296 138478 397352
rect 138478 397296 138492 397352
rect 138428 397292 138492 397296
rect 150940 397292 151004 397356
rect 183508 397352 183572 397356
rect 183508 397296 183522 397352
rect 183522 397296 183572 397352
rect 183508 397292 183572 397296
rect 237052 397292 237116 397356
rect 239260 397352 239324 397356
rect 239260 397296 239274 397352
rect 239274 397296 239324 397352
rect 239260 397292 239324 397296
rect 241652 397352 241716 397356
rect 241652 397296 241666 397352
rect 241666 397296 241716 397352
rect 241652 397292 241716 397296
rect 242940 397352 243004 397356
rect 242940 397296 242954 397352
rect 242954 397296 243004 397352
rect 242940 397292 243004 397296
rect 245332 397292 245396 397356
rect 248644 397352 248708 397356
rect 248644 397296 248658 397352
rect 248658 397296 248708 397352
rect 248644 397292 248708 397296
rect 250668 397292 250732 397356
rect 253428 397292 253492 397356
rect 253612 397352 253676 397356
rect 253612 397296 253626 397352
rect 253626 397296 253676 397352
rect 253612 397292 253676 397296
rect 256188 397352 256252 397356
rect 256188 397296 256202 397352
rect 256202 397296 256252 397352
rect 256188 397292 256252 397296
rect 260972 397352 261036 397356
rect 260972 397296 260986 397352
rect 260986 397296 261036 397352
rect 260972 397292 261036 397296
rect 262076 397352 262140 397356
rect 262076 397296 262090 397352
rect 262090 397296 262140 397352
rect 262076 397292 262140 397296
rect 263548 397352 263612 397356
rect 263548 397296 263598 397352
rect 263598 397296 263612 397352
rect 263548 397292 263612 397296
rect 271276 397292 271340 397356
rect 273300 397352 273364 397356
rect 273300 397296 273314 397352
rect 273314 397296 273364 397352
rect 273300 397292 273364 397296
rect 274404 397292 274468 397356
rect 275324 397292 275388 397356
rect 276980 397292 277044 397356
rect 278084 397352 278148 397356
rect 278084 397296 278098 397352
rect 278098 397296 278148 397352
rect 278084 397292 278148 397296
rect 290964 397292 291028 397356
rect 293356 397352 293420 397356
rect 293356 397296 293370 397352
rect 293370 397296 293420 397352
rect 293356 397292 293420 397296
rect 298508 397352 298572 397356
rect 298508 397296 298522 397352
rect 298522 397296 298572 397352
rect 298508 397292 298572 397296
rect 308628 397352 308692 397356
rect 308628 397296 308642 397352
rect 308642 397296 308692 397352
rect 308628 397292 308692 397296
rect 311020 397352 311084 397356
rect 311020 397296 311034 397352
rect 311034 397296 311084 397352
rect 311020 397292 311084 397296
rect 313412 397352 313476 397356
rect 313412 397296 313426 397352
rect 313426 397296 313476 397352
rect 313412 397292 313476 397296
rect 343220 397292 343284 397356
rect 96476 397216 96540 397220
rect 96476 397160 96490 397216
rect 96490 397160 96540 397216
rect 96476 397156 96540 397160
rect 98500 397216 98564 397220
rect 98500 397160 98514 397216
rect 98514 397160 98564 397216
rect 98500 397156 98564 397160
rect 103836 397156 103900 397220
rect 113220 397216 113284 397220
rect 113220 397160 113234 397216
rect 113234 397160 113284 397216
rect 113220 397156 113284 397160
rect 263916 397216 263980 397220
rect 263916 397160 263930 397216
rect 263930 397160 263980 397216
rect 263916 397156 263980 397160
rect 273484 397216 273548 397220
rect 273484 397160 273498 397216
rect 273498 397160 273548 397216
rect 273484 397156 273548 397160
rect 258396 396884 258460 396948
rect 76052 396748 76116 396812
rect 81940 396748 82004 396812
rect 84332 396748 84396 396812
rect 88380 396748 88444 396812
rect 90036 396748 90100 396812
rect 93716 396808 93780 396812
rect 93716 396752 93766 396808
rect 93766 396752 93780 396808
rect 93716 396748 93780 396752
rect 94636 396748 94700 396812
rect 97028 396748 97092 396812
rect 101076 396748 101140 396812
rect 106044 396808 106108 396812
rect 106044 396752 106058 396808
rect 106058 396752 106108 396808
rect 106044 396748 106108 396752
rect 107516 396748 107580 396812
rect 108804 396808 108868 396812
rect 108804 396752 108854 396808
rect 108854 396752 108868 396808
rect 108804 396748 108868 396752
rect 111012 396748 111076 396812
rect 112300 396748 112364 396812
rect 117084 396748 117148 396812
rect 118188 396748 118252 396812
rect 119108 396748 119172 396812
rect 120764 396748 120828 396812
rect 123524 396748 123588 396812
rect 125916 396748 125980 396812
rect 128676 396748 128740 396812
rect 131068 396808 131132 396812
rect 131068 396752 131082 396808
rect 131082 396752 131132 396808
rect 131068 396748 131132 396752
rect 133460 396748 133524 396812
rect 140820 396808 140884 396812
rect 140820 396752 140834 396808
rect 140834 396752 140884 396808
rect 140820 396748 140884 396752
rect 143580 396748 143644 396812
rect 145604 396748 145668 396812
rect 148548 396748 148612 396812
rect 154068 396748 154132 396812
rect 155908 396808 155972 396812
rect 155908 396752 155958 396808
rect 155958 396752 155972 396808
rect 155908 396748 155972 396752
rect 158484 396748 158548 396812
rect 160876 396748 160940 396812
rect 163452 396748 163516 396812
rect 166028 396748 166092 396812
rect 183140 396808 183204 396812
rect 183140 396752 183190 396808
rect 183190 396752 183204 396808
rect 183140 396748 183204 396752
rect 238156 396748 238220 396812
rect 240548 396748 240612 396812
rect 244228 396748 244292 396812
rect 246436 396748 246500 396812
rect 248276 396748 248340 396812
rect 250116 396748 250180 396812
rect 251220 396808 251284 396812
rect 251220 396752 251270 396808
rect 251270 396752 251284 396808
rect 251220 396748 251284 396752
rect 254532 396808 254596 396812
rect 254532 396752 254546 396808
rect 254546 396752 254596 396808
rect 254532 396748 254596 396752
rect 255820 396748 255884 396812
rect 256924 396748 256988 396812
rect 258396 396748 258460 396812
rect 259500 396808 259564 396812
rect 259500 396752 259514 396808
rect 259514 396752 259564 396808
rect 259500 396748 259564 396752
rect 262812 396748 262876 396812
rect 265940 396748 266004 396812
rect 266308 396748 266372 396812
rect 268332 396748 268396 396812
rect 269804 396748 269868 396812
rect 270908 396748 270972 396812
rect 272564 396808 272628 396812
rect 272564 396752 272578 396808
rect 272578 396752 272628 396808
rect 272564 396748 272628 396752
rect 276244 396748 276308 396812
rect 278452 396748 278516 396812
rect 279004 396748 279068 396812
rect 280844 396748 280908 396812
rect 283788 396748 283852 396812
rect 285996 396808 286060 396812
rect 285996 396752 286010 396808
rect 286010 396752 286060 396808
rect 285996 396748 286060 396752
rect 288204 396748 288268 396812
rect 295932 396748 295996 396812
rect 303476 396748 303540 396812
rect 305868 396748 305932 396812
rect 318380 396748 318444 396812
rect 320956 396748 321020 396812
rect 323348 396748 323412 396812
rect 343404 396748 343468 396812
rect 77156 396612 77220 396676
rect 90772 396612 90836 396676
rect 91508 396612 91572 396676
rect 108252 396612 108316 396676
rect 115980 396612 116044 396676
rect 247724 396672 247788 396676
rect 247724 396616 247738 396672
rect 247738 396616 247788 396672
rect 247724 396612 247788 396616
rect 252324 396612 252388 396676
rect 260604 396612 260668 396676
rect 267596 396612 267660 396676
rect 268700 396612 268764 396676
rect 219388 393348 219452 393412
rect 219204 392804 219268 392868
rect 219204 383692 219268 383756
rect 219388 383556 219452 383620
rect 219388 374172 219452 374236
rect 219388 373900 219452 373964
rect 219388 364380 219452 364444
rect 219388 364244 219452 364308
rect 219388 354724 219452 354788
rect 219388 354588 219452 354652
rect 219388 345068 219452 345132
rect 219204 344524 219268 344588
rect 219204 335412 219268 335476
rect 219204 335004 219268 335068
rect 219204 325892 219268 325956
rect 219388 325620 219452 325684
rect 219388 316236 219452 316300
rect 219388 315964 219452 316028
rect 219388 306444 219452 306508
rect 219388 306308 219452 306372
rect 219388 296788 219452 296852
rect 219388 296652 219452 296716
rect 219388 287132 219452 287196
rect 219388 286996 219452 287060
rect 219388 277476 219452 277540
rect 219388 277340 219452 277404
rect 219388 267820 219452 267884
rect 219388 267684 219452 267748
rect 219388 258300 219452 258364
rect 219388 257892 219452 257956
rect 219388 248372 219452 248436
rect 219204 247964 219268 248028
rect 219388 238852 219452 238916
rect 218652 238444 218716 238508
rect 218836 238172 218900 238236
rect 219388 238172 219452 238236
rect 226748 236812 226812 236876
rect 219204 235316 219268 235380
rect 226564 235316 226628 235380
rect 219204 235044 219268 235108
rect 218652 234228 218716 234292
rect 226196 234228 226260 234292
rect 218836 234092 218900 234156
rect 226012 234092 226076 234156
rect 228220 233412 228284 233476
rect 224908 231780 224972 231844
rect 224724 231644 224788 231708
rect 223988 230964 224052 231028
rect 219204 230828 219268 230892
rect 223804 230828 223868 230892
rect 219020 228788 219084 228852
rect 224172 228788 224236 228852
rect 224356 228652 224420 228716
rect 225276 228516 225340 228580
rect 60596 226612 60660 226676
rect 60780 226204 60844 226268
rect 60596 225932 60660 225996
rect 60780 225796 60844 225860
rect 223436 226204 223500 226268
rect 223436 225660 223500 225724
rect 226932 225660 226996 225724
rect 226012 147732 226076 147796
rect 226196 143440 226260 143444
rect 226196 143384 226210 143440
rect 226210 143384 226260 143440
rect 226196 143380 226260 143384
rect 226932 126924 226996 126988
rect 226748 113324 226812 113388
rect 228220 111828 228284 111892
rect 226564 74972 226628 75036
rect 224908 70212 224972 70276
rect 225460 70212 225524 70276
rect 224908 60692 224972 60756
rect 225460 60692 225524 60756
rect 223620 60284 223684 60348
rect 225092 60148 225156 60212
rect 224172 59740 224236 59804
rect 227668 59196 227732 59260
rect 223804 59060 223868 59124
rect 223988 59120 224052 59124
rect 223988 59064 224002 59120
rect 224002 59064 224052 59120
rect 223988 59060 224052 59064
rect 224356 59120 224420 59124
rect 224356 59064 224370 59120
rect 224370 59064 224420 59120
rect 224356 59060 224420 59064
rect 227852 58788 227916 58852
rect 226380 58380 226444 58444
rect 224908 57836 224972 57900
rect 224908 57020 224972 57084
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 687454 2414 704282
rect 1794 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 2414 687454
rect 1794 687134 2414 687218
rect 1794 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 2414 687134
rect 1794 651454 2414 686898
rect 1794 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 2414 651454
rect 1794 651134 2414 651218
rect 1794 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 2414 651134
rect 1794 615454 2414 650898
rect 1794 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 2414 615454
rect 1794 615134 2414 615218
rect 1794 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 2414 615134
rect 1794 579454 2414 614898
rect 1794 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 2414 579454
rect 1794 579134 2414 579218
rect 1794 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 2414 579134
rect 1794 543454 2414 578898
rect 1794 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 2414 543454
rect 1794 543134 2414 543218
rect 1794 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 2414 543134
rect 1794 507454 2414 542898
rect 1794 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 2414 507454
rect 1794 507134 2414 507218
rect 1794 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 2414 507134
rect 1794 471454 2414 506898
rect 1794 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 2414 471454
rect 1794 471134 2414 471218
rect 1794 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 2414 471134
rect 1794 435454 2414 470898
rect 1794 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 2414 435454
rect 1794 435134 2414 435218
rect 1794 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 2414 435134
rect 1794 399454 2414 434898
rect 1794 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 2414 399454
rect 1794 399134 2414 399218
rect 1794 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 2414 399134
rect 1794 363454 2414 398898
rect 1794 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 2414 363454
rect 1794 363134 2414 363218
rect 1794 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 2414 363134
rect 1794 327454 2414 362898
rect 1794 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 2414 327454
rect 1794 327134 2414 327218
rect 1794 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 2414 327134
rect 1794 291454 2414 326898
rect 1794 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 2414 291454
rect 1794 291134 2414 291218
rect 1794 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 2414 291134
rect 1794 255454 2414 290898
rect 1794 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 2414 255454
rect 1794 255134 2414 255218
rect 1794 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 2414 255134
rect 1794 219454 2414 254898
rect 1794 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 2414 219454
rect 1794 219134 2414 219218
rect 1794 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 2414 219134
rect 1794 183454 2414 218898
rect 1794 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 2414 183454
rect 1794 183134 2414 183218
rect 1794 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 2414 183134
rect 1794 147454 2414 182898
rect 1794 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 2414 147454
rect 1794 147134 2414 147218
rect 1794 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 2414 147134
rect 1794 111454 2414 146898
rect 1794 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 2414 111454
rect 1794 111134 2414 111218
rect 1794 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 2414 111134
rect 1794 75454 2414 110898
rect 1794 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 2414 75454
rect 1794 75134 2414 75218
rect 1794 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 2414 75134
rect 1794 39454 2414 74898
rect 1794 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 2414 39454
rect 1794 39134 2414 39218
rect 1794 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 2414 39134
rect 1794 3454 2414 38898
rect 1794 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 2414 3454
rect 1794 3134 2414 3218
rect 1794 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 2414 3134
rect 1794 -346 2414 2898
rect 1794 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 2414 -346
rect 1794 -666 2414 -582
rect 1794 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 2414 -666
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect 1794 -1894 2414 -902
rect 5514 691174 6134 706202
rect 5514 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 6134 691174
rect 5514 690854 6134 690938
rect 5514 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 6134 690854
rect 5514 655174 6134 690618
rect 5514 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 6134 655174
rect 5514 654854 6134 654938
rect 5514 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 6134 654854
rect 5514 619174 6134 654618
rect 5514 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 6134 619174
rect 5514 618854 6134 618938
rect 5514 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 6134 618854
rect 5514 583174 6134 618618
rect 5514 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 6134 583174
rect 5514 582854 6134 582938
rect 5514 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 6134 582854
rect 5514 547174 6134 582618
rect 5514 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 6134 547174
rect 5514 546854 6134 546938
rect 5514 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 6134 546854
rect 5514 511174 6134 546618
rect 5514 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 6134 511174
rect 5514 510854 6134 510938
rect 5514 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 6134 510854
rect 5514 475174 6134 510618
rect 5514 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 6134 475174
rect 5514 474854 6134 474938
rect 5514 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 6134 474854
rect 5514 439174 6134 474618
rect 5514 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 6134 439174
rect 5514 438854 6134 438938
rect 5514 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 6134 438854
rect 5514 403174 6134 438618
rect 5514 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 6134 403174
rect 5514 402854 6134 402938
rect 5514 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 6134 402854
rect 5514 367174 6134 402618
rect 5514 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 6134 367174
rect 5514 366854 6134 366938
rect 5514 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 6134 366854
rect 5514 331174 6134 366618
rect 5514 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 6134 331174
rect 5514 330854 6134 330938
rect 5514 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 6134 330854
rect 5514 295174 6134 330618
rect 5514 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 6134 295174
rect 5514 294854 6134 294938
rect 5514 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 6134 294854
rect 5514 259174 6134 294618
rect 5514 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 6134 259174
rect 5514 258854 6134 258938
rect 5514 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 6134 258854
rect 5514 223174 6134 258618
rect 5514 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 6134 223174
rect 5514 222854 6134 222938
rect 5514 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 6134 222854
rect 5514 187174 6134 222618
rect 5514 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 6134 187174
rect 5514 186854 6134 186938
rect 5514 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 6134 186854
rect 5514 151174 6134 186618
rect 5514 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 6134 151174
rect 5514 150854 6134 150938
rect 5514 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 6134 150854
rect 5514 115174 6134 150618
rect 5514 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 6134 115174
rect 5514 114854 6134 114938
rect 5514 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 6134 114854
rect 5514 79174 6134 114618
rect 5514 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 6134 79174
rect 5514 78854 6134 78938
rect 5514 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 6134 78854
rect 5514 43174 6134 78618
rect 5514 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 6134 43174
rect 5514 42854 6134 42938
rect 5514 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 6134 42854
rect 5514 7174 6134 42618
rect 5514 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 6134 7174
rect 5514 6854 6134 6938
rect 5514 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 6134 6854
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 6618
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect 9234 694894 9854 708122
rect 9234 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 9854 694894
rect 9234 694574 9854 694658
rect 9234 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 9854 694574
rect 9234 658894 9854 694338
rect 9234 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 9854 658894
rect 9234 658574 9854 658658
rect 9234 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 9854 658574
rect 9234 622894 9854 658338
rect 9234 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 9854 622894
rect 9234 622574 9854 622658
rect 9234 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 9854 622574
rect 9234 586894 9854 622338
rect 9234 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 9854 586894
rect 9234 586574 9854 586658
rect 9234 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 9854 586574
rect 9234 550894 9854 586338
rect 9234 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 9854 550894
rect 9234 550574 9854 550658
rect 9234 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 9854 550574
rect 9234 514894 9854 550338
rect 9234 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 9854 514894
rect 9234 514574 9854 514658
rect 9234 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 9854 514574
rect 9234 478894 9854 514338
rect 9234 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 9854 478894
rect 9234 478574 9854 478658
rect 9234 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 9854 478574
rect 9234 442894 9854 478338
rect 9234 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 9854 442894
rect 9234 442574 9854 442658
rect 9234 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 9854 442574
rect 9234 406894 9854 442338
rect 9234 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 9854 406894
rect 9234 406574 9854 406658
rect 9234 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 9854 406574
rect 9234 370894 9854 406338
rect 9234 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 9854 370894
rect 9234 370574 9854 370658
rect 9234 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 9854 370574
rect 9234 334894 9854 370338
rect 9234 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 9854 334894
rect 9234 334574 9854 334658
rect 9234 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 9854 334574
rect 9234 298894 9854 334338
rect 9234 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 9854 298894
rect 9234 298574 9854 298658
rect 9234 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 9854 298574
rect 9234 262894 9854 298338
rect 9234 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 9854 262894
rect 9234 262574 9854 262658
rect 9234 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 9854 262574
rect 9234 226894 9854 262338
rect 9234 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 9854 226894
rect 9234 226574 9854 226658
rect 9234 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 9854 226574
rect 9234 190894 9854 226338
rect 9234 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 9854 190894
rect 9234 190574 9854 190658
rect 9234 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 9854 190574
rect 9234 154894 9854 190338
rect 9234 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 9854 154894
rect 9234 154574 9854 154658
rect 9234 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 9854 154574
rect 9234 118894 9854 154338
rect 9234 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 9854 118894
rect 9234 118574 9854 118658
rect 9234 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 9854 118574
rect 9234 82894 9854 118338
rect 9234 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 9854 82894
rect 9234 82574 9854 82658
rect 9234 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 9854 82574
rect 9234 46894 9854 82338
rect 9234 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 9854 46894
rect 9234 46574 9854 46658
rect 9234 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 9854 46574
rect 9234 10894 9854 46338
rect 9234 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 9854 10894
rect 9234 10574 9854 10658
rect 9234 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 9854 10574
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 10338
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect 12954 698614 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 12954 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 13574 698614
rect 12954 698294 13574 698378
rect 12954 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 13574 698294
rect 12954 662614 13574 698058
rect 12954 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 13574 662614
rect 12954 662294 13574 662378
rect 12954 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 13574 662294
rect 12954 626614 13574 662058
rect 12954 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 13574 626614
rect 12954 626294 13574 626378
rect 12954 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 13574 626294
rect 12954 590614 13574 626058
rect 12954 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 13574 590614
rect 12954 590294 13574 590378
rect 12954 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 13574 590294
rect 12954 554614 13574 590058
rect 12954 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 13574 554614
rect 12954 554294 13574 554378
rect 12954 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 13574 554294
rect 12954 518614 13574 554058
rect 12954 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 13574 518614
rect 12954 518294 13574 518378
rect 12954 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 13574 518294
rect 12954 482614 13574 518058
rect 12954 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 13574 482614
rect 12954 482294 13574 482378
rect 12954 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 13574 482294
rect 12954 446614 13574 482058
rect 12954 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 13574 446614
rect 12954 446294 13574 446378
rect 12954 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 13574 446294
rect 12954 410614 13574 446058
rect 12954 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 13574 410614
rect 12954 410294 13574 410378
rect 12954 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 13574 410294
rect 12954 374614 13574 410058
rect 12954 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 13574 374614
rect 12954 374294 13574 374378
rect 12954 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 13574 374294
rect 12954 338614 13574 374058
rect 12954 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 13574 338614
rect 12954 338294 13574 338378
rect 12954 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 13574 338294
rect 12954 302614 13574 338058
rect 12954 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 13574 302614
rect 12954 302294 13574 302378
rect 12954 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 13574 302294
rect 12954 266614 13574 302058
rect 12954 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 13574 266614
rect 12954 266294 13574 266378
rect 12954 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 13574 266294
rect 12954 230614 13574 266058
rect 12954 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 13574 230614
rect 12954 230294 13574 230378
rect 12954 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 13574 230294
rect 12954 194614 13574 230058
rect 12954 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 13574 194614
rect 12954 194294 13574 194378
rect 12954 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 13574 194294
rect 12954 158614 13574 194058
rect 12954 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 13574 158614
rect 12954 158294 13574 158378
rect 12954 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 13574 158294
rect 12954 122614 13574 158058
rect 12954 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 13574 122614
rect 12954 122294 13574 122378
rect 12954 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 13574 122294
rect 12954 86614 13574 122058
rect 12954 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 13574 86614
rect 12954 86294 13574 86378
rect 12954 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 13574 86294
rect 12954 50614 13574 86058
rect 12954 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 13574 50614
rect 12954 50294 13574 50378
rect 12954 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 13574 50294
rect 12954 14614 13574 50058
rect 12954 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 13574 14614
rect 12954 14294 13574 14378
rect 12954 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 13574 14294
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 14058
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 669454 20414 705242
rect 19794 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 20414 669454
rect 19794 669134 20414 669218
rect 19794 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 20414 669134
rect 19794 633454 20414 668898
rect 19794 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 20414 633454
rect 19794 633134 20414 633218
rect 19794 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 20414 633134
rect 19794 597454 20414 632898
rect 19794 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 20414 597454
rect 19794 597134 20414 597218
rect 19794 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 20414 597134
rect 19794 561454 20414 596898
rect 19794 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 20414 561454
rect 19794 561134 20414 561218
rect 19794 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 20414 561134
rect 19794 525454 20414 560898
rect 19794 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 20414 525454
rect 19794 525134 20414 525218
rect 19794 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 20414 525134
rect 19794 489454 20414 524898
rect 19794 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 20414 489454
rect 19794 489134 20414 489218
rect 19794 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 20414 489134
rect 19794 453454 20414 488898
rect 19794 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 20414 453454
rect 19794 453134 20414 453218
rect 19794 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 20414 453134
rect 19794 417454 20414 452898
rect 19794 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 20414 417454
rect 19794 417134 20414 417218
rect 19794 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 20414 417134
rect 19794 381454 20414 416898
rect 19794 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 20414 381454
rect 19794 381134 20414 381218
rect 19794 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 20414 381134
rect 19794 345454 20414 380898
rect 19794 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 20414 345454
rect 19794 345134 20414 345218
rect 19794 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 20414 345134
rect 19794 309454 20414 344898
rect 19794 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 20414 309454
rect 19794 309134 20414 309218
rect 19794 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 20414 309134
rect 19794 273454 20414 308898
rect 19794 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 20414 273454
rect 19794 273134 20414 273218
rect 19794 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 20414 273134
rect 19794 237454 20414 272898
rect 19794 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 20414 237454
rect 19794 237134 20414 237218
rect 19794 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 20414 237134
rect 19794 201454 20414 236898
rect 19794 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 20414 201454
rect 19794 201134 20414 201218
rect 19794 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 20414 201134
rect 19794 165454 20414 200898
rect 19794 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 20414 165454
rect 19794 165134 20414 165218
rect 19794 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 20414 165134
rect 19794 129454 20414 164898
rect 19794 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 20414 129454
rect 19794 129134 20414 129218
rect 19794 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 20414 129134
rect 19794 93454 20414 128898
rect 19794 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 20414 93454
rect 19794 93134 20414 93218
rect 19794 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 20414 93134
rect 19794 57454 20414 92898
rect 19794 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 20414 57454
rect 19794 57134 20414 57218
rect 19794 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 20414 57134
rect 19794 21454 20414 56898
rect 19794 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 20414 21454
rect 19794 21134 20414 21218
rect 19794 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 20414 21134
rect 19794 -1306 20414 20898
rect 19794 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 20414 -1306
rect 19794 -1626 20414 -1542
rect 19794 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 20414 -1626
rect 19794 -1894 20414 -1862
rect 23514 673174 24134 707162
rect 23514 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 24134 673174
rect 23514 672854 24134 672938
rect 23514 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 24134 672854
rect 23514 637174 24134 672618
rect 23514 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 24134 637174
rect 23514 636854 24134 636938
rect 23514 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 24134 636854
rect 23514 601174 24134 636618
rect 23514 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 24134 601174
rect 23514 600854 24134 600938
rect 23514 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 24134 600854
rect 23514 565174 24134 600618
rect 23514 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 24134 565174
rect 23514 564854 24134 564938
rect 23514 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 24134 564854
rect 23514 529174 24134 564618
rect 23514 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 24134 529174
rect 23514 528854 24134 528938
rect 23514 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 24134 528854
rect 23514 493174 24134 528618
rect 23514 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 24134 493174
rect 23514 492854 24134 492938
rect 23514 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 24134 492854
rect 23514 457174 24134 492618
rect 23514 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 24134 457174
rect 23514 456854 24134 456938
rect 23514 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 24134 456854
rect 23514 421174 24134 456618
rect 23514 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 24134 421174
rect 23514 420854 24134 420938
rect 23514 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 24134 420854
rect 23514 385174 24134 420618
rect 23514 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 24134 385174
rect 23514 384854 24134 384938
rect 23514 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 24134 384854
rect 23514 349174 24134 384618
rect 23514 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 24134 349174
rect 23514 348854 24134 348938
rect 23514 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 24134 348854
rect 23514 313174 24134 348618
rect 23514 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 24134 313174
rect 23514 312854 24134 312938
rect 23514 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 24134 312854
rect 23514 277174 24134 312618
rect 23514 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 24134 277174
rect 23514 276854 24134 276938
rect 23514 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 24134 276854
rect 23514 241174 24134 276618
rect 23514 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 24134 241174
rect 23514 240854 24134 240938
rect 23514 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 24134 240854
rect 23514 205174 24134 240618
rect 23514 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 24134 205174
rect 23514 204854 24134 204938
rect 23514 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 24134 204854
rect 23514 169174 24134 204618
rect 23514 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 24134 169174
rect 23514 168854 24134 168938
rect 23514 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 24134 168854
rect 23514 133174 24134 168618
rect 23514 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 24134 133174
rect 23514 132854 24134 132938
rect 23514 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 24134 132854
rect 23514 97174 24134 132618
rect 23514 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 24134 97174
rect 23514 96854 24134 96938
rect 23514 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 24134 96854
rect 23514 61174 24134 96618
rect 23514 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 24134 61174
rect 23514 60854 24134 60938
rect 23514 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 24134 60854
rect 23514 25174 24134 60618
rect 23514 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 24134 25174
rect 23514 24854 24134 24938
rect 23514 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 24134 24854
rect 23514 -3226 24134 24618
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 676894 27854 709082
rect 27234 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 27854 676894
rect 27234 676574 27854 676658
rect 27234 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 27854 676574
rect 27234 640894 27854 676338
rect 27234 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 27854 640894
rect 27234 640574 27854 640658
rect 27234 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 27854 640574
rect 27234 604894 27854 640338
rect 27234 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 27854 604894
rect 27234 604574 27854 604658
rect 27234 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 27854 604574
rect 27234 568894 27854 604338
rect 27234 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 27854 568894
rect 27234 568574 27854 568658
rect 27234 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 27854 568574
rect 27234 532894 27854 568338
rect 27234 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 27854 532894
rect 27234 532574 27854 532658
rect 27234 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 27854 532574
rect 27234 496894 27854 532338
rect 27234 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 27854 496894
rect 27234 496574 27854 496658
rect 27234 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 27854 496574
rect 27234 460894 27854 496338
rect 27234 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 27854 460894
rect 27234 460574 27854 460658
rect 27234 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 27854 460574
rect 27234 424894 27854 460338
rect 27234 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 27854 424894
rect 27234 424574 27854 424658
rect 27234 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 27854 424574
rect 27234 388894 27854 424338
rect 27234 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 27854 388894
rect 27234 388574 27854 388658
rect 27234 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 27854 388574
rect 27234 352894 27854 388338
rect 27234 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 27854 352894
rect 27234 352574 27854 352658
rect 27234 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 27854 352574
rect 27234 316894 27854 352338
rect 27234 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 27854 316894
rect 27234 316574 27854 316658
rect 27234 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 27854 316574
rect 27234 280894 27854 316338
rect 27234 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 27854 280894
rect 27234 280574 27854 280658
rect 27234 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 27854 280574
rect 27234 244894 27854 280338
rect 27234 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 27854 244894
rect 27234 244574 27854 244658
rect 27234 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 27854 244574
rect 27234 208894 27854 244338
rect 27234 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 27854 208894
rect 27234 208574 27854 208658
rect 27234 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 27854 208574
rect 27234 172894 27854 208338
rect 27234 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 27854 172894
rect 27234 172574 27854 172658
rect 27234 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 27854 172574
rect 27234 136894 27854 172338
rect 27234 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 27854 136894
rect 27234 136574 27854 136658
rect 27234 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 27854 136574
rect 27234 100894 27854 136338
rect 27234 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 27854 100894
rect 27234 100574 27854 100658
rect 27234 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 27854 100574
rect 27234 64894 27854 100338
rect 27234 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 27854 64894
rect 27234 64574 27854 64658
rect 27234 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 27854 64574
rect 27234 28894 27854 64338
rect 27234 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 27854 28894
rect 27234 28574 27854 28658
rect 27234 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 27854 28574
rect 27234 -5146 27854 28338
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 30954 680614 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 30954 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 31574 680614
rect 30954 680294 31574 680378
rect 30954 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 31574 680294
rect 30954 644614 31574 680058
rect 30954 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 31574 644614
rect 30954 644294 31574 644378
rect 30954 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 31574 644294
rect 30954 608614 31574 644058
rect 30954 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 31574 608614
rect 30954 608294 31574 608378
rect 30954 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 31574 608294
rect 30954 572614 31574 608058
rect 30954 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 31574 572614
rect 30954 572294 31574 572378
rect 30954 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 31574 572294
rect 30954 536614 31574 572058
rect 30954 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 31574 536614
rect 30954 536294 31574 536378
rect 30954 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 31574 536294
rect 30954 500614 31574 536058
rect 30954 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 31574 500614
rect 30954 500294 31574 500378
rect 30954 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 31574 500294
rect 30954 464614 31574 500058
rect 30954 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 31574 464614
rect 30954 464294 31574 464378
rect 30954 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 31574 464294
rect 30954 428614 31574 464058
rect 30954 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 31574 428614
rect 30954 428294 31574 428378
rect 30954 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 31574 428294
rect 30954 392614 31574 428058
rect 30954 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 31574 392614
rect 30954 392294 31574 392378
rect 30954 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 31574 392294
rect 30954 356614 31574 392058
rect 30954 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 31574 356614
rect 30954 356294 31574 356378
rect 30954 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 31574 356294
rect 30954 320614 31574 356058
rect 30954 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 31574 320614
rect 30954 320294 31574 320378
rect 30954 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 31574 320294
rect 30954 284614 31574 320058
rect 30954 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 31574 284614
rect 30954 284294 31574 284378
rect 30954 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 31574 284294
rect 30954 248614 31574 284058
rect 30954 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 31574 248614
rect 30954 248294 31574 248378
rect 30954 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 31574 248294
rect 30954 212614 31574 248058
rect 30954 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 31574 212614
rect 30954 212294 31574 212378
rect 30954 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 31574 212294
rect 30954 176614 31574 212058
rect 30954 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 31574 176614
rect 30954 176294 31574 176378
rect 30954 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 31574 176294
rect 30954 140614 31574 176058
rect 30954 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 31574 140614
rect 30954 140294 31574 140378
rect 30954 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 31574 140294
rect 30954 104614 31574 140058
rect 30954 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 31574 104614
rect 30954 104294 31574 104378
rect 30954 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 31574 104294
rect 30954 68614 31574 104058
rect 30954 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 31574 68614
rect 30954 68294 31574 68378
rect 30954 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 31574 68294
rect 30954 32614 31574 68058
rect 30954 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 31574 32614
rect 30954 32294 31574 32378
rect 30954 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 31574 32294
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 32058
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 687454 38414 704282
rect 37794 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 38414 687454
rect 37794 687134 38414 687218
rect 37794 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 38414 687134
rect 37794 651454 38414 686898
rect 37794 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 38414 651454
rect 37794 651134 38414 651218
rect 37794 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 38414 651134
rect 37794 615454 38414 650898
rect 37794 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 38414 615454
rect 37794 615134 38414 615218
rect 37794 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 38414 615134
rect 37794 579454 38414 614898
rect 37794 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 38414 579454
rect 37794 579134 38414 579218
rect 37794 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 38414 579134
rect 37794 543454 38414 578898
rect 37794 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 38414 543454
rect 37794 543134 38414 543218
rect 37794 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 38414 543134
rect 37794 507454 38414 542898
rect 37794 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 38414 507454
rect 37794 507134 38414 507218
rect 37794 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 38414 507134
rect 37794 471454 38414 506898
rect 37794 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 38414 471454
rect 37794 471134 38414 471218
rect 37794 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 38414 471134
rect 37794 435454 38414 470898
rect 37794 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 38414 435454
rect 37794 435134 38414 435218
rect 37794 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 38414 435134
rect 37794 399454 38414 434898
rect 37794 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 38414 399454
rect 37794 399134 38414 399218
rect 37794 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 38414 399134
rect 37794 363454 38414 398898
rect 37794 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 38414 363454
rect 37794 363134 38414 363218
rect 37794 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 38414 363134
rect 37794 327454 38414 362898
rect 37794 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 38414 327454
rect 37794 327134 38414 327218
rect 37794 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 38414 327134
rect 37794 291454 38414 326898
rect 37794 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 38414 291454
rect 37794 291134 38414 291218
rect 37794 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 38414 291134
rect 37794 255454 38414 290898
rect 37794 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 38414 255454
rect 37794 255134 38414 255218
rect 37794 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 38414 255134
rect 37794 219454 38414 254898
rect 37794 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 38414 219454
rect 37794 219134 38414 219218
rect 37794 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 38414 219134
rect 37794 183454 38414 218898
rect 37794 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 38414 183454
rect 37794 183134 38414 183218
rect 37794 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 38414 183134
rect 37794 147454 38414 182898
rect 37794 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 38414 147454
rect 37794 147134 38414 147218
rect 37794 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 38414 147134
rect 37794 111454 38414 146898
rect 37794 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 38414 111454
rect 37794 111134 38414 111218
rect 37794 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 38414 111134
rect 37794 75454 38414 110898
rect 37794 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 38414 75454
rect 37794 75134 38414 75218
rect 37794 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 38414 75134
rect 37794 39454 38414 74898
rect 37794 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 38414 39454
rect 37794 39134 38414 39218
rect 37794 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 38414 39134
rect 37794 3454 38414 38898
rect 37794 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 38414 3454
rect 37794 3134 38414 3218
rect 37794 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 38414 3134
rect 37794 -346 38414 2898
rect 37794 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 38414 -346
rect 37794 -666 38414 -582
rect 37794 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 38414 -666
rect 37794 -1894 38414 -902
rect 41514 691174 42134 706202
rect 41514 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 42134 691174
rect 41514 690854 42134 690938
rect 41514 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 42134 690854
rect 41514 655174 42134 690618
rect 41514 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 42134 655174
rect 41514 654854 42134 654938
rect 41514 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 42134 654854
rect 41514 619174 42134 654618
rect 41514 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 42134 619174
rect 41514 618854 42134 618938
rect 41514 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 42134 618854
rect 41514 583174 42134 618618
rect 41514 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 42134 583174
rect 41514 582854 42134 582938
rect 41514 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 42134 582854
rect 41514 547174 42134 582618
rect 41514 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 42134 547174
rect 41514 546854 42134 546938
rect 41514 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 42134 546854
rect 41514 511174 42134 546618
rect 41514 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 42134 511174
rect 41514 510854 42134 510938
rect 41514 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 42134 510854
rect 41514 475174 42134 510618
rect 41514 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 42134 475174
rect 41514 474854 42134 474938
rect 41514 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 42134 474854
rect 41514 439174 42134 474618
rect 41514 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 42134 439174
rect 41514 438854 42134 438938
rect 41514 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 42134 438854
rect 41514 403174 42134 438618
rect 41514 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 42134 403174
rect 41514 402854 42134 402938
rect 41514 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 42134 402854
rect 41514 367174 42134 402618
rect 41514 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 42134 367174
rect 41514 366854 42134 366938
rect 41514 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 42134 366854
rect 41514 331174 42134 366618
rect 41514 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 42134 331174
rect 41514 330854 42134 330938
rect 41514 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 42134 330854
rect 41514 295174 42134 330618
rect 41514 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 42134 295174
rect 41514 294854 42134 294938
rect 41514 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 42134 294854
rect 41514 259174 42134 294618
rect 41514 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 42134 259174
rect 41514 258854 42134 258938
rect 41514 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 42134 258854
rect 41514 223174 42134 258618
rect 41514 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 42134 223174
rect 41514 222854 42134 222938
rect 41514 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 42134 222854
rect 41514 187174 42134 222618
rect 41514 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 42134 187174
rect 41514 186854 42134 186938
rect 41514 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 42134 186854
rect 41514 151174 42134 186618
rect 41514 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 42134 151174
rect 41514 150854 42134 150938
rect 41514 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 42134 150854
rect 41514 115174 42134 150618
rect 41514 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 42134 115174
rect 41514 114854 42134 114938
rect 41514 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 42134 114854
rect 41514 79174 42134 114618
rect 41514 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 42134 79174
rect 41514 78854 42134 78938
rect 41514 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 42134 78854
rect 41514 43174 42134 78618
rect 41514 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 42134 43174
rect 41514 42854 42134 42938
rect 41514 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 42134 42854
rect 41514 7174 42134 42618
rect 41514 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 42134 7174
rect 41514 6854 42134 6938
rect 41514 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 42134 6854
rect 41514 -2266 42134 6618
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 694894 45854 708122
rect 45234 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 45854 694894
rect 45234 694574 45854 694658
rect 45234 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 45854 694574
rect 45234 658894 45854 694338
rect 45234 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 45854 658894
rect 45234 658574 45854 658658
rect 45234 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 45854 658574
rect 45234 622894 45854 658338
rect 45234 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 45854 622894
rect 45234 622574 45854 622658
rect 45234 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 45854 622574
rect 45234 586894 45854 622338
rect 45234 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 45854 586894
rect 45234 586574 45854 586658
rect 45234 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 45854 586574
rect 45234 550894 45854 586338
rect 45234 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 45854 550894
rect 45234 550574 45854 550658
rect 45234 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 45854 550574
rect 45234 514894 45854 550338
rect 45234 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 45854 514894
rect 45234 514574 45854 514658
rect 45234 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 45854 514574
rect 45234 478894 45854 514338
rect 45234 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 45854 478894
rect 45234 478574 45854 478658
rect 45234 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 45854 478574
rect 45234 442894 45854 478338
rect 45234 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 45854 442894
rect 45234 442574 45854 442658
rect 45234 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 45854 442574
rect 45234 406894 45854 442338
rect 45234 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 45854 406894
rect 45234 406574 45854 406658
rect 45234 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 45854 406574
rect 45234 370894 45854 406338
rect 45234 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 45854 370894
rect 45234 370574 45854 370658
rect 45234 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 45854 370574
rect 45234 334894 45854 370338
rect 45234 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 45854 334894
rect 45234 334574 45854 334658
rect 45234 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 45854 334574
rect 45234 298894 45854 334338
rect 45234 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 45854 298894
rect 45234 298574 45854 298658
rect 45234 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 45854 298574
rect 45234 262894 45854 298338
rect 45234 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 45854 262894
rect 45234 262574 45854 262658
rect 45234 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 45854 262574
rect 45234 226894 45854 262338
rect 45234 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 45854 226894
rect 45234 226574 45854 226658
rect 45234 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 45854 226574
rect 45234 190894 45854 226338
rect 45234 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 45854 190894
rect 45234 190574 45854 190658
rect 45234 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 45854 190574
rect 45234 154894 45854 190338
rect 45234 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 45854 154894
rect 45234 154574 45854 154658
rect 45234 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 45854 154574
rect 45234 118894 45854 154338
rect 45234 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 45854 118894
rect 45234 118574 45854 118658
rect 45234 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 45854 118574
rect 45234 82894 45854 118338
rect 45234 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 45854 82894
rect 45234 82574 45854 82658
rect 45234 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 45854 82574
rect 45234 46894 45854 82338
rect 45234 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 45854 46894
rect 45234 46574 45854 46658
rect 45234 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 45854 46574
rect 45234 10894 45854 46338
rect 45234 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 45854 10894
rect 45234 10574 45854 10658
rect 45234 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 45854 10574
rect 45234 -4186 45854 10338
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 48954 698614 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 48954 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 49574 698614
rect 48954 698294 49574 698378
rect 48954 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 49574 698294
rect 48954 662614 49574 698058
rect 48954 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 49574 662614
rect 48954 662294 49574 662378
rect 48954 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 49574 662294
rect 48954 626614 49574 662058
rect 48954 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 49574 626614
rect 48954 626294 49574 626378
rect 48954 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 49574 626294
rect 48954 590614 49574 626058
rect 48954 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 49574 590614
rect 48954 590294 49574 590378
rect 48954 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 49574 590294
rect 48954 554614 49574 590058
rect 48954 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 49574 554614
rect 48954 554294 49574 554378
rect 48954 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 49574 554294
rect 48954 518614 49574 554058
rect 48954 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 49574 518614
rect 48954 518294 49574 518378
rect 48954 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 49574 518294
rect 48954 482614 49574 518058
rect 48954 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 49574 482614
rect 48954 482294 49574 482378
rect 48954 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 49574 482294
rect 48954 446614 49574 482058
rect 48954 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 49574 446614
rect 48954 446294 49574 446378
rect 48954 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 49574 446294
rect 48954 410614 49574 446058
rect 48954 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 49574 410614
rect 48954 410294 49574 410378
rect 48954 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 49574 410294
rect 48954 374614 49574 410058
rect 48954 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 49574 374614
rect 48954 374294 49574 374378
rect 48954 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 49574 374294
rect 48954 338614 49574 374058
rect 48954 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 49574 338614
rect 48954 338294 49574 338378
rect 48954 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 49574 338294
rect 48954 302614 49574 338058
rect 48954 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 49574 302614
rect 48954 302294 49574 302378
rect 48954 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 49574 302294
rect 48954 266614 49574 302058
rect 48954 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 49574 266614
rect 48954 266294 49574 266378
rect 48954 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 49574 266294
rect 48954 230614 49574 266058
rect 48954 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 49574 230614
rect 48954 230294 49574 230378
rect 48954 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 49574 230294
rect 48954 194614 49574 230058
rect 48954 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 49574 194614
rect 48954 194294 49574 194378
rect 48954 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 49574 194294
rect 48954 158614 49574 194058
rect 48954 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 49574 158614
rect 48954 158294 49574 158378
rect 48954 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 49574 158294
rect 48954 122614 49574 158058
rect 48954 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 49574 122614
rect 48954 122294 49574 122378
rect 48954 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 49574 122294
rect 48954 86614 49574 122058
rect 48954 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 49574 86614
rect 48954 86294 49574 86378
rect 48954 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 49574 86294
rect 48954 50614 49574 86058
rect 48954 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 49574 50614
rect 48954 50294 49574 50378
rect 48954 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 49574 50294
rect 48954 14614 49574 50058
rect 48954 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 49574 14614
rect 48954 14294 49574 14378
rect 48954 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 49574 14294
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 14058
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 669454 56414 705242
rect 55794 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 56414 669454
rect 55794 669134 56414 669218
rect 55794 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 56414 669134
rect 55794 633454 56414 668898
rect 55794 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 56414 633454
rect 55794 633134 56414 633218
rect 55794 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 56414 633134
rect 55794 597454 56414 632898
rect 55794 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 56414 597454
rect 55794 597134 56414 597218
rect 55794 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 56414 597134
rect 55794 561454 56414 596898
rect 55794 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 56414 561454
rect 55794 561134 56414 561218
rect 55794 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 56414 561134
rect 55794 525454 56414 560898
rect 55794 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 56414 525454
rect 55794 525134 56414 525218
rect 55794 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 56414 525134
rect 55794 489454 56414 524898
rect 55794 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 56414 489454
rect 55794 489134 56414 489218
rect 55794 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 56414 489134
rect 55794 453454 56414 488898
rect 59514 673174 60134 707162
rect 59514 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 60134 673174
rect 59514 672854 60134 672938
rect 59514 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 60134 672854
rect 59514 637174 60134 672618
rect 59514 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 60134 637174
rect 59514 636854 60134 636938
rect 59514 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 60134 636854
rect 59514 601174 60134 636618
rect 59514 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 60134 601174
rect 59514 600854 60134 600938
rect 59514 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 60134 600854
rect 59514 565174 60134 600618
rect 59514 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 60134 565174
rect 59514 564854 60134 564938
rect 59514 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 60134 564854
rect 59514 529174 60134 564618
rect 59514 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 60134 529174
rect 59514 528854 60134 528938
rect 59514 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 60134 528854
rect 59514 493174 60134 528618
rect 59514 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 60134 493174
rect 59514 492854 60134 492938
rect 59514 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 60134 492854
rect 59514 485308 60134 492618
rect 63234 676894 63854 709082
rect 63234 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 63854 676894
rect 63234 676574 63854 676658
rect 63234 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 63854 676574
rect 63234 640894 63854 676338
rect 63234 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 63854 640894
rect 63234 640574 63854 640658
rect 63234 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 63854 640574
rect 63234 604894 63854 640338
rect 63234 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 63854 604894
rect 63234 604574 63854 604658
rect 63234 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 63854 604574
rect 63234 568894 63854 604338
rect 63234 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 63854 568894
rect 63234 568574 63854 568658
rect 63234 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 63854 568574
rect 63234 532894 63854 568338
rect 63234 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 63854 532894
rect 63234 532574 63854 532658
rect 63234 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 63854 532574
rect 63234 496894 63854 532338
rect 63234 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 63854 496894
rect 63234 496574 63854 496658
rect 63234 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 63854 496574
rect 63234 485308 63854 496338
rect 66954 680614 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 66954 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 67574 680614
rect 66954 680294 67574 680378
rect 66954 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 67574 680294
rect 66954 644614 67574 680058
rect 66954 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 67574 644614
rect 66954 644294 67574 644378
rect 66954 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 67574 644294
rect 66954 608614 67574 644058
rect 66954 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 67574 608614
rect 66954 608294 67574 608378
rect 66954 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 67574 608294
rect 66954 572614 67574 608058
rect 66954 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 67574 572614
rect 66954 572294 67574 572378
rect 66954 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 67574 572294
rect 66954 536614 67574 572058
rect 66954 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 67574 536614
rect 66954 536294 67574 536378
rect 66954 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 67574 536294
rect 66954 500614 67574 536058
rect 66954 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 67574 500614
rect 66954 500294 67574 500378
rect 66954 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 67574 500294
rect 66954 485308 67574 500058
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 687454 74414 704282
rect 73794 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 74414 687454
rect 73794 687134 74414 687218
rect 73794 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 74414 687134
rect 73794 651454 74414 686898
rect 73794 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 74414 651454
rect 73794 651134 74414 651218
rect 73794 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 74414 651134
rect 73794 615454 74414 650898
rect 73794 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 74414 615454
rect 73794 615134 74414 615218
rect 73794 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 74414 615134
rect 73794 579454 74414 614898
rect 73794 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 74414 579454
rect 73794 579134 74414 579218
rect 73794 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 74414 579134
rect 73794 543454 74414 578898
rect 73794 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 74414 543454
rect 73794 543134 74414 543218
rect 73794 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 74414 543134
rect 73794 507454 74414 542898
rect 73794 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 74414 507454
rect 73794 507134 74414 507218
rect 73794 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 74414 507134
rect 73794 485308 74414 506898
rect 77514 691174 78134 706202
rect 77514 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 78134 691174
rect 77514 690854 78134 690938
rect 77514 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 78134 690854
rect 77514 655174 78134 690618
rect 77514 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 78134 655174
rect 77514 654854 78134 654938
rect 77514 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 78134 654854
rect 77514 619174 78134 654618
rect 77514 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 78134 619174
rect 77514 618854 78134 618938
rect 77514 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 78134 618854
rect 77514 583174 78134 618618
rect 77514 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 78134 583174
rect 77514 582854 78134 582938
rect 77514 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 78134 582854
rect 77514 547174 78134 582618
rect 77514 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 78134 547174
rect 77514 546854 78134 546938
rect 77514 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 78134 546854
rect 77514 511174 78134 546618
rect 77514 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 78134 511174
rect 77514 510854 78134 510938
rect 77514 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 78134 510854
rect 77514 485308 78134 510618
rect 81234 694894 81854 708122
rect 81234 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 81854 694894
rect 81234 694574 81854 694658
rect 81234 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 81854 694574
rect 81234 658894 81854 694338
rect 81234 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 81854 658894
rect 81234 658574 81854 658658
rect 81234 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 81854 658574
rect 81234 622894 81854 658338
rect 81234 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 81854 622894
rect 81234 622574 81854 622658
rect 81234 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 81854 622574
rect 81234 586894 81854 622338
rect 81234 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 81854 586894
rect 81234 586574 81854 586658
rect 81234 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 81854 586574
rect 81234 550894 81854 586338
rect 81234 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 81854 550894
rect 81234 550574 81854 550658
rect 81234 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 81854 550574
rect 81234 514894 81854 550338
rect 81234 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 81854 514894
rect 81234 514574 81854 514658
rect 81234 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 81854 514574
rect 81234 485308 81854 514338
rect 84954 698614 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 84954 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 85574 698614
rect 84954 698294 85574 698378
rect 84954 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 85574 698294
rect 84954 662614 85574 698058
rect 84954 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 85574 662614
rect 84954 662294 85574 662378
rect 84954 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 85574 662294
rect 84954 626614 85574 662058
rect 84954 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 85574 626614
rect 84954 626294 85574 626378
rect 84954 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 85574 626294
rect 84954 590614 85574 626058
rect 84954 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 85574 590614
rect 84954 590294 85574 590378
rect 84954 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 85574 590294
rect 84954 554614 85574 590058
rect 84954 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 85574 554614
rect 84954 554294 85574 554378
rect 84954 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 85574 554294
rect 84954 518614 85574 554058
rect 84954 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 85574 518614
rect 84954 518294 85574 518378
rect 84954 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 85574 518294
rect 84954 485308 85574 518058
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 669454 92414 705242
rect 91794 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 92414 669454
rect 91794 669134 92414 669218
rect 91794 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 92414 669134
rect 91794 633454 92414 668898
rect 91794 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 92414 633454
rect 91794 633134 92414 633218
rect 91794 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 92414 633134
rect 91794 597454 92414 632898
rect 91794 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 92414 597454
rect 91794 597134 92414 597218
rect 91794 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 92414 597134
rect 91794 561454 92414 596898
rect 91794 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 92414 561454
rect 91794 561134 92414 561218
rect 91794 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 92414 561134
rect 91794 525454 92414 560898
rect 91794 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 92414 525454
rect 91794 525134 92414 525218
rect 91794 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 92414 525134
rect 91794 489454 92414 524898
rect 91794 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 92414 489454
rect 91794 489134 92414 489218
rect 91794 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 92414 489134
rect 90955 487116 91021 487117
rect 90955 487052 90956 487116
rect 91020 487052 91021 487116
rect 90955 487051 91021 487052
rect 88747 485892 88813 485893
rect 88747 485828 88748 485892
rect 88812 485828 88813 485892
rect 88747 485827 88813 485828
rect 88750 483850 88810 485827
rect 88704 483790 88810 483850
rect 90958 483850 91018 487051
rect 91794 485308 92414 488898
rect 95514 673174 96134 707162
rect 95514 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 96134 673174
rect 95514 672854 96134 672938
rect 95514 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 96134 672854
rect 95514 637174 96134 672618
rect 95514 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 96134 637174
rect 95514 636854 96134 636938
rect 95514 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 96134 636854
rect 95514 601174 96134 636618
rect 95514 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 96134 601174
rect 95514 600854 96134 600938
rect 95514 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 96134 600854
rect 95514 565174 96134 600618
rect 95514 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 96134 565174
rect 95514 564854 96134 564938
rect 95514 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 96134 564854
rect 95514 529174 96134 564618
rect 95514 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 96134 529174
rect 95514 528854 96134 528938
rect 95514 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 96134 528854
rect 95514 493174 96134 528618
rect 95514 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 96134 493174
rect 95514 492854 96134 492938
rect 95514 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 96134 492854
rect 93347 486028 93413 486029
rect 93347 485964 93348 486028
rect 93412 485964 93413 486028
rect 93347 485963 93413 485964
rect 93350 483850 93410 485963
rect 95514 485308 96134 492618
rect 99234 676894 99854 709082
rect 99234 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 99854 676894
rect 99234 676574 99854 676658
rect 99234 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 99854 676574
rect 99234 640894 99854 676338
rect 99234 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 99854 640894
rect 99234 640574 99854 640658
rect 99234 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 99854 640574
rect 99234 604894 99854 640338
rect 99234 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 99854 604894
rect 99234 604574 99854 604658
rect 99234 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 99854 604574
rect 99234 568894 99854 604338
rect 99234 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 99854 568894
rect 99234 568574 99854 568658
rect 99234 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 99854 568574
rect 99234 532894 99854 568338
rect 99234 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 99854 532894
rect 99234 532574 99854 532658
rect 99234 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 99854 532574
rect 99234 496894 99854 532338
rect 99234 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 99854 496894
rect 99234 496574 99854 496658
rect 99234 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 99854 496574
rect 98499 486028 98565 486029
rect 98499 485964 98500 486028
rect 98564 485964 98565 486028
rect 98499 485963 98565 485964
rect 98502 483850 98562 485963
rect 99234 485308 99854 496338
rect 102954 680614 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 102954 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 103574 680614
rect 102954 680294 103574 680378
rect 102954 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 103574 680294
rect 102954 644614 103574 680058
rect 102954 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 103574 644614
rect 102954 644294 103574 644378
rect 102954 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 103574 644294
rect 102954 608614 103574 644058
rect 102954 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 103574 608614
rect 102954 608294 103574 608378
rect 102954 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 103574 608294
rect 102954 572614 103574 608058
rect 102954 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 103574 572614
rect 102954 572294 103574 572378
rect 102954 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 103574 572294
rect 102954 536614 103574 572058
rect 102954 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 103574 536614
rect 102954 536294 103574 536378
rect 102954 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 103574 536294
rect 102954 500614 103574 536058
rect 102954 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 103574 500614
rect 102954 500294 103574 500378
rect 102954 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 103574 500294
rect 101075 486572 101141 486573
rect 101075 486508 101076 486572
rect 101140 486508 101141 486572
rect 101075 486507 101141 486508
rect 90958 483790 91076 483850
rect 93350 483790 93524 483850
rect 88704 483202 88764 483790
rect 91016 483202 91076 483790
rect 93464 483202 93524 483790
rect 98496 483790 98562 483850
rect 101078 483850 101138 486507
rect 102954 485308 103574 500058
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 687454 110414 704282
rect 109794 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 110414 687454
rect 109794 687134 110414 687218
rect 109794 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 110414 687134
rect 109794 651454 110414 686898
rect 109794 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 110414 651454
rect 109794 651134 110414 651218
rect 109794 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 110414 651134
rect 109794 615454 110414 650898
rect 109794 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 110414 615454
rect 109794 615134 110414 615218
rect 109794 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 110414 615134
rect 109794 579454 110414 614898
rect 109794 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 110414 579454
rect 109794 579134 110414 579218
rect 109794 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 110414 579134
rect 109794 543454 110414 578898
rect 109794 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 110414 543454
rect 109794 543134 110414 543218
rect 109794 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 110414 543134
rect 109794 507454 110414 542898
rect 109794 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 110414 507454
rect 109794 507134 110414 507218
rect 109794 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 110414 507134
rect 103835 486572 103901 486573
rect 103835 486570 103836 486572
rect 103654 486510 103836 486570
rect 103654 483850 103714 486510
rect 103835 486508 103836 486510
rect 103900 486508 103901 486572
rect 103835 486507 103901 486508
rect 108619 486572 108685 486573
rect 108619 486508 108620 486572
rect 108684 486508 108685 486572
rect 108619 486507 108685 486508
rect 106227 486164 106293 486165
rect 106227 486100 106228 486164
rect 106292 486100 106293 486164
rect 106227 486099 106293 486100
rect 106230 483850 106290 486099
rect 108622 483850 108682 486507
rect 109794 485308 110414 506898
rect 113514 691174 114134 706202
rect 113514 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 114134 691174
rect 113514 690854 114134 690938
rect 113514 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 114134 690854
rect 113514 655174 114134 690618
rect 113514 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 114134 655174
rect 113514 654854 114134 654938
rect 113514 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 114134 654854
rect 113514 619174 114134 654618
rect 113514 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 114134 619174
rect 113514 618854 114134 618938
rect 113514 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 114134 618854
rect 113514 583174 114134 618618
rect 113514 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 114134 583174
rect 113514 582854 114134 582938
rect 113514 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 114134 582854
rect 113514 547174 114134 582618
rect 113514 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 114134 547174
rect 113514 546854 114134 546938
rect 113514 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 114134 546854
rect 113514 511174 114134 546618
rect 113514 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 114134 511174
rect 113514 510854 114134 510938
rect 113514 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 114134 510854
rect 111195 487252 111261 487253
rect 111195 487188 111196 487252
rect 111260 487188 111261 487252
rect 111195 487187 111261 487188
rect 111198 483850 111258 487187
rect 113514 485308 114134 510618
rect 117234 694894 117854 708122
rect 117234 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 117854 694894
rect 117234 694574 117854 694658
rect 117234 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 117854 694574
rect 117234 658894 117854 694338
rect 117234 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 117854 658894
rect 117234 658574 117854 658658
rect 117234 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 117854 658574
rect 117234 622894 117854 658338
rect 117234 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 117854 622894
rect 117234 622574 117854 622658
rect 117234 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 117854 622574
rect 117234 586894 117854 622338
rect 117234 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 117854 586894
rect 117234 586574 117854 586658
rect 117234 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 117854 586574
rect 117234 550894 117854 586338
rect 117234 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 117854 550894
rect 117234 550574 117854 550658
rect 117234 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 117854 550574
rect 117234 514894 117854 550338
rect 117234 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 117854 514894
rect 117234 514574 117854 514658
rect 117234 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 117854 514574
rect 116163 486436 116229 486437
rect 116163 486372 116164 486436
rect 116228 486372 116229 486436
rect 116163 486371 116229 486372
rect 114323 486028 114389 486029
rect 114323 485964 114324 486028
rect 114388 485964 114389 486028
rect 114323 485963 114389 485964
rect 114326 483850 114386 485963
rect 101078 483790 101140 483850
rect 96181 483444 96247 483445
rect 96181 483380 96182 483444
rect 96246 483380 96247 483444
rect 96181 483379 96247 483380
rect 96184 483202 96244 483379
rect 98496 483202 98556 483790
rect 101080 483202 101140 483790
rect 103528 483790 103714 483850
rect 106112 483790 106290 483850
rect 108560 483790 108682 483850
rect 111144 483790 111258 483850
rect 113592 483790 114386 483850
rect 116166 483850 116226 486371
rect 117234 485308 117854 514338
rect 120954 698614 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 120954 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 121574 698614
rect 120954 698294 121574 698378
rect 120954 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 121574 698294
rect 120954 662614 121574 698058
rect 120954 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 121574 662614
rect 120954 662294 121574 662378
rect 120954 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 121574 662294
rect 120954 626614 121574 662058
rect 120954 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 121574 626614
rect 120954 626294 121574 626378
rect 120954 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 121574 626294
rect 120954 590614 121574 626058
rect 120954 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 121574 590614
rect 120954 590294 121574 590378
rect 120954 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 121574 590294
rect 120954 554614 121574 590058
rect 120954 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 121574 554614
rect 120954 554294 121574 554378
rect 120954 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 121574 554294
rect 120954 518614 121574 554058
rect 120954 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 121574 518614
rect 120954 518294 121574 518378
rect 120954 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 121574 518294
rect 118555 486300 118621 486301
rect 118555 486236 118556 486300
rect 118620 486236 118621 486300
rect 118555 486235 118621 486236
rect 118558 483850 118618 486235
rect 120954 485308 121574 518058
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 669454 128414 705242
rect 127794 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 128414 669454
rect 127794 669134 128414 669218
rect 127794 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 128414 669134
rect 127794 633454 128414 668898
rect 127794 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 128414 633454
rect 127794 633134 128414 633218
rect 127794 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 128414 633134
rect 127794 597454 128414 632898
rect 127794 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 128414 597454
rect 127794 597134 128414 597218
rect 127794 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 128414 597134
rect 127794 561454 128414 596898
rect 127794 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 128414 561454
rect 127794 561134 128414 561218
rect 127794 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 128414 561134
rect 127794 525454 128414 560898
rect 127794 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 128414 525454
rect 127794 525134 128414 525218
rect 127794 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 128414 525134
rect 127794 489454 128414 524898
rect 127794 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 128414 489454
rect 127794 489134 128414 489218
rect 127794 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 128414 489134
rect 126099 486708 126165 486709
rect 126099 486644 126100 486708
rect 126164 486644 126165 486708
rect 126099 486643 126165 486644
rect 123707 486572 123773 486573
rect 123707 486508 123708 486572
rect 123772 486508 123773 486572
rect 123707 486507 123773 486508
rect 120947 485076 121013 485077
rect 120947 485012 120948 485076
rect 121012 485012 121013 485076
rect 120947 485011 121013 485012
rect 120950 483850 121010 485011
rect 123710 483850 123770 486507
rect 116166 483790 116236 483850
rect 103528 483202 103588 483790
rect 106112 483202 106172 483790
rect 108560 483202 108620 483790
rect 111144 483202 111204 483790
rect 113592 483202 113652 483790
rect 116176 483202 116236 483790
rect 118488 483790 118618 483850
rect 120936 483790 121010 483850
rect 123656 483790 123770 483850
rect 126102 483850 126162 486643
rect 127794 485308 128414 488898
rect 131514 673174 132134 707162
rect 131514 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 132134 673174
rect 131514 672854 132134 672938
rect 131514 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 132134 672854
rect 131514 637174 132134 672618
rect 131514 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 132134 637174
rect 131514 636854 132134 636938
rect 131514 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 132134 636854
rect 131514 601174 132134 636618
rect 131514 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 132134 601174
rect 131514 600854 132134 600938
rect 131514 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 132134 600854
rect 131514 565174 132134 600618
rect 131514 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 132134 565174
rect 131514 564854 132134 564938
rect 131514 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 132134 564854
rect 131514 529174 132134 564618
rect 131514 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 132134 529174
rect 131514 528854 132134 528938
rect 131514 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 132134 528854
rect 131514 493174 132134 528618
rect 131514 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 132134 493174
rect 131514 492854 132134 492938
rect 131514 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 132134 492854
rect 130883 486708 130949 486709
rect 130883 486644 130884 486708
rect 130948 486644 130949 486708
rect 130883 486643 130949 486644
rect 128491 485212 128557 485213
rect 128491 485148 128492 485212
rect 128556 485148 128557 485212
rect 128491 485147 128557 485148
rect 128494 483850 128554 485147
rect 130886 483850 130946 486643
rect 131514 485308 132134 492618
rect 135234 676894 135854 709082
rect 135234 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 135854 676894
rect 135234 676574 135854 676658
rect 135234 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 135854 676574
rect 135234 640894 135854 676338
rect 135234 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 135854 640894
rect 135234 640574 135854 640658
rect 135234 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 135854 640574
rect 135234 604894 135854 640338
rect 135234 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 135854 604894
rect 135234 604574 135854 604658
rect 135234 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 135854 604574
rect 135234 568894 135854 604338
rect 135234 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 135854 568894
rect 135234 568574 135854 568658
rect 135234 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 135854 568574
rect 135234 532894 135854 568338
rect 135234 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 135854 532894
rect 135234 532574 135854 532658
rect 135234 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 135854 532574
rect 135234 496894 135854 532338
rect 135234 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 135854 496894
rect 135234 496574 135854 496658
rect 135234 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 135854 496574
rect 135234 485308 135854 496338
rect 138954 680614 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 138954 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 139574 680614
rect 138954 680294 139574 680378
rect 138954 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 139574 680294
rect 138954 644614 139574 680058
rect 138954 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 139574 644614
rect 138954 644294 139574 644378
rect 138954 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 139574 644294
rect 138954 608614 139574 644058
rect 138954 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 139574 608614
rect 138954 608294 139574 608378
rect 138954 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 139574 608294
rect 138954 572614 139574 608058
rect 138954 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 139574 572614
rect 138954 572294 139574 572378
rect 138954 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 139574 572294
rect 138954 536614 139574 572058
rect 138954 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 139574 536614
rect 138954 536294 139574 536378
rect 138954 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 139574 536294
rect 138954 500614 139574 536058
rect 138954 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 139574 500614
rect 138954 500294 139574 500378
rect 138954 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 139574 500294
rect 138611 486980 138677 486981
rect 138611 486916 138612 486980
rect 138676 486916 138677 486980
rect 138611 486915 138677 486916
rect 136035 485348 136101 485349
rect 136035 485284 136036 485348
rect 136100 485284 136101 485348
rect 136035 485283 136101 485284
rect 133643 483852 133709 483853
rect 133643 483850 133644 483852
rect 126102 483790 126164 483850
rect 128494 483790 128612 483850
rect 130886 483790 131060 483850
rect 118488 483202 118548 483790
rect 120936 483202 120996 483790
rect 123656 483202 123716 483790
rect 126104 483202 126164 483790
rect 128552 483202 128612 483790
rect 131000 483202 131060 483790
rect 133584 483788 133644 483850
rect 133708 483788 133709 483852
rect 136038 483850 136098 485283
rect 133584 483787 133709 483788
rect 135896 483790 136098 483850
rect 138614 483850 138674 486915
rect 138954 485308 139574 500058
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 687454 146414 704282
rect 145794 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 146414 687454
rect 145794 687134 146414 687218
rect 145794 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 146414 687134
rect 145794 651454 146414 686898
rect 145794 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 146414 651454
rect 145794 651134 146414 651218
rect 145794 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 146414 651134
rect 145794 615454 146414 650898
rect 145794 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 146414 615454
rect 145794 615134 146414 615218
rect 145794 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 146414 615134
rect 145794 579454 146414 614898
rect 145794 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 146414 579454
rect 145794 579134 146414 579218
rect 145794 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 146414 579134
rect 145794 543454 146414 578898
rect 145794 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 146414 543454
rect 145794 543134 146414 543218
rect 145794 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 146414 543134
rect 145794 507454 146414 542898
rect 145794 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 146414 507454
rect 145794 507134 146414 507218
rect 145794 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 146414 507134
rect 145603 487524 145669 487525
rect 145603 487460 145604 487524
rect 145668 487460 145669 487524
rect 145603 487459 145669 487460
rect 143579 486708 143645 486709
rect 143579 486644 143580 486708
rect 143644 486644 143645 486708
rect 143579 486643 143645 486644
rect 143582 483850 143642 486643
rect 138614 483790 138676 483850
rect 133584 483202 133644 483787
rect 135896 483202 135956 483790
rect 138616 483202 138676 483790
rect 143512 483790 143642 483850
rect 145606 483850 145666 487459
rect 145794 485308 146414 506898
rect 149514 691174 150134 706202
rect 149514 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 150134 691174
rect 149514 690854 150134 690938
rect 149514 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 150134 690854
rect 149514 655174 150134 690618
rect 149514 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 150134 655174
rect 149514 654854 150134 654938
rect 149514 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 150134 654854
rect 149514 619174 150134 654618
rect 149514 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 150134 619174
rect 149514 618854 150134 618938
rect 149514 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 150134 618854
rect 149514 583174 150134 618618
rect 149514 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 150134 583174
rect 149514 582854 150134 582938
rect 149514 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 150134 582854
rect 149514 547174 150134 582618
rect 149514 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 150134 547174
rect 149514 546854 150134 546938
rect 149514 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 150134 546854
rect 149514 511174 150134 546618
rect 149514 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 150134 511174
rect 149514 510854 150134 510938
rect 149514 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 150134 510854
rect 149514 485308 150134 510618
rect 153234 694894 153854 708122
rect 153234 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 153854 694894
rect 153234 694574 153854 694658
rect 153234 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 153854 694574
rect 153234 658894 153854 694338
rect 153234 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 153854 658894
rect 153234 658574 153854 658658
rect 153234 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 153854 658574
rect 153234 622894 153854 658338
rect 153234 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 153854 622894
rect 153234 622574 153854 622658
rect 153234 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 153854 622574
rect 153234 586894 153854 622338
rect 153234 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 153854 586894
rect 153234 586574 153854 586658
rect 153234 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 153854 586574
rect 153234 550894 153854 586338
rect 153234 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 153854 550894
rect 153234 550574 153854 550658
rect 153234 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 153854 550574
rect 153234 514894 153854 550338
rect 153234 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 153854 514894
rect 153234 514574 153854 514658
rect 153234 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 153854 514574
rect 150939 486844 151005 486845
rect 150939 486780 150940 486844
rect 151004 486780 151005 486844
rect 150939 486779 151005 486780
rect 150942 483850 151002 486779
rect 153234 485308 153854 514338
rect 156954 698614 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 156954 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 157574 698614
rect 156954 698294 157574 698378
rect 156954 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 157574 698294
rect 156954 662614 157574 698058
rect 156954 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 157574 662614
rect 156954 662294 157574 662378
rect 156954 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 157574 662294
rect 156954 626614 157574 662058
rect 156954 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 157574 626614
rect 156954 626294 157574 626378
rect 156954 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 157574 626294
rect 156954 590614 157574 626058
rect 156954 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 157574 590614
rect 156954 590294 157574 590378
rect 156954 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 157574 590294
rect 156954 554614 157574 590058
rect 156954 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 157574 554614
rect 156954 554294 157574 554378
rect 156954 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 157574 554294
rect 156954 518614 157574 554058
rect 156954 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 157574 518614
rect 156954 518294 157574 518378
rect 156954 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 157574 518294
rect 156954 485308 157574 518058
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 669454 164414 705242
rect 163794 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 164414 669454
rect 163794 669134 164414 669218
rect 163794 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 164414 669134
rect 163794 633454 164414 668898
rect 163794 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 164414 633454
rect 163794 633134 164414 633218
rect 163794 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 164414 633134
rect 163794 597454 164414 632898
rect 163794 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 164414 597454
rect 163794 597134 164414 597218
rect 163794 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 164414 597134
rect 163794 561454 164414 596898
rect 163794 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 164414 561454
rect 163794 561134 164414 561218
rect 163794 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 164414 561134
rect 163794 525454 164414 560898
rect 163794 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 164414 525454
rect 163794 525134 164414 525218
rect 163794 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 164414 525134
rect 163794 489454 164414 524898
rect 163794 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 164414 489454
rect 163794 489134 164414 489218
rect 163794 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 164414 489134
rect 158483 485892 158549 485893
rect 158483 485828 158484 485892
rect 158548 485828 158549 485892
rect 158483 485827 158549 485828
rect 155907 484260 155973 484261
rect 155907 484196 155908 484260
rect 155972 484196 155973 484260
rect 155907 484195 155973 484196
rect 155910 483850 155970 484195
rect 158486 483850 158546 485827
rect 163794 485308 164414 488898
rect 167514 673174 168134 707162
rect 167514 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 168134 673174
rect 167514 672854 168134 672938
rect 167514 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 168134 672854
rect 167514 637174 168134 672618
rect 167514 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 168134 637174
rect 167514 636854 168134 636938
rect 167514 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 168134 636854
rect 167514 601174 168134 636618
rect 167514 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 168134 601174
rect 167514 600854 168134 600938
rect 167514 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 168134 600854
rect 167514 565174 168134 600618
rect 167514 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 168134 565174
rect 167514 564854 168134 564938
rect 167514 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 168134 564854
rect 167514 529174 168134 564618
rect 167514 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 168134 529174
rect 167514 528854 168134 528938
rect 167514 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 168134 528854
rect 167514 493174 168134 528618
rect 167514 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 168134 493174
rect 167514 492854 168134 492938
rect 167514 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 168134 492854
rect 166027 485756 166093 485757
rect 166027 485692 166028 485756
rect 166092 485692 166093 485756
rect 166027 485691 166093 485692
rect 161059 484124 161125 484125
rect 161059 484060 161060 484124
rect 161124 484060 161125 484124
rect 161059 484059 161125 484060
rect 161062 483850 161122 484059
rect 163267 483988 163333 483989
rect 163267 483924 163268 483988
rect 163332 483924 163333 483988
rect 163267 483923 163333 483924
rect 145606 483790 146020 483850
rect 150942 483790 151052 483850
rect 155910 483790 156084 483850
rect 141061 483444 141127 483445
rect 141061 483380 141062 483444
rect 141126 483380 141127 483444
rect 141061 483379 141127 483380
rect 141064 483202 141124 483379
rect 143512 483202 143572 483790
rect 145960 483202 146020 483790
rect 148405 483580 148471 483581
rect 148405 483516 148406 483580
rect 148470 483516 148471 483580
rect 148405 483515 148471 483516
rect 148408 483202 148468 483515
rect 150992 483202 151052 483790
rect 153573 483716 153639 483717
rect 153573 483652 153574 483716
rect 153638 483652 153639 483716
rect 153573 483651 153639 483652
rect 153576 483202 153636 483651
rect 156024 483202 156084 483790
rect 158472 483790 158546 483850
rect 161056 483790 161122 483850
rect 163270 483850 163330 483923
rect 166030 483850 166090 485691
rect 167514 485308 168134 492618
rect 171234 676894 171854 709082
rect 171234 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 171854 676894
rect 171234 676574 171854 676658
rect 171234 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 171854 676574
rect 171234 640894 171854 676338
rect 171234 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 171854 640894
rect 171234 640574 171854 640658
rect 171234 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 171854 640574
rect 171234 604894 171854 640338
rect 171234 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 171854 604894
rect 171234 604574 171854 604658
rect 171234 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 171854 604574
rect 171234 568894 171854 604338
rect 171234 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 171854 568894
rect 171234 568574 171854 568658
rect 171234 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 171854 568574
rect 171234 532894 171854 568338
rect 171234 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 171854 532894
rect 171234 532574 171854 532658
rect 171234 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 171854 532574
rect 171234 496894 171854 532338
rect 171234 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 171854 496894
rect 171234 496574 171854 496658
rect 171234 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 171854 496574
rect 171234 485308 171854 496338
rect 174954 680614 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 174954 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 175574 680614
rect 174954 680294 175574 680378
rect 174954 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 175574 680294
rect 174954 644614 175574 680058
rect 174954 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 175574 644614
rect 174954 644294 175574 644378
rect 174954 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 175574 644294
rect 174954 608614 175574 644058
rect 174954 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 175574 608614
rect 174954 608294 175574 608378
rect 174954 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 175574 608294
rect 174954 572614 175574 608058
rect 174954 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 175574 572614
rect 174954 572294 175574 572378
rect 174954 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 175574 572294
rect 174954 536614 175574 572058
rect 174954 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 175574 536614
rect 174954 536294 175574 536378
rect 174954 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 175574 536294
rect 174954 500614 175574 536058
rect 174954 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 175574 500614
rect 174954 500294 175574 500378
rect 174954 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 175574 500294
rect 174954 485308 175574 500058
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 687454 182414 704282
rect 181794 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 182414 687454
rect 181794 687134 182414 687218
rect 181794 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 182414 687134
rect 181794 651454 182414 686898
rect 181794 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 182414 651454
rect 181794 651134 182414 651218
rect 181794 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 182414 651134
rect 181794 615454 182414 650898
rect 181794 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 182414 615454
rect 181794 615134 182414 615218
rect 181794 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 182414 615134
rect 181794 579454 182414 614898
rect 181794 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 182414 579454
rect 181794 579134 182414 579218
rect 181794 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 182414 579134
rect 181794 543454 182414 578898
rect 181794 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 182414 543454
rect 181794 543134 182414 543218
rect 181794 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 182414 543134
rect 181794 507454 182414 542898
rect 181794 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 182414 507454
rect 181794 507134 182414 507218
rect 181794 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 182414 507134
rect 178355 485620 178421 485621
rect 178355 485556 178356 485620
rect 178420 485556 178421 485620
rect 178355 485555 178421 485556
rect 178358 483850 178418 485555
rect 181794 485308 182414 506898
rect 185514 691174 186134 706202
rect 185514 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 186134 691174
rect 185514 690854 186134 690938
rect 185514 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 186134 690854
rect 185514 655174 186134 690618
rect 185514 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 186134 655174
rect 185514 654854 186134 654938
rect 185514 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 186134 654854
rect 185514 619174 186134 654618
rect 185514 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 186134 619174
rect 185514 618854 186134 618938
rect 185514 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 186134 618854
rect 185514 583174 186134 618618
rect 185514 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 186134 583174
rect 185514 582854 186134 582938
rect 185514 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 186134 582854
rect 185514 547174 186134 582618
rect 185514 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 186134 547174
rect 185514 546854 186134 546938
rect 185514 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 186134 546854
rect 185514 511174 186134 546618
rect 185514 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 186134 511174
rect 185514 510854 186134 510938
rect 185514 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 186134 510854
rect 185514 485308 186134 510618
rect 189234 694894 189854 708122
rect 189234 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 189854 694894
rect 189234 694574 189854 694658
rect 189234 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 189854 694574
rect 189234 658894 189854 694338
rect 189234 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 189854 658894
rect 189234 658574 189854 658658
rect 189234 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 189854 658574
rect 189234 622894 189854 658338
rect 189234 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 189854 622894
rect 189234 622574 189854 622658
rect 189234 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 189854 622574
rect 189234 586894 189854 622338
rect 189234 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 189854 586894
rect 189234 586574 189854 586658
rect 189234 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 189854 586574
rect 189234 550894 189854 586338
rect 189234 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 189854 550894
rect 189234 550574 189854 550658
rect 189234 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 189854 550574
rect 189234 514894 189854 550338
rect 189234 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 189854 514894
rect 189234 514574 189854 514658
rect 189234 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 189854 514574
rect 189234 485308 189854 514338
rect 192954 698614 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 192954 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 193574 698614
rect 192954 698294 193574 698378
rect 192954 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 193574 698294
rect 192954 662614 193574 698058
rect 192954 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 193574 662614
rect 192954 662294 193574 662378
rect 192954 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 193574 662294
rect 192954 626614 193574 662058
rect 192954 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 193574 626614
rect 192954 626294 193574 626378
rect 192954 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 193574 626294
rect 192954 590614 193574 626058
rect 192954 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 193574 590614
rect 192954 590294 193574 590378
rect 192954 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 193574 590294
rect 192954 554614 193574 590058
rect 192954 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 193574 554614
rect 192954 554294 193574 554378
rect 192954 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 193574 554294
rect 192954 518614 193574 554058
rect 192954 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 193574 518614
rect 192954 518294 193574 518378
rect 192954 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 193574 518294
rect 192954 485308 193574 518058
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 669454 200414 705242
rect 199794 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 200414 669454
rect 199794 669134 200414 669218
rect 199794 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 200414 669134
rect 199794 633454 200414 668898
rect 199794 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 200414 633454
rect 199794 633134 200414 633218
rect 199794 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 200414 633134
rect 199794 597454 200414 632898
rect 199794 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 200414 597454
rect 199794 597134 200414 597218
rect 199794 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 200414 597134
rect 199794 561454 200414 596898
rect 199794 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 200414 561454
rect 199794 561134 200414 561218
rect 199794 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 200414 561134
rect 199794 525454 200414 560898
rect 199794 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 200414 525454
rect 199794 525134 200414 525218
rect 199794 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 200414 525134
rect 199794 489454 200414 524898
rect 199794 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 200414 489454
rect 199794 489134 200414 489218
rect 199794 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 200414 489134
rect 179643 484532 179709 484533
rect 179643 484468 179644 484532
rect 179708 484468 179709 484532
rect 179643 484467 179709 484468
rect 190867 484532 190933 484533
rect 190867 484468 190868 484532
rect 190932 484468 190933 484532
rect 190867 484467 190933 484468
rect 179646 483850 179706 484467
rect 190870 483850 190930 484467
rect 163270 483790 163428 483850
rect 166030 483790 166148 483850
rect 178358 483790 178524 483850
rect 179646 483790 179748 483850
rect 158472 483202 158532 483790
rect 161056 483202 161116 483790
rect 163368 483202 163428 483790
rect 166088 483202 166148 483790
rect 178464 483202 178524 483790
rect 179688 483202 179748 483790
rect 190840 483790 190930 483850
rect 190840 483202 190900 483790
rect 60952 471454 61300 471486
rect 60952 471218 61008 471454
rect 61244 471218 61300 471454
rect 60952 471134 61300 471218
rect 60952 470898 61008 471134
rect 61244 470898 61300 471134
rect 60952 470866 61300 470898
rect 195320 471454 195668 471486
rect 195320 471218 195376 471454
rect 195612 471218 195668 471454
rect 195320 471134 195668 471218
rect 195320 470898 195376 471134
rect 195612 470898 195668 471134
rect 195320 470866 195668 470898
rect 55794 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 56414 453454
rect 55794 453134 56414 453218
rect 55794 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 56414 453134
rect 55794 417454 56414 452898
rect 60272 453454 60620 453486
rect 60272 453218 60328 453454
rect 60564 453218 60620 453454
rect 60272 453134 60620 453218
rect 60272 452898 60328 453134
rect 60564 452898 60620 453134
rect 60272 452866 60620 452898
rect 196000 453454 196348 453486
rect 196000 453218 196056 453454
rect 196292 453218 196348 453454
rect 196000 453134 196348 453218
rect 196000 452898 196056 453134
rect 196292 452898 196348 453134
rect 196000 452866 196348 452898
rect 199794 453454 200414 488898
rect 199794 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 200414 453454
rect 199794 453134 200414 453218
rect 199794 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 200414 453134
rect 60952 435454 61300 435486
rect 60952 435218 61008 435454
rect 61244 435218 61300 435454
rect 60952 435134 61300 435218
rect 60952 434898 61008 435134
rect 61244 434898 61300 435134
rect 60952 434866 61300 434898
rect 195320 435454 195668 435486
rect 195320 435218 195376 435454
rect 195612 435218 195668 435454
rect 195320 435134 195668 435218
rect 195320 434898 195376 435134
rect 195612 434898 195668 435134
rect 195320 434866 195668 434898
rect 55794 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 56414 417454
rect 55794 417134 56414 417218
rect 55794 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 56414 417134
rect 55794 381454 56414 416898
rect 60272 417454 60620 417486
rect 60272 417218 60328 417454
rect 60564 417218 60620 417454
rect 60272 417134 60620 417218
rect 60272 416898 60328 417134
rect 60564 416898 60620 417134
rect 60272 416866 60620 416898
rect 196000 417454 196348 417486
rect 196000 417218 196056 417454
rect 196292 417218 196348 417454
rect 196000 417134 196348 417218
rect 196000 416898 196056 417134
rect 196292 416898 196348 417134
rect 196000 416866 196348 416898
rect 199794 417454 200414 452898
rect 199794 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 200414 417454
rect 199794 417134 200414 417218
rect 199794 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 200414 417134
rect 76056 399530 76116 400106
rect 76054 399470 76116 399530
rect 77144 399530 77204 400106
rect 78232 399530 78292 400106
rect 79592 399530 79652 400106
rect 80544 399530 80604 400106
rect 77144 399470 77218 399530
rect 78232 399470 78322 399530
rect 55794 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 56414 381454
rect 55794 381134 56414 381218
rect 55794 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 56414 381134
rect 55794 345454 56414 380898
rect 55794 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 56414 345454
rect 55794 345134 56414 345218
rect 55794 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 56414 345134
rect 55794 309454 56414 344898
rect 55794 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 56414 309454
rect 55794 309134 56414 309218
rect 55794 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 56414 309134
rect 55794 273454 56414 308898
rect 55794 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 56414 273454
rect 55794 273134 56414 273218
rect 55794 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 56414 273134
rect 55794 237454 56414 272898
rect 55794 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 56414 237454
rect 55794 237134 56414 237218
rect 55794 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 56414 237134
rect 55794 201454 56414 236898
rect 59514 385174 60134 398000
rect 59514 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 60134 385174
rect 59514 384854 60134 384938
rect 59514 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 60134 384854
rect 59514 349174 60134 384618
rect 59514 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 60134 349174
rect 59514 348854 60134 348938
rect 59514 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 60134 348854
rect 59514 313174 60134 348618
rect 59514 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 60134 313174
rect 59514 312854 60134 312938
rect 59514 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 60134 312854
rect 59514 277174 60134 312618
rect 59514 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 60134 277174
rect 59514 276854 60134 276938
rect 59514 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 60134 276854
rect 59514 241174 60134 276618
rect 59514 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 60134 241174
rect 59514 240854 60134 240938
rect 59514 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 60134 240854
rect 59514 228924 60134 240618
rect 63234 388894 63854 398000
rect 63234 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 63854 388894
rect 63234 388574 63854 388658
rect 63234 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 63854 388574
rect 63234 352894 63854 388338
rect 63234 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 63854 352894
rect 63234 352574 63854 352658
rect 63234 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 63854 352574
rect 63234 316894 63854 352338
rect 63234 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 63854 316894
rect 63234 316574 63854 316658
rect 63234 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 63854 316574
rect 63234 280894 63854 316338
rect 63234 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 63854 280894
rect 63234 280574 63854 280658
rect 63234 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 63854 280574
rect 63234 244894 63854 280338
rect 63234 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 63854 244894
rect 63234 244574 63854 244658
rect 63234 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 63854 244574
rect 63234 228924 63854 244338
rect 66954 392614 67574 398000
rect 66954 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 67574 392614
rect 66954 392294 67574 392378
rect 66954 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 67574 392294
rect 66954 356614 67574 392058
rect 66954 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 67574 356614
rect 66954 356294 67574 356378
rect 66954 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 67574 356294
rect 66954 320614 67574 356058
rect 66954 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 67574 320614
rect 66954 320294 67574 320378
rect 66954 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 67574 320294
rect 66954 284614 67574 320058
rect 66954 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 67574 284614
rect 66954 284294 67574 284378
rect 66954 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 67574 284294
rect 66954 248614 67574 284058
rect 66954 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 67574 248614
rect 66954 248294 67574 248378
rect 66954 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 67574 248294
rect 66954 228924 67574 248058
rect 73794 363454 74414 398000
rect 76054 396813 76114 399470
rect 76051 396812 76117 396813
rect 76051 396748 76052 396812
rect 76116 396748 76117 396812
rect 76051 396747 76117 396748
rect 77158 396677 77218 399470
rect 77155 396676 77221 396677
rect 77155 396612 77156 396676
rect 77220 396612 77221 396676
rect 77155 396611 77221 396612
rect 73794 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 74414 363454
rect 73794 363134 74414 363218
rect 73794 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 74414 363134
rect 73794 327454 74414 362898
rect 73794 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 74414 327454
rect 73794 327134 74414 327218
rect 73794 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 74414 327134
rect 73794 291454 74414 326898
rect 73794 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 74414 291454
rect 73794 291134 74414 291218
rect 73794 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 74414 291134
rect 73794 255454 74414 290898
rect 73794 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 74414 255454
rect 73794 255134 74414 255218
rect 73794 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 74414 255134
rect 73794 228924 74414 254898
rect 77514 367174 78134 398000
rect 78262 397357 78322 399470
rect 79550 399470 79652 399530
rect 80470 399470 80604 399530
rect 81768 399530 81828 400106
rect 83128 399530 83188 400106
rect 84216 399530 84276 400106
rect 85440 399530 85500 400106
rect 81768 399470 82002 399530
rect 83128 399470 83290 399530
rect 84216 399470 84394 399530
rect 79550 397357 79610 399470
rect 80470 397357 80530 399470
rect 78259 397356 78325 397357
rect 78259 397292 78260 397356
rect 78324 397292 78325 397356
rect 78259 397291 78325 397292
rect 79547 397356 79613 397357
rect 79547 397292 79548 397356
rect 79612 397292 79613 397356
rect 79547 397291 79613 397292
rect 80467 397356 80533 397357
rect 80467 397292 80468 397356
rect 80532 397292 80533 397356
rect 80467 397291 80533 397292
rect 77514 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 78134 367174
rect 77514 366854 78134 366938
rect 77514 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 78134 366854
rect 77514 331174 78134 366618
rect 77514 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 78134 331174
rect 77514 330854 78134 330938
rect 77514 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 78134 330854
rect 77514 295174 78134 330618
rect 77514 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 78134 295174
rect 77514 294854 78134 294938
rect 77514 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 78134 294854
rect 77514 259174 78134 294618
rect 77514 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 78134 259174
rect 77514 258854 78134 258938
rect 77514 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 78134 258854
rect 77514 228924 78134 258618
rect 81234 370894 81854 398000
rect 81942 396813 82002 399470
rect 83230 397357 83290 399470
rect 83227 397356 83293 397357
rect 83227 397292 83228 397356
rect 83292 397292 83293 397356
rect 83227 397291 83293 397292
rect 84334 396813 84394 399470
rect 85438 399470 85500 399530
rect 86528 399530 86588 400106
rect 87616 399530 87676 400106
rect 88296 399530 88356 400106
rect 88704 399530 88764 400106
rect 90064 399530 90124 400106
rect 86528 399470 86602 399530
rect 87616 399470 87706 399530
rect 88296 399470 88442 399530
rect 88704 399470 88810 399530
rect 85438 398173 85498 399470
rect 85435 398172 85501 398173
rect 85435 398108 85436 398172
rect 85500 398108 85501 398172
rect 85435 398107 85501 398108
rect 81939 396812 82005 396813
rect 81939 396748 81940 396812
rect 82004 396748 82005 396812
rect 81939 396747 82005 396748
rect 84331 396812 84397 396813
rect 84331 396748 84332 396812
rect 84396 396748 84397 396812
rect 84331 396747 84397 396748
rect 81234 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 81854 370894
rect 81234 370574 81854 370658
rect 81234 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 81854 370574
rect 81234 334894 81854 370338
rect 81234 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 81854 334894
rect 81234 334574 81854 334658
rect 81234 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 81854 334574
rect 81234 298894 81854 334338
rect 81234 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 81854 298894
rect 81234 298574 81854 298658
rect 81234 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 81854 298574
rect 81234 262894 81854 298338
rect 81234 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 81854 262894
rect 81234 262574 81854 262658
rect 81234 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 81854 262574
rect 81234 228924 81854 262338
rect 84954 374614 85574 398000
rect 86542 397357 86602 399470
rect 87646 397357 87706 399470
rect 86539 397356 86605 397357
rect 86539 397292 86540 397356
rect 86604 397292 86605 397356
rect 86539 397291 86605 397292
rect 87643 397356 87709 397357
rect 87643 397292 87644 397356
rect 87708 397292 87709 397356
rect 87643 397291 87709 397292
rect 88382 396813 88442 399470
rect 88750 397357 88810 399470
rect 90038 399470 90124 399530
rect 90744 399530 90804 400106
rect 91288 399530 91348 400106
rect 92376 399530 92436 400106
rect 93464 399530 93524 400106
rect 90744 399470 90834 399530
rect 91288 399470 91386 399530
rect 88747 397356 88813 397357
rect 88747 397292 88748 397356
rect 88812 397292 88813 397356
rect 88747 397291 88813 397292
rect 90038 396813 90098 399470
rect 88379 396812 88445 396813
rect 88379 396748 88380 396812
rect 88444 396748 88445 396812
rect 88379 396747 88445 396748
rect 90035 396812 90101 396813
rect 90035 396748 90036 396812
rect 90100 396748 90101 396812
rect 90035 396747 90101 396748
rect 90774 396677 90834 399470
rect 91326 397357 91386 399470
rect 91510 399470 92436 399530
rect 93350 399470 93524 399530
rect 93600 399530 93660 400106
rect 94552 399530 94612 400106
rect 95912 399530 95972 400106
rect 96048 399669 96108 400106
rect 96045 399668 96111 399669
rect 96045 399604 96046 399668
rect 96110 399604 96111 399668
rect 96045 399603 96111 399604
rect 96475 399668 96541 399669
rect 96475 399604 96476 399668
rect 96540 399604 96541 399668
rect 96475 399603 96541 399604
rect 93600 399470 93778 399530
rect 94552 399470 94698 399530
rect 95912 399470 96354 399530
rect 91323 397356 91389 397357
rect 91323 397292 91324 397356
rect 91388 397292 91389 397356
rect 91323 397291 91389 397292
rect 91510 396677 91570 399470
rect 90771 396676 90837 396677
rect 90771 396612 90772 396676
rect 90836 396612 90837 396676
rect 90771 396611 90837 396612
rect 91507 396676 91573 396677
rect 91507 396612 91508 396676
rect 91572 396612 91573 396676
rect 91507 396611 91573 396612
rect 84954 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 85574 374614
rect 84954 374294 85574 374378
rect 84954 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 85574 374294
rect 84954 338614 85574 374058
rect 84954 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 85574 338614
rect 84954 338294 85574 338378
rect 84954 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 85574 338294
rect 84954 302614 85574 338058
rect 84954 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 85574 302614
rect 84954 302294 85574 302378
rect 84954 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 85574 302294
rect 84954 266614 85574 302058
rect 84954 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 85574 266614
rect 84954 266294 85574 266378
rect 84954 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 85574 266294
rect 84954 230614 85574 266058
rect 84954 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 85574 230614
rect 84954 230294 85574 230378
rect 84954 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 85574 230294
rect 84954 228924 85574 230058
rect 91794 381454 92414 398000
rect 93350 397357 93410 399470
rect 93347 397356 93413 397357
rect 93347 397292 93348 397356
rect 93412 397292 93413 397356
rect 93347 397291 93413 397292
rect 93718 396813 93778 399470
rect 94638 396813 94698 399470
rect 93715 396812 93781 396813
rect 93715 396748 93716 396812
rect 93780 396748 93781 396812
rect 93715 396747 93781 396748
rect 94635 396812 94701 396813
rect 94635 396748 94636 396812
rect 94700 396748 94701 396812
rect 94635 396747 94701 396748
rect 91794 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 92414 381454
rect 91794 381134 92414 381218
rect 91794 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 92414 381134
rect 91794 345454 92414 380898
rect 91794 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 92414 345454
rect 91794 345134 92414 345218
rect 91794 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 92414 345134
rect 91794 309454 92414 344898
rect 91794 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 92414 309454
rect 91794 309134 92414 309218
rect 91794 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 92414 309134
rect 91794 273454 92414 308898
rect 91794 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 92414 273454
rect 91794 273134 92414 273218
rect 91794 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 92414 273134
rect 91794 237454 92414 272898
rect 91794 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 92414 237454
rect 91794 237134 92414 237218
rect 91794 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 92414 237134
rect 91794 228924 92414 236898
rect 95514 385174 96134 398000
rect 96294 397357 96354 399470
rect 96291 397356 96357 397357
rect 96291 397292 96292 397356
rect 96356 397292 96357 397356
rect 96291 397291 96357 397292
rect 96478 397221 96538 399603
rect 97000 399530 97060 400106
rect 98088 399530 98148 400106
rect 98496 399530 98556 400106
rect 99448 399530 99508 400106
rect 100672 399530 100732 400106
rect 101080 399530 101140 400106
rect 97000 399470 97090 399530
rect 98088 399470 98194 399530
rect 98496 399470 98562 399530
rect 99448 399470 100034 399530
rect 100672 399470 100770 399530
rect 96475 397220 96541 397221
rect 96475 397156 96476 397220
rect 96540 397156 96541 397220
rect 96475 397155 96541 397156
rect 97030 396813 97090 399470
rect 98134 397357 98194 399470
rect 98131 397356 98197 397357
rect 98131 397292 98132 397356
rect 98196 397292 98197 397356
rect 98131 397291 98197 397292
rect 98502 397221 98562 399470
rect 98499 397220 98565 397221
rect 98499 397156 98500 397220
rect 98564 397156 98565 397220
rect 98499 397155 98565 397156
rect 97027 396812 97093 396813
rect 97027 396748 97028 396812
rect 97092 396748 97093 396812
rect 97027 396747 97093 396748
rect 95514 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 96134 385174
rect 95514 384854 96134 384938
rect 95514 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 96134 384854
rect 95514 349174 96134 384618
rect 95514 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 96134 349174
rect 95514 348854 96134 348938
rect 95514 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 96134 348854
rect 95514 313174 96134 348618
rect 95514 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 96134 313174
rect 95514 312854 96134 312938
rect 95514 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 96134 312854
rect 95514 277174 96134 312618
rect 95514 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 96134 277174
rect 95514 276854 96134 276938
rect 95514 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 96134 276854
rect 95514 241174 96134 276618
rect 95514 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 96134 241174
rect 95514 240854 96134 240938
rect 95514 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 96134 240854
rect 95514 228924 96134 240618
rect 99234 388894 99854 398000
rect 99974 397357 100034 399470
rect 100710 397357 100770 399470
rect 101078 399470 101140 399530
rect 101760 399530 101820 400106
rect 102848 399530 102908 400106
rect 101760 399470 101874 399530
rect 99971 397356 100037 397357
rect 99971 397292 99972 397356
rect 100036 397292 100037 397356
rect 99971 397291 100037 397292
rect 100707 397356 100773 397357
rect 100707 397292 100708 397356
rect 100772 397292 100773 397356
rect 100707 397291 100773 397292
rect 101078 396813 101138 399470
rect 101814 397357 101874 399470
rect 102734 399470 102908 399530
rect 103528 399530 103588 400106
rect 103936 399530 103996 400106
rect 103528 399470 103714 399530
rect 102734 397357 102794 399470
rect 101811 397356 101877 397357
rect 101811 397292 101812 397356
rect 101876 397292 101877 397356
rect 101811 397291 101877 397292
rect 102731 397356 102797 397357
rect 102731 397292 102732 397356
rect 102796 397292 102797 397356
rect 102731 397291 102797 397292
rect 101075 396812 101141 396813
rect 101075 396748 101076 396812
rect 101140 396748 101141 396812
rect 101075 396747 101141 396748
rect 99234 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 99854 388894
rect 99234 388574 99854 388658
rect 99234 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 99854 388574
rect 99234 352894 99854 388338
rect 99234 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 99854 352894
rect 99234 352574 99854 352658
rect 99234 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 99854 352574
rect 99234 316894 99854 352338
rect 99234 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 99854 316894
rect 99234 316574 99854 316658
rect 99234 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 99854 316574
rect 99234 280894 99854 316338
rect 99234 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 99854 280894
rect 99234 280574 99854 280658
rect 99234 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 99854 280574
rect 99234 244894 99854 280338
rect 99234 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 99854 244894
rect 99234 244574 99854 244658
rect 99234 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 99854 244574
rect 99234 228924 99854 244338
rect 102954 392614 103574 398000
rect 103654 397218 103714 399470
rect 103838 399470 103996 399530
rect 105296 399530 105356 400106
rect 105976 399530 106036 400106
rect 106384 399530 106444 400106
rect 107608 399530 107668 400106
rect 108288 399530 108348 400106
rect 105296 399470 105370 399530
rect 105976 399470 106106 399530
rect 106384 399470 106474 399530
rect 103838 397357 103898 399470
rect 105310 397357 105370 399470
rect 103835 397356 103901 397357
rect 103835 397292 103836 397356
rect 103900 397292 103901 397356
rect 103835 397291 103901 397292
rect 105307 397356 105373 397357
rect 105307 397292 105308 397356
rect 105372 397292 105373 397356
rect 105307 397291 105373 397292
rect 103835 397220 103901 397221
rect 103835 397218 103836 397220
rect 103654 397158 103836 397218
rect 103835 397156 103836 397158
rect 103900 397156 103901 397220
rect 103835 397155 103901 397156
rect 106046 396813 106106 399470
rect 106414 397357 106474 399470
rect 107518 399470 107668 399530
rect 108254 399470 108348 399530
rect 108696 399530 108756 400106
rect 109784 399530 109844 400106
rect 108696 399470 108866 399530
rect 106411 397356 106477 397357
rect 106411 397292 106412 397356
rect 106476 397292 106477 397356
rect 106411 397291 106477 397292
rect 107518 396813 107578 399470
rect 106043 396812 106109 396813
rect 106043 396748 106044 396812
rect 106108 396748 106109 396812
rect 106043 396747 106109 396748
rect 107515 396812 107581 396813
rect 107515 396748 107516 396812
rect 107580 396748 107581 396812
rect 107515 396747 107581 396748
rect 108254 396677 108314 399470
rect 108806 396813 108866 399470
rect 109542 399470 109844 399530
rect 111008 399530 111068 400106
rect 111144 399530 111204 400106
rect 112232 399530 112292 400106
rect 113320 399530 113380 400106
rect 111008 399470 111074 399530
rect 111144 399470 111258 399530
rect 112232 399470 112362 399530
rect 109542 397357 109602 399470
rect 109539 397356 109605 397357
rect 109539 397292 109540 397356
rect 109604 397292 109605 397356
rect 109539 397291 109605 397292
rect 108803 396812 108869 396813
rect 108803 396748 108804 396812
rect 108868 396748 108869 396812
rect 108803 396747 108869 396748
rect 108251 396676 108317 396677
rect 108251 396612 108252 396676
rect 108316 396612 108317 396676
rect 108251 396611 108317 396612
rect 102954 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 103574 392614
rect 102954 392294 103574 392378
rect 102954 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 103574 392294
rect 102954 356614 103574 392058
rect 102954 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 103574 356614
rect 102954 356294 103574 356378
rect 102954 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 103574 356294
rect 102954 320614 103574 356058
rect 102954 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 103574 320614
rect 102954 320294 103574 320378
rect 102954 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 103574 320294
rect 102954 284614 103574 320058
rect 102954 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 103574 284614
rect 102954 284294 103574 284378
rect 102954 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 103574 284294
rect 102954 248614 103574 284058
rect 102954 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 103574 248614
rect 102954 248294 103574 248378
rect 102954 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 103574 248294
rect 102954 228924 103574 248058
rect 109794 363454 110414 398000
rect 111014 396813 111074 399470
rect 111198 397357 111258 399470
rect 111195 397356 111261 397357
rect 111195 397292 111196 397356
rect 111260 397292 111261 397356
rect 111195 397291 111261 397292
rect 112302 396813 112362 399470
rect 113222 399470 113380 399530
rect 113222 397221 113282 399470
rect 113590 398173 113650 400136
rect 114408 399530 114468 400106
rect 114408 399470 114570 399530
rect 113587 398172 113653 398173
rect 113587 398108 113588 398172
rect 113652 398108 113653 398172
rect 113587 398107 113653 398108
rect 113219 397220 113285 397221
rect 113219 397156 113220 397220
rect 113284 397156 113285 397220
rect 113219 397155 113285 397156
rect 111011 396812 111077 396813
rect 111011 396748 111012 396812
rect 111076 396748 111077 396812
rect 111011 396747 111077 396748
rect 112299 396812 112365 396813
rect 112299 396748 112300 396812
rect 112364 396748 112365 396812
rect 112299 396747 112365 396748
rect 109794 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 110414 363454
rect 109794 363134 110414 363218
rect 109794 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 110414 363134
rect 109794 327454 110414 362898
rect 109794 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 110414 327454
rect 109794 327134 110414 327218
rect 109794 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 110414 327134
rect 109794 291454 110414 326898
rect 109794 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 110414 291454
rect 109794 291134 110414 291218
rect 109794 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 110414 291134
rect 109794 255454 110414 290898
rect 109794 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 110414 255454
rect 109794 255134 110414 255218
rect 109794 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 110414 255134
rect 109794 228924 110414 254898
rect 113514 367174 114134 398000
rect 114510 397357 114570 399470
rect 115798 397357 115858 400136
rect 115982 400076 116070 400136
rect 114507 397356 114573 397357
rect 114507 397292 114508 397356
rect 114572 397292 114573 397356
rect 114507 397291 114573 397292
rect 115795 397356 115861 397357
rect 115795 397292 115796 397356
rect 115860 397292 115861 397356
rect 115795 397291 115861 397292
rect 115982 396677 116042 400076
rect 116992 399530 117052 400106
rect 118080 399530 118140 400106
rect 118488 399530 118548 400106
rect 119168 399530 119228 400106
rect 120936 399530 120996 400106
rect 116992 399470 117146 399530
rect 118080 399470 118250 399530
rect 117086 396813 117146 399470
rect 117083 396812 117149 396813
rect 117083 396748 117084 396812
rect 117148 396748 117149 396812
rect 117083 396747 117149 396748
rect 115979 396676 116045 396677
rect 115979 396612 115980 396676
rect 116044 396612 116045 396676
rect 115979 396611 116045 396612
rect 113514 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 114134 367174
rect 113514 366854 114134 366938
rect 113514 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 114134 366854
rect 113514 331174 114134 366618
rect 113514 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 114134 331174
rect 113514 330854 114134 330938
rect 113514 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 114134 330854
rect 113514 295174 114134 330618
rect 113514 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 114134 295174
rect 113514 294854 114134 294938
rect 113514 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 114134 294854
rect 113514 259174 114134 294618
rect 113514 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 114134 259174
rect 113514 258854 114134 258938
rect 113514 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 114134 258854
rect 113514 228924 114134 258618
rect 117234 370894 117854 398000
rect 118190 396813 118250 399470
rect 118374 399470 118548 399530
rect 119110 399470 119228 399530
rect 120766 399470 120996 399530
rect 123520 399530 123580 400106
rect 125968 399530 126028 400106
rect 123520 399470 123586 399530
rect 118374 397357 118434 399470
rect 118371 397356 118437 397357
rect 118371 397292 118372 397356
rect 118436 397292 118437 397356
rect 118371 397291 118437 397292
rect 119110 396813 119170 399470
rect 120766 396813 120826 399470
rect 118187 396812 118253 396813
rect 118187 396748 118188 396812
rect 118252 396748 118253 396812
rect 118187 396747 118253 396748
rect 119107 396812 119173 396813
rect 119107 396748 119108 396812
rect 119172 396748 119173 396812
rect 119107 396747 119173 396748
rect 120763 396812 120829 396813
rect 120763 396748 120764 396812
rect 120828 396748 120829 396812
rect 120763 396747 120829 396748
rect 117234 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 117854 370894
rect 117234 370574 117854 370658
rect 117234 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 117854 370574
rect 117234 334894 117854 370338
rect 117234 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 117854 334894
rect 117234 334574 117854 334658
rect 117234 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 117854 334574
rect 117234 298894 117854 334338
rect 117234 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 117854 298894
rect 117234 298574 117854 298658
rect 117234 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 117854 298574
rect 117234 262894 117854 298338
rect 117234 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 117854 262894
rect 117234 262574 117854 262658
rect 117234 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 117854 262574
rect 117234 228924 117854 262338
rect 120954 374614 121574 398000
rect 123526 396813 123586 399470
rect 125918 399470 126028 399530
rect 128280 399530 128340 400106
rect 131000 399530 131060 400106
rect 133448 399530 133508 400106
rect 135896 399530 135956 400106
rect 138480 399530 138540 400106
rect 140928 399530 140988 400106
rect 128280 399470 128554 399530
rect 131000 399470 131130 399530
rect 133448 399470 133522 399530
rect 135896 399470 136098 399530
rect 125918 396813 125978 399470
rect 123523 396812 123589 396813
rect 123523 396748 123524 396812
rect 123588 396748 123589 396812
rect 123523 396747 123589 396748
rect 125915 396812 125981 396813
rect 125915 396748 125916 396812
rect 125980 396748 125981 396812
rect 125915 396747 125981 396748
rect 120954 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 121574 374614
rect 120954 374294 121574 374378
rect 120954 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 121574 374294
rect 120954 338614 121574 374058
rect 120954 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 121574 338614
rect 120954 338294 121574 338378
rect 120954 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 121574 338294
rect 120954 302614 121574 338058
rect 120954 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 121574 302614
rect 120954 302294 121574 302378
rect 120954 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 121574 302294
rect 120954 266614 121574 302058
rect 120954 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 121574 266614
rect 120954 266294 121574 266378
rect 120954 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 121574 266294
rect 120954 230614 121574 266058
rect 120954 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 121574 230614
rect 120954 230294 121574 230378
rect 120954 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 121574 230294
rect 120954 228924 121574 230058
rect 127794 381454 128414 398000
rect 128494 396810 128554 399470
rect 131070 396813 131130 399470
rect 128675 396812 128741 396813
rect 128675 396810 128676 396812
rect 128494 396750 128676 396810
rect 128675 396748 128676 396750
rect 128740 396748 128741 396812
rect 128675 396747 128741 396748
rect 131067 396812 131133 396813
rect 131067 396748 131068 396812
rect 131132 396748 131133 396812
rect 131067 396747 131133 396748
rect 127794 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 128414 381454
rect 127794 381134 128414 381218
rect 127794 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 128414 381134
rect 127794 345454 128414 380898
rect 127794 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 128414 345454
rect 127794 345134 128414 345218
rect 127794 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 128414 345134
rect 127794 309454 128414 344898
rect 127794 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 128414 309454
rect 127794 309134 128414 309218
rect 127794 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 128414 309134
rect 127794 273454 128414 308898
rect 127794 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 128414 273454
rect 127794 273134 128414 273218
rect 127794 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 128414 273134
rect 127794 237454 128414 272898
rect 127794 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 128414 237454
rect 127794 237134 128414 237218
rect 127794 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 128414 237134
rect 127794 228924 128414 236898
rect 131514 385174 132134 398000
rect 133462 396813 133522 399470
rect 133459 396812 133525 396813
rect 133459 396748 133460 396812
rect 133524 396748 133525 396812
rect 133459 396747 133525 396748
rect 131514 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 132134 385174
rect 131514 384854 132134 384938
rect 131514 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 132134 384854
rect 131514 349174 132134 384618
rect 131514 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 132134 349174
rect 131514 348854 132134 348938
rect 131514 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 132134 348854
rect 131514 313174 132134 348618
rect 131514 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 132134 313174
rect 131514 312854 132134 312938
rect 131514 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 132134 312854
rect 131514 277174 132134 312618
rect 131514 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 132134 277174
rect 131514 276854 132134 276938
rect 131514 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 132134 276854
rect 131514 241174 132134 276618
rect 131514 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 132134 241174
rect 131514 240854 132134 240938
rect 131514 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 132134 240854
rect 131514 228924 132134 240618
rect 135234 388894 135854 398000
rect 136038 397357 136098 399470
rect 138430 399470 138540 399530
rect 140822 399470 140988 399530
rect 143512 399530 143572 400106
rect 145960 399530 146020 400106
rect 143512 399470 143642 399530
rect 138430 397357 138490 399470
rect 136035 397356 136101 397357
rect 136035 397292 136036 397356
rect 136100 397292 136101 397356
rect 136035 397291 136101 397292
rect 138427 397356 138493 397357
rect 138427 397292 138428 397356
rect 138492 397292 138493 397356
rect 138427 397291 138493 397292
rect 135234 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 135854 388894
rect 135234 388574 135854 388658
rect 135234 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 135854 388574
rect 135234 352894 135854 388338
rect 135234 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 135854 352894
rect 135234 352574 135854 352658
rect 135234 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 135854 352574
rect 135234 316894 135854 352338
rect 135234 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 135854 316894
rect 135234 316574 135854 316658
rect 135234 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 135854 316574
rect 135234 280894 135854 316338
rect 135234 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 135854 280894
rect 135234 280574 135854 280658
rect 135234 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 135854 280574
rect 135234 244894 135854 280338
rect 135234 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 135854 244894
rect 135234 244574 135854 244658
rect 135234 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 135854 244574
rect 135234 228924 135854 244338
rect 138954 392614 139574 398000
rect 140822 396813 140882 399470
rect 143582 396813 143642 399470
rect 145606 399470 146020 399530
rect 148544 399530 148604 400106
rect 150992 399530 151052 400106
rect 148544 399470 148610 399530
rect 145606 396813 145666 399470
rect 140819 396812 140885 396813
rect 140819 396748 140820 396812
rect 140884 396748 140885 396812
rect 140819 396747 140885 396748
rect 143579 396812 143645 396813
rect 143579 396748 143580 396812
rect 143644 396748 143645 396812
rect 143579 396747 143645 396748
rect 145603 396812 145669 396813
rect 145603 396748 145604 396812
rect 145668 396748 145669 396812
rect 145603 396747 145669 396748
rect 138954 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 139574 392614
rect 138954 392294 139574 392378
rect 138954 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 139574 392294
rect 138954 356614 139574 392058
rect 138954 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 139574 356614
rect 138954 356294 139574 356378
rect 138954 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 139574 356294
rect 138954 320614 139574 356058
rect 138954 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 139574 320614
rect 138954 320294 139574 320378
rect 138954 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 139574 320294
rect 138954 284614 139574 320058
rect 138954 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 139574 284614
rect 138954 284294 139574 284378
rect 138954 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 139574 284294
rect 138954 248614 139574 284058
rect 138954 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 139574 248614
rect 138954 248294 139574 248378
rect 138954 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 139574 248294
rect 138954 228924 139574 248058
rect 145794 363454 146414 398000
rect 148550 396813 148610 399470
rect 150942 399470 151052 399530
rect 153440 399530 153500 400106
rect 155888 399530 155948 400106
rect 158472 399530 158532 400106
rect 160920 399530 160980 400106
rect 153440 399470 154130 399530
rect 155888 399470 155970 399530
rect 158472 399470 158546 399530
rect 148547 396812 148613 396813
rect 148547 396748 148548 396812
rect 148612 396748 148613 396812
rect 148547 396747 148613 396748
rect 145794 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 146414 363454
rect 145794 363134 146414 363218
rect 145794 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 146414 363134
rect 145794 327454 146414 362898
rect 145794 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 146414 327454
rect 145794 327134 146414 327218
rect 145794 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 146414 327134
rect 145794 291454 146414 326898
rect 145794 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 146414 291454
rect 145794 291134 146414 291218
rect 145794 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 146414 291134
rect 145794 255454 146414 290898
rect 145794 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 146414 255454
rect 145794 255134 146414 255218
rect 145794 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 146414 255134
rect 145794 228924 146414 254898
rect 149514 367174 150134 398000
rect 150942 397357 151002 399470
rect 150939 397356 151005 397357
rect 150939 397292 150940 397356
rect 151004 397292 151005 397356
rect 150939 397291 151005 397292
rect 149514 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 150134 367174
rect 149514 366854 150134 366938
rect 149514 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 150134 366854
rect 149514 331174 150134 366618
rect 149514 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 150134 331174
rect 149514 330854 150134 330938
rect 149514 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 150134 330854
rect 149514 295174 150134 330618
rect 149514 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 150134 295174
rect 149514 294854 150134 294938
rect 149514 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 150134 294854
rect 149514 259174 150134 294618
rect 149514 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 150134 259174
rect 149514 258854 150134 258938
rect 149514 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 150134 258854
rect 149514 228924 150134 258618
rect 153234 370894 153854 398000
rect 154070 396813 154130 399470
rect 155910 396813 155970 399470
rect 154067 396812 154133 396813
rect 154067 396748 154068 396812
rect 154132 396748 154133 396812
rect 154067 396747 154133 396748
rect 155907 396812 155973 396813
rect 155907 396748 155908 396812
rect 155972 396748 155973 396812
rect 155907 396747 155973 396748
rect 153234 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 153854 370894
rect 153234 370574 153854 370658
rect 153234 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 153854 370574
rect 153234 334894 153854 370338
rect 153234 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 153854 334894
rect 153234 334574 153854 334658
rect 153234 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 153854 334574
rect 153234 298894 153854 334338
rect 153234 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 153854 298894
rect 153234 298574 153854 298658
rect 153234 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 153854 298574
rect 153234 262894 153854 298338
rect 153234 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 153854 262894
rect 153234 262574 153854 262658
rect 153234 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 153854 262574
rect 153234 228924 153854 262338
rect 156954 374614 157574 398000
rect 158486 396813 158546 399470
rect 160878 399470 160980 399530
rect 163368 399530 163428 400106
rect 165952 399530 166012 400106
rect 183224 399530 183284 400106
rect 163368 399470 163514 399530
rect 165952 399470 166090 399530
rect 160878 396813 160938 399470
rect 163454 396813 163514 399470
rect 158483 396812 158549 396813
rect 158483 396748 158484 396812
rect 158548 396748 158549 396812
rect 158483 396747 158549 396748
rect 160875 396812 160941 396813
rect 160875 396748 160876 396812
rect 160940 396748 160941 396812
rect 160875 396747 160941 396748
rect 163451 396812 163517 396813
rect 163451 396748 163452 396812
rect 163516 396748 163517 396812
rect 163451 396747 163517 396748
rect 156954 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 157574 374614
rect 156954 374294 157574 374378
rect 156954 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 157574 374294
rect 156954 338614 157574 374058
rect 156954 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 157574 338614
rect 156954 338294 157574 338378
rect 156954 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 157574 338294
rect 156954 302614 157574 338058
rect 156954 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 157574 302614
rect 156954 302294 157574 302378
rect 156954 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 157574 302294
rect 156954 266614 157574 302058
rect 156954 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 157574 266614
rect 156954 266294 157574 266378
rect 156954 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 157574 266294
rect 156954 230614 157574 266058
rect 156954 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 157574 230614
rect 156954 230294 157574 230378
rect 156954 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 157574 230294
rect 156954 228924 157574 230058
rect 163794 381454 164414 398000
rect 166030 396813 166090 399470
rect 183142 399470 183284 399530
rect 183360 399530 183420 400106
rect 183360 399470 183570 399530
rect 166027 396812 166093 396813
rect 166027 396748 166028 396812
rect 166092 396748 166093 396812
rect 166027 396747 166093 396748
rect 163794 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 164414 381454
rect 163794 381134 164414 381218
rect 163794 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 164414 381134
rect 163794 345454 164414 380898
rect 163794 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 164414 345454
rect 163794 345134 164414 345218
rect 163794 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 164414 345134
rect 163794 309454 164414 344898
rect 163794 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 164414 309454
rect 163794 309134 164414 309218
rect 163794 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 164414 309134
rect 163794 273454 164414 308898
rect 163794 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 164414 273454
rect 163794 273134 164414 273218
rect 163794 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 164414 273134
rect 163794 237454 164414 272898
rect 163794 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 164414 237454
rect 163794 237134 164414 237218
rect 163794 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 164414 237134
rect 163794 228924 164414 236898
rect 167514 385174 168134 398000
rect 167514 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 168134 385174
rect 167514 384854 168134 384938
rect 167514 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 168134 384854
rect 167514 349174 168134 384618
rect 167514 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 168134 349174
rect 167514 348854 168134 348938
rect 167514 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 168134 348854
rect 167514 313174 168134 348618
rect 167514 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 168134 313174
rect 167514 312854 168134 312938
rect 167514 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 168134 312854
rect 167514 277174 168134 312618
rect 167514 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 168134 277174
rect 167514 276854 168134 276938
rect 167514 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 168134 276854
rect 167514 241174 168134 276618
rect 167514 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 168134 241174
rect 167514 240854 168134 240938
rect 167514 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 168134 240854
rect 167514 228924 168134 240618
rect 171234 388894 171854 398000
rect 171234 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 171854 388894
rect 171234 388574 171854 388658
rect 171234 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 171854 388574
rect 171234 352894 171854 388338
rect 171234 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 171854 352894
rect 171234 352574 171854 352658
rect 171234 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 171854 352574
rect 171234 316894 171854 352338
rect 171234 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 171854 316894
rect 171234 316574 171854 316658
rect 171234 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 171854 316574
rect 171234 280894 171854 316338
rect 171234 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 171854 280894
rect 171234 280574 171854 280658
rect 171234 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 171854 280574
rect 171234 244894 171854 280338
rect 171234 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 171854 244894
rect 171234 244574 171854 244658
rect 171234 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 171854 244574
rect 171234 228924 171854 244338
rect 174954 392614 175574 398000
rect 174954 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 175574 392614
rect 174954 392294 175574 392378
rect 174954 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 175574 392294
rect 174954 356614 175574 392058
rect 174954 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 175574 356614
rect 174954 356294 175574 356378
rect 174954 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 175574 356294
rect 174954 320614 175574 356058
rect 174954 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 175574 320614
rect 174954 320294 175574 320378
rect 174954 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 175574 320294
rect 174954 284614 175574 320058
rect 174954 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 175574 284614
rect 174954 284294 175574 284378
rect 174954 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 175574 284294
rect 174954 248614 175574 284058
rect 174954 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 175574 248614
rect 174954 248294 175574 248378
rect 174954 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 175574 248294
rect 174954 228924 175574 248058
rect 181794 363454 182414 398000
rect 183142 396813 183202 399470
rect 183510 397357 183570 399470
rect 183507 397356 183573 397357
rect 183507 397292 183508 397356
rect 183572 397292 183573 397356
rect 183507 397291 183573 397292
rect 183139 396812 183205 396813
rect 183139 396748 183140 396812
rect 183204 396748 183205 396812
rect 183139 396747 183205 396748
rect 181794 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 182414 363454
rect 181794 363134 182414 363218
rect 181794 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 182414 363134
rect 181794 327454 182414 362898
rect 181794 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 182414 327454
rect 181794 327134 182414 327218
rect 181794 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 182414 327134
rect 181794 291454 182414 326898
rect 181794 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 182414 291454
rect 181794 291134 182414 291218
rect 181794 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 182414 291134
rect 181794 255454 182414 290898
rect 181794 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 182414 255454
rect 181794 255134 182414 255218
rect 181794 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 182414 255134
rect 181794 228924 182414 254898
rect 185514 367174 186134 398000
rect 185514 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 186134 367174
rect 185514 366854 186134 366938
rect 185514 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 186134 366854
rect 185514 331174 186134 366618
rect 185514 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 186134 331174
rect 185514 330854 186134 330938
rect 185514 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 186134 330854
rect 185514 295174 186134 330618
rect 185514 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 186134 295174
rect 185514 294854 186134 294938
rect 185514 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 186134 294854
rect 185514 259174 186134 294618
rect 185514 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 186134 259174
rect 185514 258854 186134 258938
rect 185514 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 186134 258854
rect 185514 228924 186134 258618
rect 189234 370894 189854 398000
rect 189234 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 189854 370894
rect 189234 370574 189854 370658
rect 189234 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 189854 370574
rect 189234 334894 189854 370338
rect 189234 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 189854 334894
rect 189234 334574 189854 334658
rect 189234 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 189854 334574
rect 189234 298894 189854 334338
rect 189234 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 189854 298894
rect 189234 298574 189854 298658
rect 189234 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 189854 298574
rect 189234 262894 189854 298338
rect 189234 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 189854 262894
rect 189234 262574 189854 262658
rect 189234 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 189854 262574
rect 189234 228924 189854 262338
rect 192954 374614 193574 398000
rect 192954 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 193574 374614
rect 192954 374294 193574 374378
rect 192954 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 193574 374294
rect 192954 338614 193574 374058
rect 192954 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 193574 338614
rect 192954 338294 193574 338378
rect 192954 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 193574 338294
rect 192954 302614 193574 338058
rect 192954 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 193574 302614
rect 192954 302294 193574 302378
rect 192954 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 193574 302294
rect 192954 266614 193574 302058
rect 192954 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 193574 266614
rect 192954 266294 193574 266378
rect 192954 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 193574 266294
rect 192954 230614 193574 266058
rect 192954 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 193574 230614
rect 192954 230294 193574 230378
rect 192954 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 193574 230294
rect 192954 228924 193574 230058
rect 199794 381454 200414 416898
rect 199794 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 200414 381454
rect 199794 381134 200414 381218
rect 199794 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 200414 381134
rect 199794 345454 200414 380898
rect 199794 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 200414 345454
rect 199794 345134 200414 345218
rect 199794 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 200414 345134
rect 199794 309454 200414 344898
rect 199794 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 200414 309454
rect 199794 309134 200414 309218
rect 199794 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 200414 309134
rect 199794 273454 200414 308898
rect 199794 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 200414 273454
rect 199794 273134 200414 273218
rect 199794 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 200414 273134
rect 199794 237454 200414 272898
rect 199794 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 200414 237454
rect 199794 237134 200414 237218
rect 199794 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 200414 237134
rect 199794 228924 200414 236898
rect 203514 673174 204134 707162
rect 203514 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 204134 673174
rect 203514 672854 204134 672938
rect 203514 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 204134 672854
rect 203514 637174 204134 672618
rect 203514 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 204134 637174
rect 203514 636854 204134 636938
rect 203514 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 204134 636854
rect 203514 601174 204134 636618
rect 203514 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 204134 601174
rect 203514 600854 204134 600938
rect 203514 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 204134 600854
rect 203514 565174 204134 600618
rect 203514 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 204134 565174
rect 203514 564854 204134 564938
rect 203514 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 204134 564854
rect 203514 529174 204134 564618
rect 203514 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 204134 529174
rect 203514 528854 204134 528938
rect 203514 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 204134 528854
rect 203514 493174 204134 528618
rect 203514 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 204134 493174
rect 203514 492854 204134 492938
rect 203514 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 204134 492854
rect 203514 457174 204134 492618
rect 203514 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 204134 457174
rect 203514 456854 204134 456938
rect 203514 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 204134 456854
rect 203514 421174 204134 456618
rect 203514 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 204134 421174
rect 203514 420854 204134 420938
rect 203514 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 204134 420854
rect 203514 385174 204134 420618
rect 203514 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 204134 385174
rect 203514 384854 204134 384938
rect 203514 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 204134 384854
rect 203514 349174 204134 384618
rect 203514 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 204134 349174
rect 203514 348854 204134 348938
rect 203514 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 204134 348854
rect 203514 313174 204134 348618
rect 203514 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 204134 313174
rect 203514 312854 204134 312938
rect 203514 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 204134 312854
rect 203514 277174 204134 312618
rect 203514 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 204134 277174
rect 203514 276854 204134 276938
rect 203514 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 204134 276854
rect 203514 241174 204134 276618
rect 203514 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 204134 241174
rect 203514 240854 204134 240938
rect 203514 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 204134 240854
rect 203514 228924 204134 240618
rect 207234 676894 207854 709082
rect 207234 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 207854 676894
rect 207234 676574 207854 676658
rect 207234 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 207854 676574
rect 207234 640894 207854 676338
rect 207234 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 207854 640894
rect 207234 640574 207854 640658
rect 207234 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 207854 640574
rect 207234 604894 207854 640338
rect 207234 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 207854 604894
rect 207234 604574 207854 604658
rect 207234 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 207854 604574
rect 207234 568894 207854 604338
rect 207234 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 207854 568894
rect 207234 568574 207854 568658
rect 207234 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 207854 568574
rect 207234 532894 207854 568338
rect 207234 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 207854 532894
rect 207234 532574 207854 532658
rect 207234 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 207854 532574
rect 207234 496894 207854 532338
rect 207234 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 207854 496894
rect 207234 496574 207854 496658
rect 207234 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 207854 496574
rect 207234 460894 207854 496338
rect 207234 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 207854 460894
rect 207234 460574 207854 460658
rect 207234 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 207854 460574
rect 207234 424894 207854 460338
rect 207234 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 207854 424894
rect 207234 424574 207854 424658
rect 207234 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 207854 424574
rect 207234 388894 207854 424338
rect 207234 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 207854 388894
rect 207234 388574 207854 388658
rect 207234 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 207854 388574
rect 207234 352894 207854 388338
rect 207234 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 207854 352894
rect 207234 352574 207854 352658
rect 207234 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 207854 352574
rect 207234 316894 207854 352338
rect 207234 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 207854 316894
rect 207234 316574 207854 316658
rect 207234 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 207854 316574
rect 207234 280894 207854 316338
rect 207234 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 207854 280894
rect 207234 280574 207854 280658
rect 207234 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 207854 280574
rect 207234 244894 207854 280338
rect 207234 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 207854 244894
rect 207234 244574 207854 244658
rect 207234 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 207854 244574
rect 207234 228924 207854 244338
rect 210954 680614 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 210954 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 211574 680614
rect 210954 680294 211574 680378
rect 210954 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 211574 680294
rect 210954 644614 211574 680058
rect 210954 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 211574 644614
rect 210954 644294 211574 644378
rect 210954 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 211574 644294
rect 210954 608614 211574 644058
rect 210954 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 211574 608614
rect 210954 608294 211574 608378
rect 210954 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 211574 608294
rect 210954 572614 211574 608058
rect 210954 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 211574 572614
rect 210954 572294 211574 572378
rect 210954 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 211574 572294
rect 210954 536614 211574 572058
rect 210954 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 211574 536614
rect 210954 536294 211574 536378
rect 210954 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 211574 536294
rect 210954 500614 211574 536058
rect 210954 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 211574 500614
rect 210954 500294 211574 500378
rect 210954 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 211574 500294
rect 210954 464614 211574 500058
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 687454 218414 704282
rect 217794 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 218414 687454
rect 217794 687134 218414 687218
rect 217794 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 218414 687134
rect 217794 651454 218414 686898
rect 217794 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 218414 651454
rect 217794 651134 218414 651218
rect 217794 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 218414 651134
rect 217794 615454 218414 650898
rect 217794 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 218414 615454
rect 217794 615134 218414 615218
rect 217794 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 218414 615134
rect 217794 579454 218414 614898
rect 217794 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 218414 579454
rect 217794 579134 218414 579218
rect 217794 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 218414 579134
rect 217794 543454 218414 578898
rect 217794 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 218414 543454
rect 217794 543134 218414 543218
rect 217794 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 218414 543134
rect 217794 507454 218414 542898
rect 217794 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 218414 507454
rect 217794 507134 218414 507218
rect 217794 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 218414 507134
rect 217547 487116 217613 487117
rect 217547 487052 217548 487116
rect 217612 487052 217613 487116
rect 217547 487051 217613 487052
rect 217550 485210 217610 487051
rect 217794 485308 218414 506898
rect 221514 691174 222134 706202
rect 221514 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 222134 691174
rect 221514 690854 222134 690938
rect 221514 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 222134 690854
rect 221514 655174 222134 690618
rect 221514 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 222134 655174
rect 221514 654854 222134 654938
rect 221514 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 222134 654854
rect 221514 619174 222134 654618
rect 221514 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 222134 619174
rect 221514 618854 222134 618938
rect 221514 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 222134 618854
rect 221514 583174 222134 618618
rect 221514 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 222134 583174
rect 221514 582854 222134 582938
rect 221514 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 222134 582854
rect 221514 547174 222134 582618
rect 221514 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 222134 547174
rect 221514 546854 222134 546938
rect 221514 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 222134 546854
rect 221514 511174 222134 546618
rect 221514 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 222134 511174
rect 221514 510854 222134 510938
rect 221514 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 222134 510854
rect 218651 491468 218717 491469
rect 218651 491404 218652 491468
rect 218716 491404 218717 491468
rect 218651 491403 218717 491404
rect 217550 485150 218162 485210
rect 218102 480317 218162 485150
rect 218099 480316 218165 480317
rect 218099 480252 218100 480316
rect 218164 480252 218165 480316
rect 218099 480251 218165 480252
rect 218467 479908 218533 479909
rect 218467 479844 218468 479908
rect 218532 479844 218533 479908
rect 218467 479843 218533 479844
rect 218470 470797 218530 479843
rect 218467 470796 218533 470797
rect 218467 470732 218468 470796
rect 218532 470732 218533 470796
rect 218467 470731 218533 470732
rect 218467 470524 218533 470525
rect 218467 470460 218468 470524
rect 218532 470460 218533 470524
rect 218467 470459 218533 470460
rect 210954 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 211574 464614
rect 210954 464294 211574 464378
rect 210954 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 211574 464294
rect 210954 428614 211574 464058
rect 218470 461005 218530 470459
rect 218467 461004 218533 461005
rect 218467 460940 218468 461004
rect 218532 460940 218533 461004
rect 218467 460939 218533 460940
rect 218467 460868 218533 460869
rect 218467 460804 218468 460868
rect 218532 460804 218533 460868
rect 218467 460803 218533 460804
rect 218470 451349 218530 460803
rect 218467 451348 218533 451349
rect 218467 451284 218468 451348
rect 218532 451284 218533 451348
rect 218467 451283 218533 451284
rect 218467 451212 218533 451213
rect 218467 451148 218468 451212
rect 218532 451148 218533 451212
rect 218467 451147 218533 451148
rect 218470 441693 218530 451147
rect 218467 441692 218533 441693
rect 218467 441628 218468 441692
rect 218532 441628 218533 441692
rect 218467 441627 218533 441628
rect 218467 441556 218533 441557
rect 218467 441492 218468 441556
rect 218532 441492 218533 441556
rect 218467 441491 218533 441492
rect 218470 432037 218530 441491
rect 218467 432036 218533 432037
rect 218467 431972 218468 432036
rect 218532 431972 218533 432036
rect 218467 431971 218533 431972
rect 218467 431900 218533 431901
rect 218467 431836 218468 431900
rect 218532 431836 218533 431900
rect 218467 431835 218533 431836
rect 210954 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 211574 428614
rect 210954 428294 211574 428378
rect 210954 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 211574 428294
rect 210954 392614 211574 428058
rect 218470 422381 218530 431835
rect 218467 422380 218533 422381
rect 218467 422316 218468 422380
rect 218532 422316 218533 422380
rect 218467 422315 218533 422316
rect 218467 422244 218533 422245
rect 218467 422180 218468 422244
rect 218532 422180 218533 422244
rect 218467 422179 218533 422180
rect 218470 412725 218530 422179
rect 218467 412724 218533 412725
rect 218467 412660 218468 412724
rect 218532 412660 218533 412724
rect 218467 412659 218533 412660
rect 218467 412588 218533 412589
rect 218467 412524 218468 412588
rect 218532 412524 218533 412588
rect 218467 412523 218533 412524
rect 218470 403069 218530 412523
rect 218467 403068 218533 403069
rect 218467 403004 218468 403068
rect 218532 403004 218533 403068
rect 218467 403003 218533 403004
rect 218467 402932 218533 402933
rect 218467 402868 218468 402932
rect 218532 402868 218533 402932
rect 218467 402867 218533 402868
rect 218470 398309 218530 402867
rect 218467 398308 218533 398309
rect 218467 398244 218468 398308
rect 218532 398244 218533 398308
rect 218467 398243 218533 398244
rect 210954 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 211574 392614
rect 210954 392294 211574 392378
rect 210954 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 211574 392294
rect 210954 356614 211574 392058
rect 210954 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 211574 356614
rect 210954 356294 211574 356378
rect 210954 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 211574 356294
rect 210954 320614 211574 356058
rect 210954 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 211574 320614
rect 210954 320294 211574 320378
rect 210954 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 211574 320294
rect 210954 284614 211574 320058
rect 210954 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 211574 284614
rect 210954 284294 211574 284378
rect 210954 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 211574 284294
rect 210954 248614 211574 284058
rect 210954 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 211574 248614
rect 210954 248294 211574 248378
rect 210954 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 211574 248294
rect 210954 228924 211574 248058
rect 217794 363454 218414 398000
rect 217794 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 218414 363454
rect 217794 363134 218414 363218
rect 217794 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 218414 363134
rect 217794 327454 218414 362898
rect 217794 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 218414 327454
rect 217794 327134 218414 327218
rect 217794 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 218414 327134
rect 217794 291454 218414 326898
rect 217794 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 218414 291454
rect 217794 291134 218414 291218
rect 217794 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 218414 291134
rect 217794 255454 218414 290898
rect 217794 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 218414 255454
rect 217794 255134 218414 255218
rect 217794 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 218414 255134
rect 217794 228924 218414 254898
rect 218654 238509 218714 491403
rect 218835 491332 218901 491333
rect 218835 491268 218836 491332
rect 218900 491268 218901 491332
rect 218835 491267 218901 491268
rect 218651 238508 218717 238509
rect 218651 238444 218652 238508
rect 218716 238444 218717 238508
rect 218651 238443 218717 238444
rect 218838 238370 218898 491267
rect 219203 490244 219269 490245
rect 219203 490180 219204 490244
rect 219268 490180 219269 490244
rect 219203 490179 219269 490180
rect 219206 489930 219266 490179
rect 219206 489870 219450 489930
rect 219390 489290 219450 489870
rect 219206 489230 219450 489290
rect 219019 485484 219085 485485
rect 219019 485420 219020 485484
rect 219084 485420 219085 485484
rect 219019 485419 219085 485420
rect 218654 238310 218898 238370
rect 218654 234293 218714 238310
rect 218835 238236 218901 238237
rect 218835 238172 218836 238236
rect 218900 238172 218901 238236
rect 218835 238171 218901 238172
rect 218651 234292 218717 234293
rect 218651 234228 218652 234292
rect 218716 234228 218717 234292
rect 218651 234227 218717 234228
rect 218838 234157 218898 238171
rect 218835 234156 218901 234157
rect 218835 234092 218836 234156
rect 218900 234092 218901 234156
rect 218835 234091 218901 234092
rect 219022 228853 219082 485419
rect 219206 479909 219266 489230
rect 221514 485308 222134 510618
rect 225234 694894 225854 708122
rect 225234 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 225854 694894
rect 225234 694574 225854 694658
rect 225234 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 225854 694574
rect 225234 658894 225854 694338
rect 225234 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 225854 658894
rect 225234 658574 225854 658658
rect 225234 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 225854 658574
rect 225234 622894 225854 658338
rect 225234 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 225854 622894
rect 225234 622574 225854 622658
rect 225234 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 225854 622574
rect 225234 586894 225854 622338
rect 225234 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 225854 586894
rect 225234 586574 225854 586658
rect 225234 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 225854 586574
rect 225234 550894 225854 586338
rect 225234 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 225854 550894
rect 225234 550574 225854 550658
rect 225234 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 225854 550574
rect 225234 514894 225854 550338
rect 225234 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 225854 514894
rect 225234 514574 225854 514658
rect 225234 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 225854 514574
rect 225234 485308 225854 514338
rect 228954 698614 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 228954 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 229574 698614
rect 228954 698294 229574 698378
rect 228954 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 229574 698294
rect 228954 662614 229574 698058
rect 228954 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 229574 662614
rect 228954 662294 229574 662378
rect 228954 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 229574 662294
rect 228954 626614 229574 662058
rect 228954 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 229574 626614
rect 228954 626294 229574 626378
rect 228954 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 229574 626294
rect 228954 590614 229574 626058
rect 228954 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 229574 590614
rect 228954 590294 229574 590378
rect 228954 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 229574 590294
rect 228954 554614 229574 590058
rect 228954 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 229574 554614
rect 228954 554294 229574 554378
rect 228954 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 229574 554294
rect 228954 518614 229574 554058
rect 228954 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 229574 518614
rect 228954 518294 229574 518378
rect 228954 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 229574 518294
rect 228954 485308 229574 518058
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 669454 236414 705242
rect 235794 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 236414 669454
rect 235794 669134 236414 669218
rect 235794 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 236414 669134
rect 235794 633454 236414 668898
rect 235794 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 236414 633454
rect 235794 633134 236414 633218
rect 235794 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 236414 633134
rect 235794 597454 236414 632898
rect 235794 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 236414 597454
rect 235794 597134 236414 597218
rect 235794 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 236414 597134
rect 235794 561454 236414 596898
rect 235794 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 236414 561454
rect 235794 561134 236414 561218
rect 235794 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 236414 561134
rect 235794 525454 236414 560898
rect 235794 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 236414 525454
rect 235794 525134 236414 525218
rect 235794 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 236414 525134
rect 235794 489454 236414 524898
rect 235794 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 236414 489454
rect 235794 489134 236414 489218
rect 235794 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 236414 489134
rect 235794 485308 236414 488898
rect 239514 673174 240134 707162
rect 239514 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 240134 673174
rect 239514 672854 240134 672938
rect 239514 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 240134 672854
rect 239514 637174 240134 672618
rect 239514 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 240134 637174
rect 239514 636854 240134 636938
rect 239514 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 240134 636854
rect 239514 601174 240134 636618
rect 239514 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 240134 601174
rect 239514 600854 240134 600938
rect 239514 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 240134 600854
rect 239514 565174 240134 600618
rect 239514 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 240134 565174
rect 239514 564854 240134 564938
rect 239514 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 240134 564854
rect 239514 529174 240134 564618
rect 239514 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 240134 529174
rect 239514 528854 240134 528938
rect 239514 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 240134 528854
rect 239514 493174 240134 528618
rect 239514 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 240134 493174
rect 239514 492854 240134 492938
rect 239514 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 240134 492854
rect 239514 485308 240134 492618
rect 243234 676894 243854 709082
rect 243234 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 243854 676894
rect 243234 676574 243854 676658
rect 243234 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 243854 676574
rect 243234 640894 243854 676338
rect 243234 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 243854 640894
rect 243234 640574 243854 640658
rect 243234 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 243854 640574
rect 243234 604894 243854 640338
rect 243234 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 243854 604894
rect 243234 604574 243854 604658
rect 243234 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 243854 604574
rect 243234 568894 243854 604338
rect 243234 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 243854 568894
rect 243234 568574 243854 568658
rect 243234 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 243854 568574
rect 243234 532894 243854 568338
rect 243234 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 243854 532894
rect 243234 532574 243854 532658
rect 243234 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 243854 532574
rect 243234 496894 243854 532338
rect 243234 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 243854 496894
rect 243234 496574 243854 496658
rect 243234 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 243854 496574
rect 243234 485308 243854 496338
rect 246954 680614 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 246954 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 247574 680614
rect 246954 680294 247574 680378
rect 246954 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 247574 680294
rect 246954 644614 247574 680058
rect 246954 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 247574 644614
rect 246954 644294 247574 644378
rect 246954 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 247574 644294
rect 246954 608614 247574 644058
rect 246954 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 247574 608614
rect 246954 608294 247574 608378
rect 246954 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 247574 608294
rect 246954 572614 247574 608058
rect 246954 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 247574 572614
rect 246954 572294 247574 572378
rect 246954 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 247574 572294
rect 246954 536614 247574 572058
rect 246954 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 247574 536614
rect 246954 536294 247574 536378
rect 246954 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 247574 536294
rect 246954 500614 247574 536058
rect 246954 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 247574 500614
rect 246954 500294 247574 500378
rect 246954 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 247574 500294
rect 246954 485308 247574 500058
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 687454 254414 704282
rect 253794 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 254414 687454
rect 253794 687134 254414 687218
rect 253794 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 254414 687134
rect 253794 651454 254414 686898
rect 253794 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 254414 651454
rect 253794 651134 254414 651218
rect 253794 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 254414 651134
rect 253794 615454 254414 650898
rect 253794 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 254414 615454
rect 253794 615134 254414 615218
rect 253794 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 254414 615134
rect 253794 579454 254414 614898
rect 253794 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 254414 579454
rect 253794 579134 254414 579218
rect 253794 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 254414 579134
rect 253794 543454 254414 578898
rect 253794 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 254414 543454
rect 253794 543134 254414 543218
rect 253794 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 254414 543134
rect 253794 507454 254414 542898
rect 253794 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 254414 507454
rect 253794 507134 254414 507218
rect 253794 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 254414 507134
rect 248643 486844 248709 486845
rect 248643 486780 248644 486844
rect 248708 486780 248709 486844
rect 248643 486779 248709 486780
rect 219939 485076 220005 485077
rect 219939 485012 219940 485076
rect 220004 485012 220005 485076
rect 219939 485011 220005 485012
rect 219571 484260 219637 484261
rect 219571 484196 219572 484260
rect 219636 484196 219637 484260
rect 219571 484195 219637 484196
rect 219387 480316 219453 480317
rect 219387 480252 219388 480316
rect 219452 480252 219453 480316
rect 219387 480251 219453 480252
rect 219203 479908 219269 479909
rect 219203 479844 219204 479908
rect 219268 479844 219269 479908
rect 219203 479843 219269 479844
rect 219390 479770 219450 480251
rect 219206 479710 219450 479770
rect 219206 470930 219266 479710
rect 219206 470870 219450 470930
rect 219203 470796 219269 470797
rect 219203 470732 219204 470796
rect 219268 470732 219269 470796
rect 219203 470731 219269 470732
rect 219206 392869 219266 470731
rect 219390 470525 219450 470870
rect 219387 470524 219453 470525
rect 219387 470460 219388 470524
rect 219452 470460 219453 470524
rect 219387 470459 219453 470460
rect 219387 461004 219453 461005
rect 219387 460940 219388 461004
rect 219452 460940 219453 461004
rect 219387 460939 219453 460940
rect 219390 460869 219450 460939
rect 219387 460868 219453 460869
rect 219387 460804 219388 460868
rect 219452 460804 219453 460868
rect 219387 460803 219453 460804
rect 219387 451348 219453 451349
rect 219387 451284 219388 451348
rect 219452 451284 219453 451348
rect 219387 451283 219453 451284
rect 219390 451213 219450 451283
rect 219387 451212 219453 451213
rect 219387 451148 219388 451212
rect 219452 451148 219453 451212
rect 219387 451147 219453 451148
rect 219387 441692 219453 441693
rect 219387 441628 219388 441692
rect 219452 441628 219453 441692
rect 219387 441627 219453 441628
rect 219390 441557 219450 441627
rect 219387 441556 219453 441557
rect 219387 441492 219388 441556
rect 219452 441492 219453 441556
rect 219387 441491 219453 441492
rect 219387 432036 219453 432037
rect 219387 431972 219388 432036
rect 219452 431972 219453 432036
rect 219387 431971 219453 431972
rect 219390 431901 219450 431971
rect 219387 431900 219453 431901
rect 219387 431836 219388 431900
rect 219452 431836 219453 431900
rect 219387 431835 219453 431836
rect 219387 422380 219453 422381
rect 219387 422316 219388 422380
rect 219452 422316 219453 422380
rect 219387 422315 219453 422316
rect 219390 422245 219450 422315
rect 219387 422244 219453 422245
rect 219387 422180 219388 422244
rect 219452 422180 219453 422244
rect 219387 422179 219453 422180
rect 219387 412724 219453 412725
rect 219387 412660 219388 412724
rect 219452 412660 219453 412724
rect 219387 412659 219453 412660
rect 219390 412589 219450 412659
rect 219387 412588 219453 412589
rect 219387 412524 219388 412588
rect 219452 412524 219453 412588
rect 219387 412523 219453 412524
rect 219574 403341 219634 484195
rect 219755 483444 219821 483445
rect 219755 483380 219756 483444
rect 219820 483380 219821 483444
rect 219755 483379 219821 483380
rect 219571 403340 219637 403341
rect 219571 403276 219572 403340
rect 219636 403276 219637 403340
rect 219571 403275 219637 403276
rect 219571 403204 219637 403205
rect 219571 403140 219572 403204
rect 219636 403140 219637 403204
rect 219571 403139 219637 403140
rect 219387 403068 219453 403069
rect 219387 403004 219388 403068
rect 219452 403004 219453 403068
rect 219387 403003 219453 403004
rect 219390 402933 219450 403003
rect 219387 402932 219453 402933
rect 219387 402868 219388 402932
rect 219452 402868 219453 402932
rect 219387 402867 219453 402868
rect 219574 399941 219634 403139
rect 219571 399940 219637 399941
rect 219571 399876 219572 399940
rect 219636 399876 219637 399940
rect 219571 399875 219637 399876
rect 219758 398037 219818 483379
rect 219942 398173 220002 485011
rect 248646 483850 248706 486779
rect 253427 485892 253493 485893
rect 253427 485828 253428 485892
rect 253492 485828 253493 485892
rect 253427 485827 253493 485828
rect 251035 485212 251101 485213
rect 251035 485148 251036 485212
rect 251100 485148 251101 485212
rect 251035 485147 251101 485148
rect 251038 483850 251098 485147
rect 248646 483790 248764 483850
rect 248704 483202 248764 483790
rect 251016 483790 251098 483850
rect 253430 483850 253490 485827
rect 253794 485308 254414 506898
rect 257514 691174 258134 706202
rect 257514 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 258134 691174
rect 257514 690854 258134 690938
rect 257514 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 258134 690854
rect 257514 655174 258134 690618
rect 257514 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 258134 655174
rect 257514 654854 258134 654938
rect 257514 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 258134 654854
rect 257514 619174 258134 654618
rect 257514 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 258134 619174
rect 257514 618854 258134 618938
rect 257514 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 258134 618854
rect 257514 583174 258134 618618
rect 257514 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 258134 583174
rect 257514 582854 258134 582938
rect 257514 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 258134 582854
rect 257514 547174 258134 582618
rect 257514 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 258134 547174
rect 257514 546854 258134 546938
rect 257514 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 258134 546854
rect 257514 511174 258134 546618
rect 257514 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 258134 511174
rect 257514 510854 258134 510938
rect 257514 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 258134 510854
rect 256187 485892 256253 485893
rect 256187 485828 256188 485892
rect 256252 485828 256253 485892
rect 256187 485827 256253 485828
rect 256190 483850 256250 485827
rect 257514 485308 258134 510618
rect 261234 694894 261854 708122
rect 261234 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 261854 694894
rect 261234 694574 261854 694658
rect 261234 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 261854 694574
rect 261234 658894 261854 694338
rect 261234 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 261854 658894
rect 261234 658574 261854 658658
rect 261234 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 261854 658574
rect 261234 622894 261854 658338
rect 261234 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 261854 622894
rect 261234 622574 261854 622658
rect 261234 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 261854 622574
rect 261234 586894 261854 622338
rect 261234 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 261854 586894
rect 261234 586574 261854 586658
rect 261234 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 261854 586574
rect 261234 550894 261854 586338
rect 261234 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 261854 550894
rect 261234 550574 261854 550658
rect 261234 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 261854 550574
rect 261234 514894 261854 550338
rect 261234 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 261854 514894
rect 261234 514574 261854 514658
rect 261234 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 261854 514574
rect 260971 485620 261037 485621
rect 260971 485556 260972 485620
rect 261036 485556 261037 485620
rect 260971 485555 261037 485556
rect 258395 483988 258461 483989
rect 258395 483924 258396 483988
rect 258460 483924 258461 483988
rect 258395 483923 258461 483924
rect 253430 483790 253524 483850
rect 251016 483202 251076 483790
rect 253464 483202 253524 483790
rect 256184 483790 256250 483850
rect 258398 483850 258458 483923
rect 260974 483850 261034 485555
rect 261234 485308 261854 514338
rect 264954 698614 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 264954 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 265574 698614
rect 264954 698294 265574 698378
rect 264954 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 265574 698294
rect 264954 662614 265574 698058
rect 264954 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 265574 662614
rect 264954 662294 265574 662378
rect 264954 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 265574 662294
rect 264954 626614 265574 662058
rect 264954 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 265574 626614
rect 264954 626294 265574 626378
rect 264954 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 265574 626294
rect 264954 590614 265574 626058
rect 264954 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 265574 590614
rect 264954 590294 265574 590378
rect 264954 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 265574 590294
rect 264954 554614 265574 590058
rect 264954 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 265574 554614
rect 264954 554294 265574 554378
rect 264954 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 265574 554294
rect 264954 518614 265574 554058
rect 264954 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 265574 518614
rect 264954 518294 265574 518378
rect 264954 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 265574 518294
rect 263547 485892 263613 485893
rect 263547 485828 263548 485892
rect 263612 485828 263613 485892
rect 263547 485827 263613 485828
rect 263550 483850 263610 485827
rect 264954 485308 265574 518058
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 669454 272414 705242
rect 271794 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 272414 669454
rect 271794 669134 272414 669218
rect 271794 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 272414 669134
rect 271794 633454 272414 668898
rect 271794 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 272414 633454
rect 271794 633134 272414 633218
rect 271794 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 272414 633134
rect 271794 597454 272414 632898
rect 271794 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 272414 597454
rect 271794 597134 272414 597218
rect 271794 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 272414 597134
rect 271794 561454 272414 596898
rect 271794 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 272414 561454
rect 271794 561134 272414 561218
rect 271794 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 272414 561134
rect 271794 525454 272414 560898
rect 271794 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 272414 525454
rect 271794 525134 272414 525218
rect 271794 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 272414 525134
rect 271794 489454 272414 524898
rect 271794 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 272414 489454
rect 271794 489134 272414 489218
rect 271794 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 272414 489134
rect 271091 487524 271157 487525
rect 271091 487460 271092 487524
rect 271156 487460 271157 487524
rect 271091 487459 271157 487460
rect 266123 486844 266189 486845
rect 266123 486780 266124 486844
rect 266188 486780 266189 486844
rect 266123 486779 266189 486780
rect 266126 483850 266186 486779
rect 268515 484940 268581 484941
rect 268515 484876 268516 484940
rect 268580 484876 268581 484940
rect 268515 484875 268581 484876
rect 258398 483790 258556 483850
rect 260974 483790 261140 483850
rect 256184 483202 256244 483790
rect 258496 483202 258556 483790
rect 261080 483202 261140 483790
rect 263528 483790 263610 483850
rect 266112 483790 266186 483850
rect 268518 483850 268578 484875
rect 271094 483850 271154 487459
rect 271794 485308 272414 488898
rect 275514 673174 276134 707162
rect 275514 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 276134 673174
rect 275514 672854 276134 672938
rect 275514 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 276134 672854
rect 275514 637174 276134 672618
rect 275514 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 276134 637174
rect 275514 636854 276134 636938
rect 275514 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 276134 636854
rect 275514 601174 276134 636618
rect 275514 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 276134 601174
rect 275514 600854 276134 600938
rect 275514 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 276134 600854
rect 275514 565174 276134 600618
rect 275514 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 276134 565174
rect 275514 564854 276134 564938
rect 275514 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 276134 564854
rect 275514 529174 276134 564618
rect 275514 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 276134 529174
rect 275514 528854 276134 528938
rect 275514 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 276134 528854
rect 275514 493174 276134 528618
rect 275514 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 276134 493174
rect 275514 492854 276134 492938
rect 275514 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 276134 492854
rect 275514 485308 276134 492618
rect 279234 676894 279854 709082
rect 279234 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 279854 676894
rect 279234 676574 279854 676658
rect 279234 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 279854 676574
rect 279234 640894 279854 676338
rect 279234 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 279854 640894
rect 279234 640574 279854 640658
rect 279234 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 279854 640574
rect 279234 604894 279854 640338
rect 279234 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 279854 604894
rect 279234 604574 279854 604658
rect 279234 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 279854 604574
rect 279234 568894 279854 604338
rect 279234 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 279854 568894
rect 279234 568574 279854 568658
rect 279234 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 279854 568574
rect 279234 532894 279854 568338
rect 279234 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 279854 532894
rect 279234 532574 279854 532658
rect 279234 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 279854 532574
rect 279234 496894 279854 532338
rect 279234 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 279854 496894
rect 279234 496574 279854 496658
rect 279234 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 279854 496574
rect 276243 485892 276309 485893
rect 276243 485828 276244 485892
rect 276308 485828 276309 485892
rect 276243 485827 276309 485828
rect 273483 484124 273549 484125
rect 273483 484060 273484 484124
rect 273548 484060 273549 484124
rect 273483 484059 273549 484060
rect 273486 483850 273546 484059
rect 276246 483850 276306 485827
rect 279234 485308 279854 496338
rect 282954 680614 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 282954 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 283574 680614
rect 282954 680294 283574 680378
rect 282954 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 283574 680294
rect 282954 644614 283574 680058
rect 282954 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 283574 644614
rect 282954 644294 283574 644378
rect 282954 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 283574 644294
rect 282954 608614 283574 644058
rect 282954 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 283574 608614
rect 282954 608294 283574 608378
rect 282954 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 283574 608294
rect 282954 572614 283574 608058
rect 282954 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 283574 572614
rect 282954 572294 283574 572378
rect 282954 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 283574 572294
rect 282954 536614 283574 572058
rect 282954 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 283574 536614
rect 282954 536294 283574 536378
rect 282954 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 283574 536294
rect 282954 500614 283574 536058
rect 282954 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 283574 500614
rect 282954 500294 283574 500378
rect 282954 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 283574 500294
rect 282954 485308 283574 500058
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 687454 290414 704282
rect 289794 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 290414 687454
rect 289794 687134 290414 687218
rect 289794 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 290414 687134
rect 289794 651454 290414 686898
rect 289794 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 290414 651454
rect 289794 651134 290414 651218
rect 289794 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 290414 651134
rect 289794 615454 290414 650898
rect 289794 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 290414 615454
rect 289794 615134 290414 615218
rect 289794 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 290414 615134
rect 289794 579454 290414 614898
rect 289794 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 290414 579454
rect 289794 579134 290414 579218
rect 289794 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 290414 579134
rect 289794 543454 290414 578898
rect 289794 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 290414 543454
rect 289794 543134 290414 543218
rect 289794 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 290414 543134
rect 289794 507454 290414 542898
rect 289794 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 290414 507454
rect 289794 507134 290414 507218
rect 289794 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 290414 507134
rect 283787 486708 283853 486709
rect 283787 486644 283788 486708
rect 283852 486644 283853 486708
rect 283787 486643 283853 486644
rect 278451 484804 278517 484805
rect 278451 484740 278452 484804
rect 278516 484740 278517 484804
rect 278451 484739 278517 484740
rect 268518 483790 268620 483850
rect 271094 483790 271204 483850
rect 273486 483790 273652 483850
rect 263528 483202 263588 483790
rect 266112 483202 266172 483790
rect 268560 483202 268620 483790
rect 271144 483202 271204 483790
rect 273592 483202 273652 483790
rect 276176 483790 276306 483850
rect 278454 483850 278514 484739
rect 280933 483852 280999 483853
rect 278454 483790 278548 483850
rect 276176 483202 276236 483790
rect 278488 483202 278548 483790
rect 280933 483788 280934 483852
rect 280998 483788 280999 483852
rect 283790 483850 283850 486643
rect 288571 486572 288637 486573
rect 288571 486508 288572 486572
rect 288636 486508 288637 486572
rect 288571 486507 288637 486508
rect 288574 483850 288634 486507
rect 289794 485308 290414 506898
rect 293514 691174 294134 706202
rect 293514 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 294134 691174
rect 293514 690854 294134 690938
rect 293514 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 294134 690854
rect 293514 655174 294134 690618
rect 293514 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 294134 655174
rect 293514 654854 294134 654938
rect 293514 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 294134 654854
rect 293514 619174 294134 654618
rect 293514 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 294134 619174
rect 293514 618854 294134 618938
rect 293514 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 294134 618854
rect 293514 583174 294134 618618
rect 293514 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 294134 583174
rect 293514 582854 294134 582938
rect 293514 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 294134 582854
rect 293514 547174 294134 582618
rect 293514 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 294134 547174
rect 293514 546854 294134 546938
rect 293514 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 294134 546854
rect 293514 511174 294134 546618
rect 293514 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 294134 511174
rect 293514 510854 294134 510938
rect 293514 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 294134 510854
rect 293514 485308 294134 510618
rect 297234 694894 297854 708122
rect 297234 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 297854 694894
rect 297234 694574 297854 694658
rect 297234 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 297854 694574
rect 297234 658894 297854 694338
rect 297234 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 297854 658894
rect 297234 658574 297854 658658
rect 297234 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 297854 658574
rect 297234 622894 297854 658338
rect 297234 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 297854 622894
rect 297234 622574 297854 622658
rect 297234 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 297854 622574
rect 297234 586894 297854 622338
rect 297234 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 297854 586894
rect 297234 586574 297854 586658
rect 297234 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 297854 586574
rect 297234 550894 297854 586338
rect 297234 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 297854 550894
rect 297234 550574 297854 550658
rect 297234 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 297854 550574
rect 297234 514894 297854 550338
rect 297234 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 297854 514894
rect 297234 514574 297854 514658
rect 297234 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 297854 514574
rect 297234 485308 297854 514338
rect 300954 698614 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 300954 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 301574 698614
rect 300954 698294 301574 698378
rect 300954 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 301574 698294
rect 300954 662614 301574 698058
rect 300954 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 301574 662614
rect 300954 662294 301574 662378
rect 300954 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 301574 662294
rect 300954 626614 301574 662058
rect 300954 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 301574 626614
rect 300954 626294 301574 626378
rect 300954 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 301574 626294
rect 300954 590614 301574 626058
rect 300954 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 301574 590614
rect 300954 590294 301574 590378
rect 300954 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 301574 590294
rect 300954 554614 301574 590058
rect 300954 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 301574 554614
rect 300954 554294 301574 554378
rect 300954 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 301574 554294
rect 300954 518614 301574 554058
rect 300954 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 301574 518614
rect 300954 518294 301574 518378
rect 300954 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 301574 518294
rect 300954 485308 301574 518058
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 669454 308414 705242
rect 307794 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 308414 669454
rect 307794 669134 308414 669218
rect 307794 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 308414 669134
rect 307794 633454 308414 668898
rect 307794 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 308414 633454
rect 307794 633134 308414 633218
rect 307794 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 308414 633134
rect 307794 597454 308414 632898
rect 307794 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 308414 597454
rect 307794 597134 308414 597218
rect 307794 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 308414 597134
rect 307794 561454 308414 596898
rect 307794 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 308414 561454
rect 307794 561134 308414 561218
rect 307794 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 308414 561134
rect 307794 525454 308414 560898
rect 307794 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 308414 525454
rect 307794 525134 308414 525218
rect 307794 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 308414 525134
rect 307794 489454 308414 524898
rect 307794 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 308414 489454
rect 307794 489134 308414 489218
rect 307794 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 308414 489134
rect 305867 486436 305933 486437
rect 305867 486372 305868 486436
rect 305932 486372 305933 486436
rect 305867 486371 305933 486372
rect 303475 485892 303541 485893
rect 303475 485828 303476 485892
rect 303540 485828 303541 485892
rect 303475 485827 303541 485828
rect 295931 485076 295997 485077
rect 295931 485012 295932 485076
rect 295996 485012 295997 485076
rect 295931 485011 295997 485012
rect 301083 485076 301149 485077
rect 301083 485012 301084 485076
rect 301148 485012 301149 485076
rect 301083 485011 301149 485012
rect 295934 483850 295994 485011
rect 298507 484532 298573 484533
rect 298507 484468 298508 484532
rect 298572 484468 298573 484532
rect 298507 484467 298573 484468
rect 280933 483787 280999 483788
rect 283656 483790 283850 483850
rect 288552 483790 288634 483850
rect 295896 483790 295994 483850
rect 298510 483850 298570 484467
rect 301086 483850 301146 485011
rect 298510 483790 298676 483850
rect 280936 483202 280996 483787
rect 283656 483202 283716 483790
rect 286101 483716 286167 483717
rect 286101 483652 286102 483716
rect 286166 483652 286167 483716
rect 286101 483651 286167 483652
rect 286104 483202 286164 483651
rect 288552 483202 288612 483790
rect 290997 483580 291063 483581
rect 290997 483516 290998 483580
rect 291062 483516 291063 483580
rect 290997 483515 291063 483516
rect 291000 483202 291060 483515
rect 293581 483444 293647 483445
rect 293581 483380 293582 483444
rect 293646 483380 293647 483444
rect 293581 483379 293647 483380
rect 293584 483202 293644 483379
rect 295896 483202 295956 483790
rect 298616 483202 298676 483790
rect 301064 483790 301146 483850
rect 303478 483850 303538 485827
rect 305870 483850 305930 486371
rect 307794 485308 308414 488898
rect 311514 673174 312134 707162
rect 311514 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 312134 673174
rect 311514 672854 312134 672938
rect 311514 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 312134 672854
rect 311514 637174 312134 672618
rect 311514 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 312134 637174
rect 311514 636854 312134 636938
rect 311514 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 312134 636854
rect 311514 601174 312134 636618
rect 311514 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 312134 601174
rect 311514 600854 312134 600938
rect 311514 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 312134 600854
rect 311514 565174 312134 600618
rect 311514 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 312134 565174
rect 311514 564854 312134 564938
rect 311514 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 312134 564854
rect 311514 529174 312134 564618
rect 311514 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 312134 529174
rect 311514 528854 312134 528938
rect 311514 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 312134 528854
rect 311514 493174 312134 528618
rect 311514 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 312134 493174
rect 311514 492854 312134 492938
rect 311514 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 312134 492854
rect 311514 485308 312134 492618
rect 315234 676894 315854 709082
rect 315234 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 315854 676894
rect 315234 676574 315854 676658
rect 315234 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 315854 676574
rect 315234 640894 315854 676338
rect 315234 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 315854 640894
rect 315234 640574 315854 640658
rect 315234 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 315854 640574
rect 315234 604894 315854 640338
rect 315234 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 315854 604894
rect 315234 604574 315854 604658
rect 315234 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 315854 604574
rect 315234 568894 315854 604338
rect 315234 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 315854 568894
rect 315234 568574 315854 568658
rect 315234 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 315854 568574
rect 315234 532894 315854 568338
rect 315234 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 315854 532894
rect 315234 532574 315854 532658
rect 315234 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 315854 532574
rect 315234 496894 315854 532338
rect 315234 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 315854 496894
rect 315234 496574 315854 496658
rect 315234 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 315854 496574
rect 313595 486300 313661 486301
rect 313595 486236 313596 486300
rect 313660 486236 313661 486300
rect 313595 486235 313661 486236
rect 308259 485212 308325 485213
rect 308259 485148 308260 485212
rect 308324 485148 308325 485212
rect 308259 485147 308325 485148
rect 308262 483850 308322 485147
rect 311019 484668 311085 484669
rect 311019 484604 311020 484668
rect 311084 484604 311085 484668
rect 311019 484603 311085 484604
rect 311022 483850 311082 484603
rect 313598 483850 313658 486235
rect 315234 485308 315854 496338
rect 318954 680614 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 318954 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 319574 680614
rect 318954 680294 319574 680378
rect 318954 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 319574 680294
rect 318954 644614 319574 680058
rect 318954 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 319574 644614
rect 318954 644294 319574 644378
rect 318954 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 319574 644294
rect 318954 608614 319574 644058
rect 318954 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 319574 608614
rect 318954 608294 319574 608378
rect 318954 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 319574 608294
rect 318954 572614 319574 608058
rect 318954 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 319574 572614
rect 318954 572294 319574 572378
rect 318954 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 319574 572294
rect 318954 536614 319574 572058
rect 318954 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 319574 536614
rect 318954 536294 319574 536378
rect 318954 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 319574 536294
rect 318954 500614 319574 536058
rect 318954 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 319574 500614
rect 318954 500294 319574 500378
rect 318954 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 319574 500294
rect 318379 486164 318445 486165
rect 318379 486100 318380 486164
rect 318444 486100 318445 486164
rect 318379 486099 318445 486100
rect 316171 483852 316237 483853
rect 316171 483850 316172 483852
rect 303478 483790 303572 483850
rect 305870 483790 306020 483850
rect 308262 483790 308468 483850
rect 301064 483202 301124 483790
rect 303512 483202 303572 483790
rect 305960 483202 306020 483790
rect 308408 483202 308468 483790
rect 310992 483790 311082 483850
rect 313576 483790 313658 483850
rect 316024 483790 316172 483850
rect 310992 483202 311052 483790
rect 313576 483202 313636 483790
rect 316024 483202 316084 483790
rect 316171 483788 316172 483790
rect 316236 483788 316237 483852
rect 318382 483850 318442 486099
rect 318954 485308 319574 500058
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 687454 326414 704282
rect 325794 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 326414 687454
rect 325794 687134 326414 687218
rect 325794 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 326414 687134
rect 325794 651454 326414 686898
rect 325794 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 326414 651454
rect 325794 651134 326414 651218
rect 325794 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 326414 651134
rect 325794 615454 326414 650898
rect 325794 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 326414 615454
rect 325794 615134 326414 615218
rect 325794 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 326414 615134
rect 325794 579454 326414 614898
rect 325794 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 326414 579454
rect 325794 579134 326414 579218
rect 325794 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 326414 579134
rect 325794 543454 326414 578898
rect 325794 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 326414 543454
rect 325794 543134 326414 543218
rect 325794 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 326414 543134
rect 325794 507454 326414 542898
rect 325794 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 326414 507454
rect 325794 507134 326414 507218
rect 325794 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 326414 507134
rect 323347 486028 323413 486029
rect 323347 485964 323348 486028
rect 323412 485964 323413 486028
rect 323347 485963 323413 485964
rect 323350 483850 323410 485963
rect 325794 485308 326414 506898
rect 329514 691174 330134 706202
rect 329514 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 330134 691174
rect 329514 690854 330134 690938
rect 329514 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 330134 690854
rect 329514 655174 330134 690618
rect 329514 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 330134 655174
rect 329514 654854 330134 654938
rect 329514 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 330134 654854
rect 329514 619174 330134 654618
rect 329514 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 330134 619174
rect 329514 618854 330134 618938
rect 329514 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 330134 618854
rect 329514 583174 330134 618618
rect 329514 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 330134 583174
rect 329514 582854 330134 582938
rect 329514 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 330134 582854
rect 329514 547174 330134 582618
rect 329514 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 330134 547174
rect 329514 546854 330134 546938
rect 329514 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 330134 546854
rect 329514 511174 330134 546618
rect 329514 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 330134 511174
rect 329514 510854 330134 510938
rect 329514 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 330134 510854
rect 326659 486980 326725 486981
rect 326659 486916 326660 486980
rect 326724 486916 326725 486980
rect 326659 486915 326725 486916
rect 326662 483850 326722 486915
rect 329514 485308 330134 510618
rect 333234 694894 333854 708122
rect 333234 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 333854 694894
rect 333234 694574 333854 694658
rect 333234 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 333854 694574
rect 333234 658894 333854 694338
rect 333234 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 333854 658894
rect 333234 658574 333854 658658
rect 333234 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 333854 658574
rect 333234 622894 333854 658338
rect 333234 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 333854 622894
rect 333234 622574 333854 622658
rect 333234 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 333854 622574
rect 333234 586894 333854 622338
rect 333234 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 333854 586894
rect 333234 586574 333854 586658
rect 333234 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 333854 586574
rect 333234 550894 333854 586338
rect 333234 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 333854 550894
rect 333234 550574 333854 550658
rect 333234 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 333854 550574
rect 333234 514894 333854 550338
rect 333234 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 333854 514894
rect 333234 514574 333854 514658
rect 333234 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 333854 514574
rect 333234 485308 333854 514338
rect 336954 698614 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 336954 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 337574 698614
rect 336954 698294 337574 698378
rect 336954 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 337574 698294
rect 336954 662614 337574 698058
rect 336954 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 337574 662614
rect 336954 662294 337574 662378
rect 336954 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 337574 662294
rect 336954 626614 337574 662058
rect 336954 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 337574 626614
rect 336954 626294 337574 626378
rect 336954 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 337574 626294
rect 336954 590614 337574 626058
rect 336954 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 337574 590614
rect 336954 590294 337574 590378
rect 336954 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 337574 590294
rect 336954 554614 337574 590058
rect 336954 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 337574 554614
rect 336954 554294 337574 554378
rect 336954 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 337574 554294
rect 336954 518614 337574 554058
rect 336954 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 337574 518614
rect 336954 518294 337574 518378
rect 336954 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 337574 518294
rect 336954 485308 337574 518058
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 669454 344414 705242
rect 343794 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 344414 669454
rect 343794 669134 344414 669218
rect 343794 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 344414 669134
rect 343794 633454 344414 668898
rect 343794 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 344414 633454
rect 343794 633134 344414 633218
rect 343794 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 344414 633134
rect 343794 597454 344414 632898
rect 343794 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 344414 597454
rect 343794 597134 344414 597218
rect 343794 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 344414 597134
rect 343794 561454 344414 596898
rect 343794 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 344414 561454
rect 343794 561134 344414 561218
rect 343794 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 344414 561134
rect 343794 525454 344414 560898
rect 343794 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 344414 525454
rect 343794 525134 344414 525218
rect 343794 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 344414 525134
rect 343794 489454 344414 524898
rect 343794 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 344414 489454
rect 343794 489134 344414 489218
rect 343794 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 344414 489134
rect 339723 486436 339789 486437
rect 339723 486372 339724 486436
rect 339788 486372 339789 486436
rect 339723 486371 339789 486372
rect 338435 485892 338501 485893
rect 338435 485828 338436 485892
rect 338500 485828 338501 485892
rect 338435 485827 338501 485828
rect 318382 483790 318532 483850
rect 323350 483790 323428 483850
rect 316171 483787 316237 483788
rect 318472 483202 318532 483790
rect 321053 483444 321119 483445
rect 321053 483380 321054 483444
rect 321118 483380 321119 483444
rect 321053 483379 321119 483380
rect 321056 483202 321116 483379
rect 323368 483202 323428 483790
rect 326088 483790 326722 483850
rect 338438 483850 338498 485827
rect 339726 483850 339786 486371
rect 343794 485308 344414 488898
rect 347514 673174 348134 707162
rect 347514 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 348134 673174
rect 347514 672854 348134 672938
rect 347514 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 348134 672854
rect 347514 637174 348134 672618
rect 347514 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 348134 637174
rect 347514 636854 348134 636938
rect 347514 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 348134 636854
rect 347514 601174 348134 636618
rect 347514 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 348134 601174
rect 347514 600854 348134 600938
rect 347514 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 348134 600854
rect 347514 565174 348134 600618
rect 347514 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 348134 565174
rect 347514 564854 348134 564938
rect 347514 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 348134 564854
rect 347514 529174 348134 564618
rect 347514 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 348134 529174
rect 347514 528854 348134 528938
rect 347514 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 348134 528854
rect 347514 493174 348134 528618
rect 347514 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 348134 493174
rect 347514 492854 348134 492938
rect 347514 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 348134 492854
rect 347514 485308 348134 492618
rect 351234 676894 351854 709082
rect 351234 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 351854 676894
rect 351234 676574 351854 676658
rect 351234 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 351854 676574
rect 351234 640894 351854 676338
rect 351234 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 351854 640894
rect 351234 640574 351854 640658
rect 351234 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 351854 640574
rect 351234 604894 351854 640338
rect 351234 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 351854 604894
rect 351234 604574 351854 604658
rect 351234 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 351854 604574
rect 351234 568894 351854 604338
rect 351234 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 351854 568894
rect 351234 568574 351854 568658
rect 351234 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 351854 568574
rect 351234 532894 351854 568338
rect 351234 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 351854 532894
rect 351234 532574 351854 532658
rect 351234 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 351854 532574
rect 351234 496894 351854 532338
rect 351234 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 351854 496894
rect 351234 496574 351854 496658
rect 351234 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 351854 496574
rect 350763 486436 350829 486437
rect 350763 486372 350764 486436
rect 350828 486372 350829 486436
rect 350763 486371 350829 486372
rect 338438 483790 338524 483850
rect 326088 483202 326148 483790
rect 338464 483202 338524 483790
rect 339688 483790 339786 483850
rect 350766 483850 350826 486371
rect 351234 485308 351854 496338
rect 354954 680614 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 354954 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 355574 680614
rect 354954 680294 355574 680378
rect 354954 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 355574 680294
rect 354954 644614 355574 680058
rect 354954 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 355574 644614
rect 354954 644294 355574 644378
rect 354954 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 355574 644294
rect 354954 608614 355574 644058
rect 354954 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 355574 608614
rect 354954 608294 355574 608378
rect 354954 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 355574 608294
rect 354954 572614 355574 608058
rect 354954 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 355574 572614
rect 354954 572294 355574 572378
rect 354954 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 355574 572294
rect 354954 536614 355574 572058
rect 354954 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 355574 536614
rect 354954 536294 355574 536378
rect 354954 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 355574 536294
rect 354954 500614 355574 536058
rect 354954 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 355574 500614
rect 354954 500294 355574 500378
rect 354954 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 355574 500294
rect 354954 485308 355574 500058
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 687454 362414 704282
rect 361794 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 362414 687454
rect 361794 687134 362414 687218
rect 361794 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 362414 687134
rect 361794 651454 362414 686898
rect 361794 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 362414 651454
rect 361794 651134 362414 651218
rect 361794 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 362414 651134
rect 361794 615454 362414 650898
rect 361794 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 362414 615454
rect 361794 615134 362414 615218
rect 361794 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 362414 615134
rect 361794 579454 362414 614898
rect 361794 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 362414 579454
rect 361794 579134 362414 579218
rect 361794 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 362414 579134
rect 361794 543454 362414 578898
rect 361794 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 362414 543454
rect 361794 543134 362414 543218
rect 361794 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 362414 543134
rect 361794 507454 362414 542898
rect 361794 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 362414 507454
rect 361794 507134 362414 507218
rect 361794 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 362414 507134
rect 350766 483790 350900 483850
rect 339688 483202 339748 483790
rect 350840 483202 350900 483790
rect 220952 471454 221300 471486
rect 220952 471218 221008 471454
rect 221244 471218 221300 471454
rect 220952 471134 221300 471218
rect 220952 470898 221008 471134
rect 221244 470898 221300 471134
rect 220952 470866 221300 470898
rect 355320 471454 355668 471486
rect 355320 471218 355376 471454
rect 355612 471218 355668 471454
rect 355320 471134 355668 471218
rect 355320 470898 355376 471134
rect 355612 470898 355668 471134
rect 355320 470866 355668 470898
rect 361794 471454 362414 506898
rect 361794 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 362414 471454
rect 361794 471134 362414 471218
rect 361794 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 362414 471134
rect 220272 453454 220620 453486
rect 220272 453218 220328 453454
rect 220564 453218 220620 453454
rect 220272 453134 220620 453218
rect 220272 452898 220328 453134
rect 220564 452898 220620 453134
rect 220272 452866 220620 452898
rect 356000 453454 356348 453486
rect 356000 453218 356056 453454
rect 356292 453218 356348 453454
rect 356000 453134 356348 453218
rect 356000 452898 356056 453134
rect 356292 452898 356348 453134
rect 356000 452866 356348 452898
rect 220952 435454 221300 435486
rect 220952 435218 221008 435454
rect 221244 435218 221300 435454
rect 220952 435134 221300 435218
rect 220952 434898 221008 435134
rect 221244 434898 221300 435134
rect 220952 434866 221300 434898
rect 355320 435454 355668 435486
rect 355320 435218 355376 435454
rect 355612 435218 355668 435454
rect 355320 435134 355668 435218
rect 355320 434898 355376 435134
rect 355612 434898 355668 435134
rect 355320 434866 355668 434898
rect 361794 435454 362414 470898
rect 361794 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 362414 435454
rect 361794 435134 362414 435218
rect 361794 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 362414 435134
rect 220272 417454 220620 417486
rect 220272 417218 220328 417454
rect 220564 417218 220620 417454
rect 220272 417134 220620 417218
rect 220272 416898 220328 417134
rect 220564 416898 220620 417134
rect 220272 416866 220620 416898
rect 356000 417454 356348 417486
rect 356000 417218 356056 417454
rect 356292 417218 356348 417454
rect 356000 417134 356348 417218
rect 356000 416898 356056 417134
rect 356292 416898 356348 417134
rect 356000 416866 356348 416898
rect 223619 399532 223685 399533
rect 223619 399468 223620 399532
rect 223684 399468 223685 399532
rect 236056 399530 236116 400106
rect 237144 399530 237204 400106
rect 238232 399530 238292 400106
rect 239592 399530 239652 400106
rect 223619 399467 223685 399468
rect 235950 399470 236116 399530
rect 237054 399470 237204 399530
rect 238158 399470 238292 399530
rect 239262 399470 239652 399530
rect 240544 399530 240604 400106
rect 241768 399530 241828 400106
rect 243128 399530 243188 400106
rect 240544 399470 240610 399530
rect 219939 398172 220005 398173
rect 219939 398108 219940 398172
rect 220004 398108 220005 398172
rect 219939 398107 220005 398108
rect 219755 398036 219821 398037
rect 219755 397972 219756 398036
rect 219820 397972 219821 398036
rect 219755 397971 219821 397972
rect 219387 393412 219453 393413
rect 219387 393348 219388 393412
rect 219452 393348 219453 393412
rect 219387 393347 219453 393348
rect 219203 392868 219269 392869
rect 219203 392804 219204 392868
rect 219268 392804 219269 392868
rect 219203 392803 219269 392804
rect 219390 392730 219450 393347
rect 219206 392670 219450 392730
rect 219206 383890 219266 392670
rect 219206 383830 219450 383890
rect 219203 383756 219269 383757
rect 219203 383692 219204 383756
rect 219268 383692 219269 383756
rect 219203 383691 219269 383692
rect 219206 344589 219266 383691
rect 219390 383621 219450 383830
rect 219387 383620 219453 383621
rect 219387 383556 219388 383620
rect 219452 383556 219453 383620
rect 219387 383555 219453 383556
rect 219387 374236 219453 374237
rect 219387 374172 219388 374236
rect 219452 374172 219453 374236
rect 219387 374171 219453 374172
rect 219390 373965 219450 374171
rect 219387 373964 219453 373965
rect 219387 373900 219388 373964
rect 219452 373900 219453 373964
rect 219387 373899 219453 373900
rect 221514 367174 222134 398000
rect 221514 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 222134 367174
rect 221514 366854 222134 366938
rect 221514 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 222134 366854
rect 219387 364444 219453 364445
rect 219387 364380 219388 364444
rect 219452 364380 219453 364444
rect 219387 364379 219453 364380
rect 219390 364309 219450 364379
rect 219387 364308 219453 364309
rect 219387 364244 219388 364308
rect 219452 364244 219453 364308
rect 219387 364243 219453 364244
rect 219387 354788 219453 354789
rect 219387 354724 219388 354788
rect 219452 354724 219453 354788
rect 219387 354723 219453 354724
rect 219390 354653 219450 354723
rect 219387 354652 219453 354653
rect 219387 354588 219388 354652
rect 219452 354588 219453 354652
rect 219387 354587 219453 354588
rect 219387 345132 219453 345133
rect 219387 345068 219388 345132
rect 219452 345068 219453 345132
rect 219387 345067 219453 345068
rect 219203 344588 219269 344589
rect 219203 344524 219204 344588
rect 219268 344524 219269 344588
rect 219203 344523 219269 344524
rect 219390 344450 219450 345067
rect 219206 344390 219450 344450
rect 219206 335610 219266 344390
rect 219206 335550 219450 335610
rect 219203 335476 219269 335477
rect 219203 335412 219204 335476
rect 219268 335412 219269 335476
rect 219203 335411 219269 335412
rect 219206 335069 219266 335411
rect 219203 335068 219269 335069
rect 219203 335004 219204 335068
rect 219268 335004 219269 335068
rect 219203 335003 219269 335004
rect 219390 334930 219450 335550
rect 219206 334870 219450 334930
rect 219206 326090 219266 334870
rect 221514 331174 222134 366618
rect 221514 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 222134 331174
rect 221514 330854 222134 330938
rect 221514 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 222134 330854
rect 219206 326030 219450 326090
rect 219203 325956 219269 325957
rect 219203 325892 219204 325956
rect 219268 325892 219269 325956
rect 219203 325891 219269 325892
rect 219206 248029 219266 325891
rect 219390 325685 219450 326030
rect 219387 325684 219453 325685
rect 219387 325620 219388 325684
rect 219452 325620 219453 325684
rect 219387 325619 219453 325620
rect 219387 316300 219453 316301
rect 219387 316236 219388 316300
rect 219452 316236 219453 316300
rect 219387 316235 219453 316236
rect 219390 316029 219450 316235
rect 219387 316028 219453 316029
rect 219387 315964 219388 316028
rect 219452 315964 219453 316028
rect 219387 315963 219453 315964
rect 219387 306508 219453 306509
rect 219387 306444 219388 306508
rect 219452 306444 219453 306508
rect 219387 306443 219453 306444
rect 219390 306373 219450 306443
rect 219387 306372 219453 306373
rect 219387 306308 219388 306372
rect 219452 306308 219453 306372
rect 219387 306307 219453 306308
rect 219387 296852 219453 296853
rect 219387 296788 219388 296852
rect 219452 296788 219453 296852
rect 219387 296787 219453 296788
rect 219390 296717 219450 296787
rect 219387 296716 219453 296717
rect 219387 296652 219388 296716
rect 219452 296652 219453 296716
rect 219387 296651 219453 296652
rect 221514 295174 222134 330618
rect 221514 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 222134 295174
rect 221514 294854 222134 294938
rect 221514 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 222134 294854
rect 219387 287196 219453 287197
rect 219387 287132 219388 287196
rect 219452 287132 219453 287196
rect 219387 287131 219453 287132
rect 219390 287061 219450 287131
rect 219387 287060 219453 287061
rect 219387 286996 219388 287060
rect 219452 286996 219453 287060
rect 219387 286995 219453 286996
rect 219387 277540 219453 277541
rect 219387 277476 219388 277540
rect 219452 277476 219453 277540
rect 219387 277475 219453 277476
rect 219390 277405 219450 277475
rect 219387 277404 219453 277405
rect 219387 277340 219388 277404
rect 219452 277340 219453 277404
rect 219387 277339 219453 277340
rect 219387 267884 219453 267885
rect 219387 267820 219388 267884
rect 219452 267820 219453 267884
rect 219387 267819 219453 267820
rect 219390 267749 219450 267819
rect 219387 267748 219453 267749
rect 219387 267684 219388 267748
rect 219452 267684 219453 267748
rect 219387 267683 219453 267684
rect 221514 259174 222134 294618
rect 221514 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 222134 259174
rect 221514 258854 222134 258938
rect 221514 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 222134 258854
rect 219387 258364 219453 258365
rect 219387 258300 219388 258364
rect 219452 258300 219453 258364
rect 219387 258299 219453 258300
rect 219390 257957 219450 258299
rect 219387 257956 219453 257957
rect 219387 257892 219388 257956
rect 219452 257892 219453 257956
rect 219387 257891 219453 257892
rect 219387 248436 219453 248437
rect 219387 248372 219388 248436
rect 219452 248372 219453 248436
rect 219387 248371 219453 248372
rect 219203 248028 219269 248029
rect 219203 247964 219204 248028
rect 219268 247964 219269 248028
rect 219203 247963 219269 247964
rect 219390 247890 219450 248371
rect 219206 247830 219450 247890
rect 219206 235381 219266 247830
rect 219387 238916 219453 238917
rect 219387 238852 219388 238916
rect 219452 238852 219453 238916
rect 219387 238851 219453 238852
rect 219390 238237 219450 238851
rect 219387 238236 219453 238237
rect 219387 238172 219388 238236
rect 219452 238172 219453 238236
rect 219387 238171 219453 238172
rect 219203 235380 219269 235381
rect 219203 235316 219204 235380
rect 219268 235316 219269 235380
rect 219203 235315 219269 235316
rect 219203 235108 219269 235109
rect 219203 235044 219204 235108
rect 219268 235044 219269 235108
rect 219203 235043 219269 235044
rect 219206 230893 219266 235043
rect 219203 230892 219269 230893
rect 219203 230828 219204 230892
rect 219268 230828 219269 230892
rect 219203 230827 219269 230828
rect 221514 228924 222134 258618
rect 219019 228852 219085 228853
rect 219019 228788 219020 228852
rect 219084 228788 219085 228852
rect 219019 228787 219085 228788
rect 60595 226676 60661 226677
rect 60595 226612 60596 226676
rect 60660 226612 60661 226676
rect 60595 226611 60661 226612
rect 60598 225997 60658 226611
rect 60779 226268 60845 226269
rect 60779 226204 60780 226268
rect 60844 226204 60845 226268
rect 60779 226203 60845 226204
rect 223435 226268 223501 226269
rect 223435 226204 223436 226268
rect 223500 226204 223501 226268
rect 223435 226203 223501 226204
rect 60595 225996 60661 225997
rect 60595 225932 60596 225996
rect 60660 225932 60661 225996
rect 60595 225931 60661 225932
rect 60782 225861 60842 226203
rect 60779 225860 60845 225861
rect 60779 225796 60780 225860
rect 60844 225796 60845 225860
rect 60779 225795 60845 225796
rect 223438 225725 223498 226203
rect 223435 225724 223501 225725
rect 223435 225660 223436 225724
rect 223500 225660 223501 225724
rect 223435 225659 223501 225660
rect 64208 219454 64528 219486
rect 64208 219218 64250 219454
rect 64486 219218 64528 219454
rect 64208 219134 64528 219218
rect 64208 218898 64250 219134
rect 64486 218898 64528 219134
rect 64208 218866 64528 218898
rect 94928 219454 95248 219486
rect 94928 219218 94970 219454
rect 95206 219218 95248 219454
rect 94928 219134 95248 219218
rect 94928 218898 94970 219134
rect 95206 218898 95248 219134
rect 94928 218866 95248 218898
rect 125648 219454 125968 219486
rect 125648 219218 125690 219454
rect 125926 219218 125968 219454
rect 125648 219134 125968 219218
rect 125648 218898 125690 219134
rect 125926 218898 125968 219134
rect 125648 218866 125968 218898
rect 156368 219454 156688 219486
rect 156368 219218 156410 219454
rect 156646 219218 156688 219454
rect 156368 219134 156688 219218
rect 156368 218898 156410 219134
rect 156646 218898 156688 219134
rect 156368 218866 156688 218898
rect 187088 219454 187408 219486
rect 187088 219218 187130 219454
rect 187366 219218 187408 219454
rect 187088 219134 187408 219218
rect 187088 218898 187130 219134
rect 187366 218898 187408 219134
rect 187088 218866 187408 218898
rect 217808 219454 218128 219486
rect 217808 219218 217850 219454
rect 218086 219218 218128 219454
rect 217808 219134 218128 219218
rect 217808 218898 217850 219134
rect 218086 218898 218128 219134
rect 217808 218866 218128 218898
rect 55794 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 56414 201454
rect 55794 201134 56414 201218
rect 55794 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 56414 201134
rect 55794 165454 56414 200898
rect 79568 201454 79888 201486
rect 79568 201218 79610 201454
rect 79846 201218 79888 201454
rect 79568 201134 79888 201218
rect 79568 200898 79610 201134
rect 79846 200898 79888 201134
rect 79568 200866 79888 200898
rect 110288 201454 110608 201486
rect 110288 201218 110330 201454
rect 110566 201218 110608 201454
rect 110288 201134 110608 201218
rect 110288 200898 110330 201134
rect 110566 200898 110608 201134
rect 110288 200866 110608 200898
rect 141008 201454 141328 201486
rect 141008 201218 141050 201454
rect 141286 201218 141328 201454
rect 141008 201134 141328 201218
rect 141008 200898 141050 201134
rect 141286 200898 141328 201134
rect 141008 200866 141328 200898
rect 171728 201454 172048 201486
rect 171728 201218 171770 201454
rect 172006 201218 172048 201454
rect 171728 201134 172048 201218
rect 171728 200898 171770 201134
rect 172006 200898 172048 201134
rect 171728 200866 172048 200898
rect 202448 201454 202768 201486
rect 202448 201218 202490 201454
rect 202726 201218 202768 201454
rect 202448 201134 202768 201218
rect 202448 200898 202490 201134
rect 202726 200898 202768 201134
rect 202448 200866 202768 200898
rect 64208 183454 64528 183486
rect 64208 183218 64250 183454
rect 64486 183218 64528 183454
rect 64208 183134 64528 183218
rect 64208 182898 64250 183134
rect 64486 182898 64528 183134
rect 64208 182866 64528 182898
rect 94928 183454 95248 183486
rect 94928 183218 94970 183454
rect 95206 183218 95248 183454
rect 94928 183134 95248 183218
rect 94928 182898 94970 183134
rect 95206 182898 95248 183134
rect 94928 182866 95248 182898
rect 125648 183454 125968 183486
rect 125648 183218 125690 183454
rect 125926 183218 125968 183454
rect 125648 183134 125968 183218
rect 125648 182898 125690 183134
rect 125926 182898 125968 183134
rect 125648 182866 125968 182898
rect 156368 183454 156688 183486
rect 156368 183218 156410 183454
rect 156646 183218 156688 183454
rect 156368 183134 156688 183218
rect 156368 182898 156410 183134
rect 156646 182898 156688 183134
rect 156368 182866 156688 182898
rect 187088 183454 187408 183486
rect 187088 183218 187130 183454
rect 187366 183218 187408 183454
rect 187088 183134 187408 183218
rect 187088 182898 187130 183134
rect 187366 182898 187408 183134
rect 187088 182866 187408 182898
rect 217808 183454 218128 183486
rect 217808 183218 217850 183454
rect 218086 183218 218128 183454
rect 217808 183134 218128 183218
rect 217808 182898 217850 183134
rect 218086 182898 218128 183134
rect 217808 182866 218128 182898
rect 55794 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 56414 165454
rect 55794 165134 56414 165218
rect 55794 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 56414 165134
rect 55794 129454 56414 164898
rect 79568 165454 79888 165486
rect 79568 165218 79610 165454
rect 79846 165218 79888 165454
rect 79568 165134 79888 165218
rect 79568 164898 79610 165134
rect 79846 164898 79888 165134
rect 79568 164866 79888 164898
rect 110288 165454 110608 165486
rect 110288 165218 110330 165454
rect 110566 165218 110608 165454
rect 110288 165134 110608 165218
rect 110288 164898 110330 165134
rect 110566 164898 110608 165134
rect 110288 164866 110608 164898
rect 141008 165454 141328 165486
rect 141008 165218 141050 165454
rect 141286 165218 141328 165454
rect 141008 165134 141328 165218
rect 141008 164898 141050 165134
rect 141286 164898 141328 165134
rect 141008 164866 141328 164898
rect 171728 165454 172048 165486
rect 171728 165218 171770 165454
rect 172006 165218 172048 165454
rect 171728 165134 172048 165218
rect 171728 164898 171770 165134
rect 172006 164898 172048 165134
rect 171728 164866 172048 164898
rect 202448 165454 202768 165486
rect 202448 165218 202490 165454
rect 202726 165218 202768 165454
rect 202448 165134 202768 165218
rect 202448 164898 202490 165134
rect 202726 164898 202768 165134
rect 202448 164866 202768 164898
rect 64208 147454 64528 147486
rect 64208 147218 64250 147454
rect 64486 147218 64528 147454
rect 64208 147134 64528 147218
rect 64208 146898 64250 147134
rect 64486 146898 64528 147134
rect 64208 146866 64528 146898
rect 94928 147454 95248 147486
rect 94928 147218 94970 147454
rect 95206 147218 95248 147454
rect 94928 147134 95248 147218
rect 94928 146898 94970 147134
rect 95206 146898 95248 147134
rect 94928 146866 95248 146898
rect 125648 147454 125968 147486
rect 125648 147218 125690 147454
rect 125926 147218 125968 147454
rect 125648 147134 125968 147218
rect 125648 146898 125690 147134
rect 125926 146898 125968 147134
rect 125648 146866 125968 146898
rect 156368 147454 156688 147486
rect 156368 147218 156410 147454
rect 156646 147218 156688 147454
rect 156368 147134 156688 147218
rect 156368 146898 156410 147134
rect 156646 146898 156688 147134
rect 156368 146866 156688 146898
rect 187088 147454 187408 147486
rect 187088 147218 187130 147454
rect 187366 147218 187408 147454
rect 187088 147134 187408 147218
rect 187088 146898 187130 147134
rect 187366 146898 187408 147134
rect 187088 146866 187408 146898
rect 217808 147454 218128 147486
rect 217808 147218 217850 147454
rect 218086 147218 218128 147454
rect 217808 147134 218128 147218
rect 217808 146898 217850 147134
rect 218086 146898 218128 147134
rect 217808 146866 218128 146898
rect 55794 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 56414 129454
rect 55794 129134 56414 129218
rect 55794 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 56414 129134
rect 55794 93454 56414 128898
rect 79568 129454 79888 129486
rect 79568 129218 79610 129454
rect 79846 129218 79888 129454
rect 79568 129134 79888 129218
rect 79568 128898 79610 129134
rect 79846 128898 79888 129134
rect 79568 128866 79888 128898
rect 110288 129454 110608 129486
rect 110288 129218 110330 129454
rect 110566 129218 110608 129454
rect 110288 129134 110608 129218
rect 110288 128898 110330 129134
rect 110566 128898 110608 129134
rect 110288 128866 110608 128898
rect 141008 129454 141328 129486
rect 141008 129218 141050 129454
rect 141286 129218 141328 129454
rect 141008 129134 141328 129218
rect 141008 128898 141050 129134
rect 141286 128898 141328 129134
rect 141008 128866 141328 128898
rect 171728 129454 172048 129486
rect 171728 129218 171770 129454
rect 172006 129218 172048 129454
rect 171728 129134 172048 129218
rect 171728 128898 171770 129134
rect 172006 128898 172048 129134
rect 171728 128866 172048 128898
rect 202448 129454 202768 129486
rect 202448 129218 202490 129454
rect 202726 129218 202768 129454
rect 202448 129134 202768 129218
rect 202448 128898 202490 129134
rect 202726 128898 202768 129134
rect 202448 128866 202768 128898
rect 64208 111454 64528 111486
rect 64208 111218 64250 111454
rect 64486 111218 64528 111454
rect 64208 111134 64528 111218
rect 64208 110898 64250 111134
rect 64486 110898 64528 111134
rect 64208 110866 64528 110898
rect 94928 111454 95248 111486
rect 94928 111218 94970 111454
rect 95206 111218 95248 111454
rect 94928 111134 95248 111218
rect 94928 110898 94970 111134
rect 95206 110898 95248 111134
rect 94928 110866 95248 110898
rect 125648 111454 125968 111486
rect 125648 111218 125690 111454
rect 125926 111218 125968 111454
rect 125648 111134 125968 111218
rect 125648 110898 125690 111134
rect 125926 110898 125968 111134
rect 125648 110866 125968 110898
rect 156368 111454 156688 111486
rect 156368 111218 156410 111454
rect 156646 111218 156688 111454
rect 156368 111134 156688 111218
rect 156368 110898 156410 111134
rect 156646 110898 156688 111134
rect 156368 110866 156688 110898
rect 187088 111454 187408 111486
rect 187088 111218 187130 111454
rect 187366 111218 187408 111454
rect 187088 111134 187408 111218
rect 187088 110898 187130 111134
rect 187366 110898 187408 111134
rect 187088 110866 187408 110898
rect 217808 111454 218128 111486
rect 217808 111218 217850 111454
rect 218086 111218 218128 111454
rect 217808 111134 218128 111218
rect 217808 110898 217850 111134
rect 218086 110898 218128 111134
rect 217808 110866 218128 110898
rect 55794 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 56414 93454
rect 55794 93134 56414 93218
rect 55794 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 56414 93134
rect 55794 57454 56414 92898
rect 79568 93454 79888 93486
rect 79568 93218 79610 93454
rect 79846 93218 79888 93454
rect 79568 93134 79888 93218
rect 79568 92898 79610 93134
rect 79846 92898 79888 93134
rect 79568 92866 79888 92898
rect 110288 93454 110608 93486
rect 110288 93218 110330 93454
rect 110566 93218 110608 93454
rect 110288 93134 110608 93218
rect 110288 92898 110330 93134
rect 110566 92898 110608 93134
rect 110288 92866 110608 92898
rect 141008 93454 141328 93486
rect 141008 93218 141050 93454
rect 141286 93218 141328 93454
rect 141008 93134 141328 93218
rect 141008 92898 141050 93134
rect 141286 92898 141328 93134
rect 141008 92866 141328 92898
rect 171728 93454 172048 93486
rect 171728 93218 171770 93454
rect 172006 93218 172048 93454
rect 171728 93134 172048 93218
rect 171728 92898 171770 93134
rect 172006 92898 172048 93134
rect 171728 92866 172048 92898
rect 202448 93454 202768 93486
rect 202448 93218 202490 93454
rect 202726 93218 202768 93454
rect 202448 93134 202768 93218
rect 202448 92898 202490 93134
rect 202726 92898 202768 93134
rect 202448 92866 202768 92898
rect 64208 75454 64528 75486
rect 64208 75218 64250 75454
rect 64486 75218 64528 75454
rect 64208 75134 64528 75218
rect 64208 74898 64250 75134
rect 64486 74898 64528 75134
rect 64208 74866 64528 74898
rect 94928 75454 95248 75486
rect 94928 75218 94970 75454
rect 95206 75218 95248 75454
rect 94928 75134 95248 75218
rect 94928 74898 94970 75134
rect 95206 74898 95248 75134
rect 94928 74866 95248 74898
rect 125648 75454 125968 75486
rect 125648 75218 125690 75454
rect 125926 75218 125968 75454
rect 125648 75134 125968 75218
rect 125648 74898 125690 75134
rect 125926 74898 125968 75134
rect 125648 74866 125968 74898
rect 156368 75454 156688 75486
rect 156368 75218 156410 75454
rect 156646 75218 156688 75454
rect 156368 75134 156688 75218
rect 156368 74898 156410 75134
rect 156646 74898 156688 75134
rect 156368 74866 156688 74898
rect 187088 75454 187408 75486
rect 187088 75218 187130 75454
rect 187366 75218 187408 75454
rect 187088 75134 187408 75218
rect 187088 74898 187130 75134
rect 187366 74898 187408 75134
rect 187088 74866 187408 74898
rect 217808 75454 218128 75486
rect 217808 75218 217850 75454
rect 218086 75218 218128 75454
rect 217808 75134 218128 75218
rect 217808 74898 217850 75134
rect 218086 74898 218128 75134
rect 217808 74866 218128 74898
rect 223622 60349 223682 399467
rect 226379 398308 226445 398309
rect 226379 398244 226380 398308
rect 226444 398244 226445 398308
rect 226379 398243 226445 398244
rect 225234 370894 225854 398000
rect 225234 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 225854 370894
rect 225234 370574 225854 370658
rect 225234 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 225854 370574
rect 225234 334894 225854 370338
rect 225234 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 225854 334894
rect 225234 334574 225854 334658
rect 225234 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 225854 334574
rect 225234 298894 225854 334338
rect 225234 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 225854 298894
rect 225234 298574 225854 298658
rect 225234 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 225854 298574
rect 225234 262894 225854 298338
rect 225234 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 225854 262894
rect 225234 262574 225854 262658
rect 225234 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 225854 262574
rect 224726 232190 225154 232250
rect 224726 231709 224786 232190
rect 224907 231844 224973 231845
rect 224907 231780 224908 231844
rect 224972 231780 224973 231844
rect 224907 231779 224973 231780
rect 224723 231708 224789 231709
rect 224723 231644 224724 231708
rect 224788 231644 224789 231708
rect 224723 231643 224789 231644
rect 223987 231028 224053 231029
rect 223987 230964 223988 231028
rect 224052 230964 224053 231028
rect 223987 230963 224053 230964
rect 223803 230892 223869 230893
rect 223803 230828 223804 230892
rect 223868 230828 223869 230892
rect 223803 230827 223869 230828
rect 223619 60348 223685 60349
rect 223619 60284 223620 60348
rect 223684 60284 223685 60348
rect 223619 60283 223685 60284
rect 223806 59125 223866 230827
rect 223990 59125 224050 230963
rect 224171 228852 224237 228853
rect 224171 228788 224172 228852
rect 224236 228788 224237 228852
rect 224171 228787 224237 228788
rect 224174 59805 224234 228787
rect 224355 228716 224421 228717
rect 224355 228652 224356 228716
rect 224420 228652 224421 228716
rect 224355 228651 224421 228652
rect 224171 59804 224237 59805
rect 224171 59740 224172 59804
rect 224236 59740 224237 59804
rect 224171 59739 224237 59740
rect 224358 59125 224418 228651
rect 224910 70277 224970 231779
rect 224907 70276 224973 70277
rect 224907 70212 224908 70276
rect 224972 70212 224973 70276
rect 224907 70211 224973 70212
rect 224907 60756 224973 60757
rect 224907 60692 224908 60756
rect 224972 60692 224973 60756
rect 224907 60691 224973 60692
rect 223803 59124 223869 59125
rect 223803 59060 223804 59124
rect 223868 59060 223869 59124
rect 223803 59059 223869 59060
rect 223987 59124 224053 59125
rect 223987 59060 223988 59124
rect 224052 59060 224053 59124
rect 223987 59059 224053 59060
rect 224355 59124 224421 59125
rect 224355 59060 224356 59124
rect 224420 59060 224421 59124
rect 224355 59059 224421 59060
rect 55794 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 56414 57454
rect 55794 57134 56414 57218
rect 55794 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 56414 57134
rect 55794 21454 56414 56898
rect 55794 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 56414 21454
rect 55794 21134 56414 21218
rect 55794 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 56414 21134
rect 55794 -1306 56414 20898
rect 55794 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 56414 -1306
rect 55794 -1626 56414 -1542
rect 55794 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 56414 -1626
rect 55794 -1894 56414 -1862
rect 59514 25174 60134 58000
rect 59514 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 60134 25174
rect 59514 24854 60134 24938
rect 59514 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 60134 24854
rect 59514 -3226 60134 24618
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 28894 63854 58000
rect 63234 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 63854 28894
rect 63234 28574 63854 28658
rect 63234 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 63854 28574
rect 63234 -5146 63854 28338
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 66954 32614 67574 58000
rect 66954 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 67574 32614
rect 66954 32294 67574 32378
rect 66954 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 67574 32294
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 32058
rect 73794 39454 74414 58000
rect 73794 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 74414 39454
rect 73794 39134 74414 39218
rect 73794 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 74414 39134
rect 73794 3454 74414 38898
rect 73794 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 74414 3454
rect 73794 3134 74414 3218
rect 73794 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 74414 3134
rect 73794 -346 74414 2898
rect 73794 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 74414 -346
rect 73794 -666 74414 -582
rect 73794 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 74414 -666
rect 73794 -1894 74414 -902
rect 77514 43174 78134 58000
rect 77514 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 78134 43174
rect 77514 42854 78134 42938
rect 77514 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 78134 42854
rect 77514 7174 78134 42618
rect 77514 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 78134 7174
rect 77514 6854 78134 6938
rect 77514 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 78134 6854
rect 77514 -2266 78134 6618
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 46894 81854 58000
rect 81234 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 81854 46894
rect 81234 46574 81854 46658
rect 81234 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 81854 46574
rect 81234 10894 81854 46338
rect 81234 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 81854 10894
rect 81234 10574 81854 10658
rect 81234 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 81854 10574
rect 81234 -4186 81854 10338
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 84954 50614 85574 58000
rect 84954 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 85574 50614
rect 84954 50294 85574 50378
rect 84954 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 85574 50294
rect 84954 14614 85574 50058
rect 84954 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 85574 14614
rect 84954 14294 85574 14378
rect 84954 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 85574 14294
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 14058
rect 91794 57454 92414 58000
rect 91794 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 92414 57454
rect 91794 57134 92414 57218
rect 91794 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 92414 57134
rect 91794 21454 92414 56898
rect 91794 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 92414 21454
rect 91794 21134 92414 21218
rect 91794 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 92414 21134
rect 91794 -1306 92414 20898
rect 91794 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 92414 -1306
rect 91794 -1626 92414 -1542
rect 91794 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 92414 -1626
rect 91794 -1894 92414 -1862
rect 95514 25174 96134 58000
rect 95514 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 96134 25174
rect 95514 24854 96134 24938
rect 95514 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 96134 24854
rect 95514 -3226 96134 24618
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 28894 99854 58000
rect 99234 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 99854 28894
rect 99234 28574 99854 28658
rect 99234 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 99854 28574
rect 99234 -5146 99854 28338
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 102954 32614 103574 58000
rect 102954 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 103574 32614
rect 102954 32294 103574 32378
rect 102954 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 103574 32294
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 32058
rect 109794 39454 110414 58000
rect 109794 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 110414 39454
rect 109794 39134 110414 39218
rect 109794 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 110414 39134
rect 109794 3454 110414 38898
rect 109794 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 110414 3454
rect 109794 3134 110414 3218
rect 109794 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 110414 3134
rect 109794 -346 110414 2898
rect 109794 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 110414 -346
rect 109794 -666 110414 -582
rect 109794 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 110414 -666
rect 109794 -1894 110414 -902
rect 113514 43174 114134 58000
rect 113514 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 114134 43174
rect 113514 42854 114134 42938
rect 113514 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 114134 42854
rect 113514 7174 114134 42618
rect 113514 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 114134 7174
rect 113514 6854 114134 6938
rect 113514 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 114134 6854
rect 113514 -2266 114134 6618
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 46894 117854 58000
rect 117234 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 117854 46894
rect 117234 46574 117854 46658
rect 117234 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 117854 46574
rect 117234 10894 117854 46338
rect 117234 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 117854 10894
rect 117234 10574 117854 10658
rect 117234 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 117854 10574
rect 117234 -4186 117854 10338
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 120954 50614 121574 58000
rect 120954 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 121574 50614
rect 120954 50294 121574 50378
rect 120954 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 121574 50294
rect 120954 14614 121574 50058
rect 120954 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 121574 14614
rect 120954 14294 121574 14378
rect 120954 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 121574 14294
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 14058
rect 127794 57454 128414 58000
rect 127794 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 128414 57454
rect 127794 57134 128414 57218
rect 127794 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 128414 57134
rect 127794 21454 128414 56898
rect 127794 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 128414 21454
rect 127794 21134 128414 21218
rect 127794 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 128414 21134
rect 127794 -1306 128414 20898
rect 127794 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 128414 -1306
rect 127794 -1626 128414 -1542
rect 127794 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 128414 -1626
rect 127794 -1894 128414 -1862
rect 131514 25174 132134 58000
rect 131514 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 132134 25174
rect 131514 24854 132134 24938
rect 131514 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 132134 24854
rect 131514 -3226 132134 24618
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 28894 135854 58000
rect 135234 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 135854 28894
rect 135234 28574 135854 28658
rect 135234 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 135854 28574
rect 135234 -5146 135854 28338
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 138954 32614 139574 58000
rect 138954 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 139574 32614
rect 138954 32294 139574 32378
rect 138954 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 139574 32294
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 32058
rect 145794 39454 146414 58000
rect 145794 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 146414 39454
rect 145794 39134 146414 39218
rect 145794 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 146414 39134
rect 145794 3454 146414 38898
rect 145794 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 146414 3454
rect 145794 3134 146414 3218
rect 145794 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 146414 3134
rect 145794 -346 146414 2898
rect 145794 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 146414 -346
rect 145794 -666 146414 -582
rect 145794 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 146414 -666
rect 145794 -1894 146414 -902
rect 149514 43174 150134 58000
rect 149514 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 150134 43174
rect 149514 42854 150134 42938
rect 149514 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 150134 42854
rect 149514 7174 150134 42618
rect 149514 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 150134 7174
rect 149514 6854 150134 6938
rect 149514 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 150134 6854
rect 149514 -2266 150134 6618
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 46894 153854 58000
rect 153234 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 153854 46894
rect 153234 46574 153854 46658
rect 153234 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 153854 46574
rect 153234 10894 153854 46338
rect 153234 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 153854 10894
rect 153234 10574 153854 10658
rect 153234 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 153854 10574
rect 153234 -4186 153854 10338
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 156954 50614 157574 58000
rect 156954 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 157574 50614
rect 156954 50294 157574 50378
rect 156954 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 157574 50294
rect 156954 14614 157574 50058
rect 156954 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 157574 14614
rect 156954 14294 157574 14378
rect 156954 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 157574 14294
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 14058
rect 163794 57454 164414 58000
rect 163794 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 164414 57454
rect 163794 57134 164414 57218
rect 163794 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 164414 57134
rect 163794 21454 164414 56898
rect 163794 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 164414 21454
rect 163794 21134 164414 21218
rect 163794 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 164414 21134
rect 163794 -1306 164414 20898
rect 163794 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 164414 -1306
rect 163794 -1626 164414 -1542
rect 163794 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 164414 -1626
rect 163794 -1894 164414 -1862
rect 167514 25174 168134 58000
rect 167514 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 168134 25174
rect 167514 24854 168134 24938
rect 167514 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 168134 24854
rect 167514 -3226 168134 24618
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 28894 171854 58000
rect 171234 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 171854 28894
rect 171234 28574 171854 28658
rect 171234 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 171854 28574
rect 171234 -5146 171854 28338
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 174954 32614 175574 58000
rect 174954 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 175574 32614
rect 174954 32294 175574 32378
rect 174954 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 175574 32294
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 32058
rect 181794 39454 182414 58000
rect 181794 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 182414 39454
rect 181794 39134 182414 39218
rect 181794 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 182414 39134
rect 181794 3454 182414 38898
rect 181794 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 182414 3454
rect 181794 3134 182414 3218
rect 181794 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 182414 3134
rect 181794 -346 182414 2898
rect 181794 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 182414 -346
rect 181794 -666 182414 -582
rect 181794 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 182414 -666
rect 181794 -1894 182414 -902
rect 185514 43174 186134 58000
rect 185514 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 186134 43174
rect 185514 42854 186134 42938
rect 185514 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 186134 42854
rect 185514 7174 186134 42618
rect 185514 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 186134 7174
rect 185514 6854 186134 6938
rect 185514 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 186134 6854
rect 185514 -2266 186134 6618
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 46894 189854 58000
rect 189234 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 189854 46894
rect 189234 46574 189854 46658
rect 189234 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 189854 46574
rect 189234 10894 189854 46338
rect 189234 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 189854 10894
rect 189234 10574 189854 10658
rect 189234 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 189854 10574
rect 189234 -4186 189854 10338
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 192954 50614 193574 58000
rect 192954 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 193574 50614
rect 192954 50294 193574 50378
rect 192954 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 193574 50294
rect 192954 14614 193574 50058
rect 192954 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 193574 14614
rect 192954 14294 193574 14378
rect 192954 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 193574 14294
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 14058
rect 199794 57454 200414 58000
rect 199794 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 200414 57454
rect 199794 57134 200414 57218
rect 199794 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 200414 57134
rect 199794 21454 200414 56898
rect 199794 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 200414 21454
rect 199794 21134 200414 21218
rect 199794 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 200414 21134
rect 199794 -1306 200414 20898
rect 199794 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 200414 -1306
rect 199794 -1626 200414 -1542
rect 199794 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 200414 -1626
rect 199794 -1894 200414 -1862
rect 203514 25174 204134 58000
rect 203514 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 204134 25174
rect 203514 24854 204134 24938
rect 203514 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 204134 24854
rect 203514 -3226 204134 24618
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 28894 207854 58000
rect 207234 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 207854 28894
rect 207234 28574 207854 28658
rect 207234 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 207854 28574
rect 207234 -5146 207854 28338
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 210954 32614 211574 58000
rect 210954 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 211574 32614
rect 210954 32294 211574 32378
rect 210954 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 211574 32294
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 32058
rect 217794 39454 218414 58000
rect 217794 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 218414 39454
rect 217794 39134 218414 39218
rect 217794 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 218414 39134
rect 217794 3454 218414 38898
rect 217794 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 218414 3454
rect 217794 3134 218414 3218
rect 217794 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 218414 3134
rect 217794 -346 218414 2898
rect 217794 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 218414 -346
rect 217794 -666 218414 -582
rect 217794 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 218414 -666
rect 217794 -1894 218414 -902
rect 221514 43174 222134 58000
rect 224910 57901 224970 60691
rect 225094 60213 225154 232190
rect 225234 228924 225854 262338
rect 226195 234292 226261 234293
rect 226195 234228 226196 234292
rect 226260 234228 226261 234292
rect 226195 234227 226261 234228
rect 226011 234156 226077 234157
rect 226011 234092 226012 234156
rect 226076 234092 226077 234156
rect 226011 234091 226077 234092
rect 225275 228580 225341 228581
rect 225275 228516 225276 228580
rect 225340 228516 225341 228580
rect 225275 228515 225341 228516
rect 225091 60212 225157 60213
rect 225091 60148 225092 60212
rect 225156 60148 225157 60212
rect 225091 60147 225157 60148
rect 225278 58170 225338 228515
rect 226014 147797 226074 234091
rect 226011 147796 226077 147797
rect 226011 147732 226012 147796
rect 226076 147732 226077 147796
rect 226011 147731 226077 147732
rect 226198 143445 226258 234227
rect 226195 143444 226261 143445
rect 226195 143380 226196 143444
rect 226260 143380 226261 143444
rect 226195 143379 226261 143380
rect 225459 70276 225525 70277
rect 225459 70212 225460 70276
rect 225524 70212 225525 70276
rect 225459 70211 225525 70212
rect 225462 60757 225522 70211
rect 225459 60756 225525 60757
rect 225459 60692 225460 60756
rect 225524 60692 225525 60756
rect 225459 60691 225525 60692
rect 226382 58445 226442 398243
rect 235950 398173 236010 399470
rect 227851 398172 227917 398173
rect 227851 398108 227852 398172
rect 227916 398108 227917 398172
rect 227851 398107 227917 398108
rect 235947 398172 236013 398173
rect 235947 398108 235948 398172
rect 236012 398108 236013 398172
rect 235947 398107 236013 398108
rect 227667 397900 227733 397901
rect 227667 397836 227668 397900
rect 227732 397836 227733 397900
rect 227667 397835 227733 397836
rect 226747 236876 226813 236877
rect 226747 236812 226748 236876
rect 226812 236812 226813 236876
rect 226747 236811 226813 236812
rect 226563 235380 226629 235381
rect 226563 235316 226564 235380
rect 226628 235316 226629 235380
rect 226563 235315 226629 235316
rect 226566 75037 226626 235315
rect 226750 113389 226810 236811
rect 226931 225724 226997 225725
rect 226931 225660 226932 225724
rect 226996 225660 226997 225724
rect 226931 225659 226997 225660
rect 226934 126989 226994 225659
rect 226931 126988 226997 126989
rect 226931 126924 226932 126988
rect 226996 126924 226997 126988
rect 226931 126923 226997 126924
rect 226747 113388 226813 113389
rect 226747 113324 226748 113388
rect 226812 113324 226813 113388
rect 226747 113323 226813 113324
rect 226563 75036 226629 75037
rect 226563 74972 226564 75036
rect 226628 74972 226629 75036
rect 226563 74971 226629 74972
rect 227670 59261 227730 397835
rect 227667 59260 227733 59261
rect 227667 59196 227668 59260
rect 227732 59196 227733 59260
rect 227667 59195 227733 59196
rect 227854 58853 227914 398107
rect 228954 374614 229574 398000
rect 228954 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 229574 374614
rect 228954 374294 229574 374378
rect 228954 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 229574 374294
rect 228954 338614 229574 374058
rect 228954 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 229574 338614
rect 228954 338294 229574 338378
rect 228954 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 229574 338294
rect 228954 302614 229574 338058
rect 228954 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 229574 302614
rect 228954 302294 229574 302378
rect 228954 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 229574 302294
rect 228954 266614 229574 302058
rect 228954 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 229574 266614
rect 228954 266294 229574 266378
rect 228954 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 229574 266294
rect 228219 233476 228285 233477
rect 228219 233412 228220 233476
rect 228284 233412 228285 233476
rect 228219 233411 228285 233412
rect 228222 111893 228282 233411
rect 228954 230614 229574 266058
rect 228954 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 229574 230614
rect 228954 230294 229574 230378
rect 228954 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 229574 230294
rect 228954 194614 229574 230058
rect 228954 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 229574 194614
rect 228954 194294 229574 194378
rect 228954 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 229574 194294
rect 228954 158614 229574 194058
rect 228954 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 229574 158614
rect 228954 158294 229574 158378
rect 228954 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 229574 158294
rect 228954 122614 229574 158058
rect 228954 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 229574 122614
rect 228954 122294 229574 122378
rect 228954 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 229574 122294
rect 228219 111892 228285 111893
rect 228219 111828 228220 111892
rect 228284 111828 228285 111892
rect 228219 111827 228285 111828
rect 228954 86614 229574 122058
rect 228954 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 229574 86614
rect 228954 86294 229574 86378
rect 228954 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 229574 86294
rect 227851 58852 227917 58853
rect 227851 58788 227852 58852
rect 227916 58788 227917 58852
rect 227851 58787 227917 58788
rect 226379 58444 226445 58445
rect 226379 58380 226380 58444
rect 226444 58380 226445 58444
rect 226379 58379 226445 58380
rect 225094 58110 225338 58170
rect 224907 57900 224973 57901
rect 224907 57836 224908 57900
rect 224972 57836 224973 57900
rect 224907 57835 224973 57836
rect 225094 57490 225154 58110
rect 224910 57430 225154 57490
rect 224910 57085 224970 57430
rect 224907 57084 224973 57085
rect 224907 57020 224908 57084
rect 224972 57020 224973 57084
rect 224907 57019 224973 57020
rect 221514 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 222134 43174
rect 221514 42854 222134 42938
rect 221514 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 222134 42854
rect 221514 7174 222134 42618
rect 221514 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 222134 7174
rect 221514 6854 222134 6938
rect 221514 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 222134 6854
rect 221514 -2266 222134 6618
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 46894 225854 58000
rect 225234 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 225854 46894
rect 225234 46574 225854 46658
rect 225234 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 225854 46574
rect 225234 10894 225854 46338
rect 225234 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 225854 10894
rect 225234 10574 225854 10658
rect 225234 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 225854 10574
rect 225234 -4186 225854 10338
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 228954 50614 229574 86058
rect 228954 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 229574 50614
rect 228954 50294 229574 50378
rect 228954 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 229574 50294
rect 228954 14614 229574 50058
rect 228954 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 229574 14614
rect 228954 14294 229574 14378
rect 228954 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 229574 14294
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 14058
rect 235794 381454 236414 398000
rect 237054 397357 237114 399470
rect 237051 397356 237117 397357
rect 237051 397292 237052 397356
rect 237116 397292 237117 397356
rect 237051 397291 237117 397292
rect 238158 396813 238218 399470
rect 239262 397357 239322 399470
rect 239259 397356 239325 397357
rect 239259 397292 239260 397356
rect 239324 397292 239325 397356
rect 239259 397291 239325 397292
rect 238155 396812 238221 396813
rect 238155 396748 238156 396812
rect 238220 396748 238221 396812
rect 238155 396747 238221 396748
rect 235794 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 236414 381454
rect 235794 381134 236414 381218
rect 235794 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 236414 381134
rect 235794 345454 236414 380898
rect 235794 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 236414 345454
rect 235794 345134 236414 345218
rect 235794 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 236414 345134
rect 235794 309454 236414 344898
rect 235794 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 236414 309454
rect 235794 309134 236414 309218
rect 235794 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 236414 309134
rect 235794 273454 236414 308898
rect 235794 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 236414 273454
rect 235794 273134 236414 273218
rect 235794 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 236414 273134
rect 235794 237454 236414 272898
rect 235794 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 236414 237454
rect 235794 237134 236414 237218
rect 235794 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 236414 237134
rect 235794 201454 236414 236898
rect 235794 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 236414 201454
rect 235794 201134 236414 201218
rect 235794 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 236414 201134
rect 235794 165454 236414 200898
rect 235794 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 236414 165454
rect 235794 165134 236414 165218
rect 235794 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 236414 165134
rect 235794 129454 236414 164898
rect 235794 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 236414 129454
rect 235794 129134 236414 129218
rect 235794 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 236414 129134
rect 235794 93454 236414 128898
rect 235794 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 236414 93454
rect 235794 93134 236414 93218
rect 235794 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 236414 93134
rect 235794 57454 236414 92898
rect 235794 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 236414 57454
rect 235794 57134 236414 57218
rect 235794 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 236414 57134
rect 235794 21454 236414 56898
rect 235794 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 236414 21454
rect 235794 21134 236414 21218
rect 235794 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 236414 21134
rect 235794 -1306 236414 20898
rect 235794 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 236414 -1306
rect 235794 -1626 236414 -1542
rect 235794 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 236414 -1626
rect 235794 -1894 236414 -1862
rect 239514 385174 240134 398000
rect 240550 396813 240610 399470
rect 241654 399470 241828 399530
rect 242942 399470 243188 399530
rect 244216 399530 244276 400106
rect 245440 399530 245500 400106
rect 246528 399530 246588 400106
rect 244216 399470 244290 399530
rect 241654 397357 241714 399470
rect 242942 397357 243002 399470
rect 241651 397356 241717 397357
rect 241651 397292 241652 397356
rect 241716 397292 241717 397356
rect 241651 397291 241717 397292
rect 242939 397356 243005 397357
rect 242939 397292 242940 397356
rect 243004 397292 243005 397356
rect 242939 397291 243005 397292
rect 240547 396812 240613 396813
rect 240547 396748 240548 396812
rect 240612 396748 240613 396812
rect 240547 396747 240613 396748
rect 239514 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 240134 385174
rect 239514 384854 240134 384938
rect 239514 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 240134 384854
rect 239514 349174 240134 384618
rect 239514 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 240134 349174
rect 239514 348854 240134 348938
rect 239514 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 240134 348854
rect 239514 313174 240134 348618
rect 239514 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 240134 313174
rect 239514 312854 240134 312938
rect 239514 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 240134 312854
rect 239514 277174 240134 312618
rect 239514 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 240134 277174
rect 239514 276854 240134 276938
rect 239514 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 240134 276854
rect 239514 241174 240134 276618
rect 239514 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 240134 241174
rect 239514 240854 240134 240938
rect 239514 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 240134 240854
rect 239514 205174 240134 240618
rect 239514 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 240134 205174
rect 239514 204854 240134 204938
rect 239514 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 240134 204854
rect 239514 169174 240134 204618
rect 239514 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 240134 169174
rect 239514 168854 240134 168938
rect 239514 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 240134 168854
rect 239514 133174 240134 168618
rect 239514 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 240134 133174
rect 239514 132854 240134 132938
rect 239514 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 240134 132854
rect 239514 97174 240134 132618
rect 239514 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 240134 97174
rect 239514 96854 240134 96938
rect 239514 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 240134 96854
rect 239514 61174 240134 96618
rect 239514 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 240134 61174
rect 239514 60854 240134 60938
rect 239514 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 240134 60854
rect 239514 25174 240134 60618
rect 239514 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 240134 25174
rect 239514 24854 240134 24938
rect 239514 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 240134 24854
rect 239514 -3226 240134 24618
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 388894 243854 398000
rect 244230 396813 244290 399470
rect 245334 399470 245500 399530
rect 246438 399470 246588 399530
rect 247616 399530 247676 400106
rect 248296 399530 248356 400106
rect 248704 399530 248764 400106
rect 247616 399470 247786 399530
rect 245334 397357 245394 399470
rect 245331 397356 245397 397357
rect 245331 397292 245332 397356
rect 245396 397292 245397 397356
rect 245331 397291 245397 397292
rect 246438 396813 246498 399470
rect 244227 396812 244293 396813
rect 244227 396748 244228 396812
rect 244292 396748 244293 396812
rect 244227 396747 244293 396748
rect 246435 396812 246501 396813
rect 246435 396748 246436 396812
rect 246500 396748 246501 396812
rect 246435 396747 246501 396748
rect 243234 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 243854 388894
rect 243234 388574 243854 388658
rect 243234 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 243854 388574
rect 243234 352894 243854 388338
rect 243234 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 243854 352894
rect 243234 352574 243854 352658
rect 243234 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 243854 352574
rect 243234 316894 243854 352338
rect 243234 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 243854 316894
rect 243234 316574 243854 316658
rect 243234 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 243854 316574
rect 243234 280894 243854 316338
rect 243234 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 243854 280894
rect 243234 280574 243854 280658
rect 243234 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 243854 280574
rect 243234 244894 243854 280338
rect 243234 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 243854 244894
rect 243234 244574 243854 244658
rect 243234 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 243854 244574
rect 243234 208894 243854 244338
rect 243234 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 243854 208894
rect 243234 208574 243854 208658
rect 243234 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 243854 208574
rect 243234 172894 243854 208338
rect 243234 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 243854 172894
rect 243234 172574 243854 172658
rect 243234 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 243854 172574
rect 243234 136894 243854 172338
rect 243234 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 243854 136894
rect 243234 136574 243854 136658
rect 243234 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 243854 136574
rect 243234 100894 243854 136338
rect 243234 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 243854 100894
rect 243234 100574 243854 100658
rect 243234 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 243854 100574
rect 243234 64894 243854 100338
rect 243234 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 243854 64894
rect 243234 64574 243854 64658
rect 243234 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 243854 64574
rect 243234 28894 243854 64338
rect 243234 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 243854 28894
rect 243234 28574 243854 28658
rect 243234 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 243854 28574
rect 243234 -5146 243854 28338
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 246954 392614 247574 398000
rect 247726 396677 247786 399470
rect 248278 399470 248356 399530
rect 248646 399470 248764 399530
rect 250064 399530 250124 400106
rect 250744 399530 250804 400106
rect 251288 399530 251348 400106
rect 252376 399530 252436 400106
rect 253464 399530 253524 400106
rect 250064 399470 250178 399530
rect 248278 396813 248338 399470
rect 248646 397357 248706 399470
rect 248643 397356 248709 397357
rect 248643 397292 248644 397356
rect 248708 397292 248709 397356
rect 248643 397291 248709 397292
rect 250118 396813 250178 399470
rect 250670 399470 250804 399530
rect 251222 399470 251348 399530
rect 252326 399470 252436 399530
rect 253430 399470 253524 399530
rect 253600 399530 253660 400106
rect 254552 399530 254612 400106
rect 255912 399530 255972 400106
rect 253600 399470 253674 399530
rect 250670 397357 250730 399470
rect 250667 397356 250733 397357
rect 250667 397292 250668 397356
rect 250732 397292 250733 397356
rect 250667 397291 250733 397292
rect 251222 396813 251282 399470
rect 248275 396812 248341 396813
rect 248275 396748 248276 396812
rect 248340 396748 248341 396812
rect 248275 396747 248341 396748
rect 250115 396812 250181 396813
rect 250115 396748 250116 396812
rect 250180 396748 250181 396812
rect 250115 396747 250181 396748
rect 251219 396812 251285 396813
rect 251219 396748 251220 396812
rect 251284 396748 251285 396812
rect 251219 396747 251285 396748
rect 252326 396677 252386 399470
rect 253430 397357 253490 399470
rect 253614 397357 253674 399470
rect 254534 399470 254612 399530
rect 255822 399470 255972 399530
rect 256048 399530 256108 400106
rect 257000 399530 257060 400106
rect 256048 399470 256250 399530
rect 253427 397356 253493 397357
rect 253427 397292 253428 397356
rect 253492 397292 253493 397356
rect 253427 397291 253493 397292
rect 253611 397356 253677 397357
rect 253611 397292 253612 397356
rect 253676 397292 253677 397356
rect 253611 397291 253677 397292
rect 247723 396676 247789 396677
rect 247723 396612 247724 396676
rect 247788 396612 247789 396676
rect 247723 396611 247789 396612
rect 252323 396676 252389 396677
rect 252323 396612 252324 396676
rect 252388 396612 252389 396676
rect 252323 396611 252389 396612
rect 246954 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 247574 392614
rect 246954 392294 247574 392378
rect 246954 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 247574 392294
rect 246954 356614 247574 392058
rect 246954 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 247574 356614
rect 246954 356294 247574 356378
rect 246954 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 247574 356294
rect 246954 320614 247574 356058
rect 246954 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 247574 320614
rect 246954 320294 247574 320378
rect 246954 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 247574 320294
rect 246954 284614 247574 320058
rect 246954 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 247574 284614
rect 246954 284294 247574 284378
rect 246954 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 247574 284294
rect 246954 248614 247574 284058
rect 246954 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 247574 248614
rect 246954 248294 247574 248378
rect 246954 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 247574 248294
rect 246954 212614 247574 248058
rect 246954 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 247574 212614
rect 246954 212294 247574 212378
rect 246954 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 247574 212294
rect 246954 176614 247574 212058
rect 246954 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 247574 176614
rect 246954 176294 247574 176378
rect 246954 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 247574 176294
rect 246954 140614 247574 176058
rect 246954 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 247574 140614
rect 246954 140294 247574 140378
rect 246954 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 247574 140294
rect 246954 104614 247574 140058
rect 246954 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 247574 104614
rect 246954 104294 247574 104378
rect 246954 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 247574 104294
rect 246954 68614 247574 104058
rect 246954 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 247574 68614
rect 246954 68294 247574 68378
rect 246954 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 247574 68294
rect 246954 32614 247574 68058
rect 246954 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 247574 32614
rect 246954 32294 247574 32378
rect 246954 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 247574 32294
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 32058
rect 253794 363454 254414 398000
rect 254534 396813 254594 399470
rect 255822 396813 255882 399470
rect 256190 397357 256250 399470
rect 256926 399470 257060 399530
rect 258088 399530 258148 400106
rect 258496 399530 258556 400106
rect 258088 399470 258274 399530
rect 256187 397356 256253 397357
rect 256187 397292 256188 397356
rect 256252 397292 256253 397356
rect 256187 397291 256253 397292
rect 256926 396813 256986 399470
rect 254531 396812 254597 396813
rect 254531 396748 254532 396812
rect 254596 396748 254597 396812
rect 254531 396747 254597 396748
rect 255819 396812 255885 396813
rect 255819 396748 255820 396812
rect 255884 396748 255885 396812
rect 255819 396747 255885 396748
rect 256923 396812 256989 396813
rect 256923 396748 256924 396812
rect 256988 396748 256989 396812
rect 256923 396747 256989 396748
rect 253794 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 254414 363454
rect 253794 363134 254414 363218
rect 253794 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 254414 363134
rect 253794 327454 254414 362898
rect 253794 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 254414 327454
rect 253794 327134 254414 327218
rect 253794 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 254414 327134
rect 253794 291454 254414 326898
rect 253794 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 254414 291454
rect 253794 291134 254414 291218
rect 253794 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 254414 291134
rect 253794 255454 254414 290898
rect 253794 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 254414 255454
rect 253794 255134 254414 255218
rect 253794 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 254414 255134
rect 253794 219454 254414 254898
rect 253794 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 254414 219454
rect 253794 219134 254414 219218
rect 253794 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 254414 219134
rect 253794 183454 254414 218898
rect 253794 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 254414 183454
rect 253794 183134 254414 183218
rect 253794 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 254414 183134
rect 253794 147454 254414 182898
rect 253794 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 254414 147454
rect 253794 147134 254414 147218
rect 253794 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 254414 147134
rect 253794 111454 254414 146898
rect 253794 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 254414 111454
rect 253794 111134 254414 111218
rect 253794 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 254414 111134
rect 253794 75454 254414 110898
rect 253794 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 254414 75454
rect 253794 75134 254414 75218
rect 253794 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 254414 75134
rect 253794 39454 254414 74898
rect 253794 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 254414 39454
rect 253794 39134 254414 39218
rect 253794 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 254414 39134
rect 253794 3454 254414 38898
rect 253794 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 254414 3454
rect 253794 3134 254414 3218
rect 253794 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 254414 3134
rect 253794 -346 254414 2898
rect 253794 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 254414 -346
rect 253794 -666 254414 -582
rect 253794 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 254414 -666
rect 253794 -1894 254414 -902
rect 257514 367174 258134 398000
rect 258214 396810 258274 399470
rect 258398 399470 258556 399530
rect 259448 399530 259508 400106
rect 260672 399530 260732 400106
rect 261080 399530 261140 400106
rect 259448 399470 259562 399530
rect 258398 396949 258458 399470
rect 258395 396948 258461 396949
rect 258395 396884 258396 396948
rect 258460 396884 258461 396948
rect 258395 396883 258461 396884
rect 259502 396813 259562 399470
rect 260606 399470 260732 399530
rect 260974 399470 261140 399530
rect 261760 399530 261820 400106
rect 262848 399530 262908 400106
rect 261760 399470 262138 399530
rect 258395 396812 258461 396813
rect 258395 396810 258396 396812
rect 258214 396750 258396 396810
rect 258395 396748 258396 396750
rect 258460 396748 258461 396812
rect 258395 396747 258461 396748
rect 259499 396812 259565 396813
rect 259499 396748 259500 396812
rect 259564 396748 259565 396812
rect 259499 396747 259565 396748
rect 260606 396677 260666 399470
rect 260974 397357 261034 399470
rect 260971 397356 261037 397357
rect 260971 397292 260972 397356
rect 261036 397292 261037 397356
rect 260971 397291 261037 397292
rect 260603 396676 260669 396677
rect 260603 396612 260604 396676
rect 260668 396612 260669 396676
rect 260603 396611 260669 396612
rect 257514 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 258134 367174
rect 257514 366854 258134 366938
rect 257514 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 258134 366854
rect 257514 331174 258134 366618
rect 257514 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 258134 331174
rect 257514 330854 258134 330938
rect 257514 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 258134 330854
rect 257514 295174 258134 330618
rect 257514 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 258134 295174
rect 257514 294854 258134 294938
rect 257514 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 258134 294854
rect 257514 259174 258134 294618
rect 257514 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 258134 259174
rect 257514 258854 258134 258938
rect 257514 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 258134 258854
rect 257514 223174 258134 258618
rect 257514 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 258134 223174
rect 257514 222854 258134 222938
rect 257514 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 258134 222854
rect 257514 187174 258134 222618
rect 257514 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 258134 187174
rect 257514 186854 258134 186938
rect 257514 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 258134 186854
rect 257514 151174 258134 186618
rect 257514 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 258134 151174
rect 257514 150854 258134 150938
rect 257514 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 258134 150854
rect 257514 115174 258134 150618
rect 257514 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 258134 115174
rect 257514 114854 258134 114938
rect 257514 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 258134 114854
rect 257514 79174 258134 114618
rect 257514 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 258134 79174
rect 257514 78854 258134 78938
rect 257514 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 258134 78854
rect 257514 43174 258134 78618
rect 257514 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 258134 43174
rect 257514 42854 258134 42938
rect 257514 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 258134 42854
rect 257514 7174 258134 42618
rect 257514 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 258134 7174
rect 257514 6854 258134 6938
rect 257514 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 258134 6854
rect 257514 -2266 258134 6618
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 370894 261854 398000
rect 262078 397357 262138 399470
rect 262814 399470 262908 399530
rect 263528 399530 263588 400106
rect 263936 399530 263996 400106
rect 265296 399530 265356 400106
rect 265976 399530 266036 400106
rect 266384 399530 266444 400106
rect 267608 399530 267668 400106
rect 263528 399470 263610 399530
rect 262075 397356 262141 397357
rect 262075 397292 262076 397356
rect 262140 397292 262141 397356
rect 262075 397291 262141 397292
rect 262814 396813 262874 399470
rect 263550 397357 263610 399470
rect 263918 399470 263996 399530
rect 265206 399470 265356 399530
rect 265942 399470 266036 399530
rect 266310 399470 266444 399530
rect 267598 399470 267668 399530
rect 268288 399530 268348 400106
rect 268696 399530 268756 400106
rect 269784 399530 269844 400106
rect 271008 399530 271068 400106
rect 268288 399470 268394 399530
rect 268696 399470 268762 399530
rect 269784 399470 269866 399530
rect 263547 397356 263613 397357
rect 263547 397292 263548 397356
rect 263612 397292 263613 397356
rect 263547 397291 263613 397292
rect 263918 397221 263978 399470
rect 265206 398173 265266 399470
rect 265203 398172 265269 398173
rect 265203 398108 265204 398172
rect 265268 398108 265269 398172
rect 265203 398107 265269 398108
rect 263915 397220 263981 397221
rect 263915 397156 263916 397220
rect 263980 397156 263981 397220
rect 263915 397155 263981 397156
rect 262811 396812 262877 396813
rect 262811 396748 262812 396812
rect 262876 396748 262877 396812
rect 262811 396747 262877 396748
rect 261234 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 261854 370894
rect 261234 370574 261854 370658
rect 261234 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 261854 370574
rect 261234 334894 261854 370338
rect 261234 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 261854 334894
rect 261234 334574 261854 334658
rect 261234 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 261854 334574
rect 261234 298894 261854 334338
rect 261234 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 261854 298894
rect 261234 298574 261854 298658
rect 261234 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 261854 298574
rect 261234 262894 261854 298338
rect 261234 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 261854 262894
rect 261234 262574 261854 262658
rect 261234 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 261854 262574
rect 261234 226894 261854 262338
rect 261234 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 261854 226894
rect 261234 226574 261854 226658
rect 261234 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 261854 226574
rect 261234 190894 261854 226338
rect 261234 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 261854 190894
rect 261234 190574 261854 190658
rect 261234 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 261854 190574
rect 261234 154894 261854 190338
rect 261234 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 261854 154894
rect 261234 154574 261854 154658
rect 261234 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 261854 154574
rect 261234 118894 261854 154338
rect 261234 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 261854 118894
rect 261234 118574 261854 118658
rect 261234 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 261854 118574
rect 261234 82894 261854 118338
rect 261234 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 261854 82894
rect 261234 82574 261854 82658
rect 261234 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 261854 82574
rect 261234 46894 261854 82338
rect 261234 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 261854 46894
rect 261234 46574 261854 46658
rect 261234 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 261854 46574
rect 261234 10894 261854 46338
rect 261234 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 261854 10894
rect 261234 10574 261854 10658
rect 261234 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 261854 10574
rect 261234 -4186 261854 10338
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 264954 374614 265574 398000
rect 265942 396813 266002 399470
rect 266310 396813 266370 399470
rect 265939 396812 266005 396813
rect 265939 396748 265940 396812
rect 266004 396748 266005 396812
rect 265939 396747 266005 396748
rect 266307 396812 266373 396813
rect 266307 396748 266308 396812
rect 266372 396748 266373 396812
rect 266307 396747 266373 396748
rect 267598 396677 267658 399470
rect 268334 396813 268394 399470
rect 268331 396812 268397 396813
rect 268331 396748 268332 396812
rect 268396 396748 268397 396812
rect 268331 396747 268397 396748
rect 268702 396677 268762 399470
rect 269806 396813 269866 399470
rect 270910 399470 271068 399530
rect 271144 399530 271204 400106
rect 272232 399530 272292 400106
rect 273320 399530 273380 400106
rect 273592 399530 273652 400106
rect 274408 399530 274468 400106
rect 275768 399530 275828 400106
rect 271144 399470 271338 399530
rect 272232 399470 272626 399530
rect 270910 396813 270970 399470
rect 271278 397357 271338 399470
rect 271275 397356 271341 397357
rect 271275 397292 271276 397356
rect 271340 397292 271341 397356
rect 271275 397291 271341 397292
rect 269803 396812 269869 396813
rect 269803 396748 269804 396812
rect 269868 396748 269869 396812
rect 269803 396747 269869 396748
rect 270907 396812 270973 396813
rect 270907 396748 270908 396812
rect 270972 396748 270973 396812
rect 270907 396747 270973 396748
rect 267595 396676 267661 396677
rect 267595 396612 267596 396676
rect 267660 396612 267661 396676
rect 267595 396611 267661 396612
rect 268699 396676 268765 396677
rect 268699 396612 268700 396676
rect 268764 396612 268765 396676
rect 268699 396611 268765 396612
rect 264954 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 265574 374614
rect 264954 374294 265574 374378
rect 264954 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 265574 374294
rect 264954 338614 265574 374058
rect 264954 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 265574 338614
rect 264954 338294 265574 338378
rect 264954 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 265574 338294
rect 264954 302614 265574 338058
rect 264954 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 265574 302614
rect 264954 302294 265574 302378
rect 264954 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 265574 302294
rect 264954 266614 265574 302058
rect 264954 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 265574 266614
rect 264954 266294 265574 266378
rect 264954 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 265574 266294
rect 264954 230614 265574 266058
rect 264954 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 265574 230614
rect 264954 230294 265574 230378
rect 264954 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 265574 230294
rect 264954 194614 265574 230058
rect 264954 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 265574 194614
rect 264954 194294 265574 194378
rect 264954 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 265574 194294
rect 264954 158614 265574 194058
rect 264954 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 265574 158614
rect 264954 158294 265574 158378
rect 264954 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 265574 158294
rect 264954 122614 265574 158058
rect 264954 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 265574 122614
rect 264954 122294 265574 122378
rect 264954 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 265574 122294
rect 264954 86614 265574 122058
rect 264954 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 265574 86614
rect 264954 86294 265574 86378
rect 264954 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 265574 86294
rect 264954 50614 265574 86058
rect 264954 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 265574 50614
rect 264954 50294 265574 50378
rect 264954 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 265574 50294
rect 264954 14614 265574 50058
rect 264954 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 265574 14614
rect 264954 14294 265574 14378
rect 264954 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 265574 14294
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 14058
rect 271794 381454 272414 398000
rect 272566 396813 272626 399470
rect 273302 399470 273380 399530
rect 273486 399470 273652 399530
rect 274406 399470 274468 399530
rect 275326 399470 275828 399530
rect 276040 399530 276100 400106
rect 276992 399530 277052 400106
rect 276040 399470 276306 399530
rect 273302 397357 273362 399470
rect 273299 397356 273365 397357
rect 273299 397292 273300 397356
rect 273364 397292 273365 397356
rect 273299 397291 273365 397292
rect 273486 397221 273546 399470
rect 274406 397357 274466 399470
rect 275326 397357 275386 399470
rect 274403 397356 274469 397357
rect 274403 397292 274404 397356
rect 274468 397292 274469 397356
rect 274403 397291 274469 397292
rect 275323 397356 275389 397357
rect 275323 397292 275324 397356
rect 275388 397292 275389 397356
rect 275323 397291 275389 397292
rect 273483 397220 273549 397221
rect 273483 397156 273484 397220
rect 273548 397156 273549 397220
rect 273483 397155 273549 397156
rect 272563 396812 272629 396813
rect 272563 396748 272564 396812
rect 272628 396748 272629 396812
rect 272563 396747 272629 396748
rect 271794 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 272414 381454
rect 271794 381134 272414 381218
rect 271794 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 272414 381134
rect 271794 345454 272414 380898
rect 271794 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 272414 345454
rect 271794 345134 272414 345218
rect 271794 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 272414 345134
rect 271794 309454 272414 344898
rect 271794 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 272414 309454
rect 271794 309134 272414 309218
rect 271794 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 272414 309134
rect 271794 273454 272414 308898
rect 271794 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 272414 273454
rect 271794 273134 272414 273218
rect 271794 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 272414 273134
rect 271794 237454 272414 272898
rect 271794 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 272414 237454
rect 271794 237134 272414 237218
rect 271794 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 272414 237134
rect 271794 201454 272414 236898
rect 271794 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 272414 201454
rect 271794 201134 272414 201218
rect 271794 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 272414 201134
rect 271794 165454 272414 200898
rect 271794 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 272414 165454
rect 271794 165134 272414 165218
rect 271794 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 272414 165134
rect 271794 129454 272414 164898
rect 271794 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 272414 129454
rect 271794 129134 272414 129218
rect 271794 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 272414 129134
rect 271794 93454 272414 128898
rect 271794 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 272414 93454
rect 271794 93134 272414 93218
rect 271794 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 272414 93134
rect 271794 57454 272414 92898
rect 271794 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 272414 57454
rect 271794 57134 272414 57218
rect 271794 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 272414 57134
rect 271794 21454 272414 56898
rect 271794 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 272414 21454
rect 271794 21134 272414 21218
rect 271794 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 272414 21134
rect 271794 -1306 272414 20898
rect 271794 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 272414 -1306
rect 271794 -1626 272414 -1542
rect 271794 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 272414 -1626
rect 271794 -1894 272414 -1862
rect 275514 385174 276134 398000
rect 276246 396813 276306 399470
rect 276982 399470 277052 399530
rect 278080 399530 278140 400106
rect 278488 399530 278548 400106
rect 279168 399530 279228 400106
rect 280936 399530 280996 400106
rect 278080 399470 278146 399530
rect 276982 397357 277042 399470
rect 278086 397357 278146 399470
rect 278454 399470 278548 399530
rect 279006 399470 279228 399530
rect 280846 399470 280996 399530
rect 283520 399530 283580 400106
rect 285968 399530 286028 400106
rect 288280 399530 288340 400106
rect 291000 399530 291060 400106
rect 293448 399530 293508 400106
rect 283520 399470 283850 399530
rect 285968 399470 286058 399530
rect 276979 397356 277045 397357
rect 276979 397292 276980 397356
rect 277044 397292 277045 397356
rect 276979 397291 277045 397292
rect 278083 397356 278149 397357
rect 278083 397292 278084 397356
rect 278148 397292 278149 397356
rect 278083 397291 278149 397292
rect 278454 396813 278514 399470
rect 279006 396813 279066 399470
rect 276243 396812 276309 396813
rect 276243 396748 276244 396812
rect 276308 396748 276309 396812
rect 276243 396747 276309 396748
rect 278451 396812 278517 396813
rect 278451 396748 278452 396812
rect 278516 396748 278517 396812
rect 278451 396747 278517 396748
rect 279003 396812 279069 396813
rect 279003 396748 279004 396812
rect 279068 396748 279069 396812
rect 279003 396747 279069 396748
rect 275514 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 276134 385174
rect 275514 384854 276134 384938
rect 275514 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 276134 384854
rect 275514 349174 276134 384618
rect 275514 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 276134 349174
rect 275514 348854 276134 348938
rect 275514 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 276134 348854
rect 275514 313174 276134 348618
rect 275514 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 276134 313174
rect 275514 312854 276134 312938
rect 275514 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 276134 312854
rect 275514 277174 276134 312618
rect 275514 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 276134 277174
rect 275514 276854 276134 276938
rect 275514 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 276134 276854
rect 275514 241174 276134 276618
rect 275514 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 276134 241174
rect 275514 240854 276134 240938
rect 275514 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 276134 240854
rect 275514 205174 276134 240618
rect 275514 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 276134 205174
rect 275514 204854 276134 204938
rect 275514 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 276134 204854
rect 275514 169174 276134 204618
rect 275514 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 276134 169174
rect 275514 168854 276134 168938
rect 275514 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 276134 168854
rect 275514 133174 276134 168618
rect 275514 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 276134 133174
rect 275514 132854 276134 132938
rect 275514 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 276134 132854
rect 275514 97174 276134 132618
rect 275514 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 276134 97174
rect 275514 96854 276134 96938
rect 275514 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 276134 96854
rect 275514 61174 276134 96618
rect 275514 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 276134 61174
rect 275514 60854 276134 60938
rect 275514 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 276134 60854
rect 275514 25174 276134 60618
rect 275514 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 276134 25174
rect 275514 24854 276134 24938
rect 275514 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 276134 24854
rect 275514 -3226 276134 24618
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 388894 279854 398000
rect 280846 396813 280906 399470
rect 280843 396812 280909 396813
rect 280843 396748 280844 396812
rect 280908 396748 280909 396812
rect 280843 396747 280909 396748
rect 279234 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 279854 388894
rect 279234 388574 279854 388658
rect 279234 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 279854 388574
rect 279234 352894 279854 388338
rect 279234 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 279854 352894
rect 279234 352574 279854 352658
rect 279234 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 279854 352574
rect 279234 316894 279854 352338
rect 279234 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 279854 316894
rect 279234 316574 279854 316658
rect 279234 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 279854 316574
rect 279234 280894 279854 316338
rect 279234 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 279854 280894
rect 279234 280574 279854 280658
rect 279234 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 279854 280574
rect 279234 244894 279854 280338
rect 279234 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 279854 244894
rect 279234 244574 279854 244658
rect 279234 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 279854 244574
rect 279234 208894 279854 244338
rect 279234 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 279854 208894
rect 279234 208574 279854 208658
rect 279234 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 279854 208574
rect 279234 172894 279854 208338
rect 279234 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 279854 172894
rect 279234 172574 279854 172658
rect 279234 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 279854 172574
rect 279234 136894 279854 172338
rect 279234 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 279854 136894
rect 279234 136574 279854 136658
rect 279234 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 279854 136574
rect 279234 100894 279854 136338
rect 279234 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 279854 100894
rect 279234 100574 279854 100658
rect 279234 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 279854 100574
rect 279234 64894 279854 100338
rect 279234 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 279854 64894
rect 279234 64574 279854 64658
rect 279234 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 279854 64574
rect 279234 28894 279854 64338
rect 279234 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 279854 28894
rect 279234 28574 279854 28658
rect 279234 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 279854 28574
rect 279234 -5146 279854 28338
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 282954 392614 283574 398000
rect 283790 396813 283850 399470
rect 285998 396813 286058 399470
rect 288206 399470 288340 399530
rect 290966 399470 291060 399530
rect 293358 399470 293508 399530
rect 295896 399530 295956 400106
rect 298480 399530 298540 400106
rect 300928 399530 300988 400106
rect 303512 399530 303572 400106
rect 305960 399530 306020 400106
rect 295896 399470 295994 399530
rect 298480 399470 298570 399530
rect 288206 396813 288266 399470
rect 283787 396812 283853 396813
rect 283787 396748 283788 396812
rect 283852 396748 283853 396812
rect 283787 396747 283853 396748
rect 285995 396812 286061 396813
rect 285995 396748 285996 396812
rect 286060 396748 286061 396812
rect 285995 396747 286061 396748
rect 288203 396812 288269 396813
rect 288203 396748 288204 396812
rect 288268 396748 288269 396812
rect 288203 396747 288269 396748
rect 282954 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 283574 392614
rect 282954 392294 283574 392378
rect 282954 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 283574 392294
rect 282954 356614 283574 392058
rect 282954 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 283574 356614
rect 282954 356294 283574 356378
rect 282954 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 283574 356294
rect 282954 320614 283574 356058
rect 282954 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 283574 320614
rect 282954 320294 283574 320378
rect 282954 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 283574 320294
rect 282954 284614 283574 320058
rect 282954 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 283574 284614
rect 282954 284294 283574 284378
rect 282954 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 283574 284294
rect 282954 248614 283574 284058
rect 282954 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 283574 248614
rect 282954 248294 283574 248378
rect 282954 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 283574 248294
rect 282954 212614 283574 248058
rect 282954 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 283574 212614
rect 282954 212294 283574 212378
rect 282954 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 283574 212294
rect 282954 176614 283574 212058
rect 282954 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 283574 176614
rect 282954 176294 283574 176378
rect 282954 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 283574 176294
rect 282954 140614 283574 176058
rect 282954 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 283574 140614
rect 282954 140294 283574 140378
rect 282954 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 283574 140294
rect 282954 104614 283574 140058
rect 282954 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 283574 104614
rect 282954 104294 283574 104378
rect 282954 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 283574 104294
rect 282954 68614 283574 104058
rect 282954 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 283574 68614
rect 282954 68294 283574 68378
rect 282954 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 283574 68294
rect 282954 32614 283574 68058
rect 282954 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 283574 32614
rect 282954 32294 283574 32378
rect 282954 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 283574 32294
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 32058
rect 289794 363454 290414 398000
rect 290966 397357 291026 399470
rect 293358 397357 293418 399470
rect 290963 397356 291029 397357
rect 290963 397292 290964 397356
rect 291028 397292 291029 397356
rect 290963 397291 291029 397292
rect 293355 397356 293421 397357
rect 293355 397292 293356 397356
rect 293420 397292 293421 397356
rect 293355 397291 293421 397292
rect 289794 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 290414 363454
rect 289794 363134 290414 363218
rect 289794 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 290414 363134
rect 289794 327454 290414 362898
rect 289794 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 290414 327454
rect 289794 327134 290414 327218
rect 289794 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 290414 327134
rect 289794 291454 290414 326898
rect 289794 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 290414 291454
rect 289794 291134 290414 291218
rect 289794 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 290414 291134
rect 289794 255454 290414 290898
rect 289794 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 290414 255454
rect 289794 255134 290414 255218
rect 289794 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 290414 255134
rect 289794 219454 290414 254898
rect 289794 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 290414 219454
rect 289794 219134 290414 219218
rect 289794 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 290414 219134
rect 289794 183454 290414 218898
rect 289794 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 290414 183454
rect 289794 183134 290414 183218
rect 289794 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 290414 183134
rect 289794 147454 290414 182898
rect 289794 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 290414 147454
rect 289794 147134 290414 147218
rect 289794 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 290414 147134
rect 289794 111454 290414 146898
rect 289794 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 290414 111454
rect 289794 111134 290414 111218
rect 289794 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 290414 111134
rect 289794 75454 290414 110898
rect 289794 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 290414 75454
rect 289794 75134 290414 75218
rect 289794 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 290414 75134
rect 289794 39454 290414 74898
rect 289794 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 290414 39454
rect 289794 39134 290414 39218
rect 289794 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 290414 39134
rect 289794 3454 290414 38898
rect 289794 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 290414 3454
rect 289794 3134 290414 3218
rect 289794 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 290414 3134
rect 289794 -346 290414 2898
rect 289794 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 290414 -346
rect 289794 -666 290414 -582
rect 289794 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 290414 -666
rect 289794 -1894 290414 -902
rect 293514 367174 294134 398000
rect 295934 396813 295994 399470
rect 295931 396812 295997 396813
rect 295931 396748 295932 396812
rect 295996 396748 295997 396812
rect 295931 396747 295997 396748
rect 293514 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 294134 367174
rect 293514 366854 294134 366938
rect 293514 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 294134 366854
rect 293514 331174 294134 366618
rect 293514 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 294134 331174
rect 293514 330854 294134 330938
rect 293514 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 294134 330854
rect 293514 295174 294134 330618
rect 293514 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 294134 295174
rect 293514 294854 294134 294938
rect 293514 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 294134 294854
rect 293514 259174 294134 294618
rect 293514 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 294134 259174
rect 293514 258854 294134 258938
rect 293514 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 294134 258854
rect 293514 223174 294134 258618
rect 293514 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 294134 223174
rect 293514 222854 294134 222938
rect 293514 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 294134 222854
rect 293514 187174 294134 222618
rect 293514 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 294134 187174
rect 293514 186854 294134 186938
rect 293514 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 294134 186854
rect 293514 151174 294134 186618
rect 293514 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 294134 151174
rect 293514 150854 294134 150938
rect 293514 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 294134 150854
rect 293514 115174 294134 150618
rect 293514 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 294134 115174
rect 293514 114854 294134 114938
rect 293514 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 294134 114854
rect 293514 79174 294134 114618
rect 293514 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 294134 79174
rect 293514 78854 294134 78938
rect 293514 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 294134 78854
rect 293514 43174 294134 78618
rect 293514 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 294134 43174
rect 293514 42854 294134 42938
rect 293514 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 294134 42854
rect 293514 7174 294134 42618
rect 293514 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 294134 7174
rect 293514 6854 294134 6938
rect 293514 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 294134 6854
rect 293514 -2266 294134 6618
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 370894 297854 398000
rect 298510 397357 298570 399470
rect 300902 399470 300988 399530
rect 303478 399470 303572 399530
rect 305870 399470 306020 399530
rect 308544 399530 308604 400106
rect 310992 399530 311052 400106
rect 313440 399530 313500 400106
rect 315888 399530 315948 400106
rect 318472 399530 318532 400106
rect 308544 399470 308690 399530
rect 310992 399470 311082 399530
rect 300902 398173 300962 399470
rect 300899 398172 300965 398173
rect 300899 398108 300900 398172
rect 300964 398108 300965 398172
rect 300899 398107 300965 398108
rect 298507 397356 298573 397357
rect 298507 397292 298508 397356
rect 298572 397292 298573 397356
rect 298507 397291 298573 397292
rect 297234 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 297854 370894
rect 297234 370574 297854 370658
rect 297234 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 297854 370574
rect 297234 334894 297854 370338
rect 297234 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 297854 334894
rect 297234 334574 297854 334658
rect 297234 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 297854 334574
rect 297234 298894 297854 334338
rect 297234 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 297854 298894
rect 297234 298574 297854 298658
rect 297234 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 297854 298574
rect 297234 262894 297854 298338
rect 297234 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 297854 262894
rect 297234 262574 297854 262658
rect 297234 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 297854 262574
rect 297234 226894 297854 262338
rect 297234 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 297854 226894
rect 297234 226574 297854 226658
rect 297234 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 297854 226574
rect 297234 190894 297854 226338
rect 297234 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 297854 190894
rect 297234 190574 297854 190658
rect 297234 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 297854 190574
rect 297234 154894 297854 190338
rect 297234 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 297854 154894
rect 297234 154574 297854 154658
rect 297234 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 297854 154574
rect 297234 118894 297854 154338
rect 297234 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 297854 118894
rect 297234 118574 297854 118658
rect 297234 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 297854 118574
rect 297234 82894 297854 118338
rect 297234 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 297854 82894
rect 297234 82574 297854 82658
rect 297234 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 297854 82574
rect 297234 46894 297854 82338
rect 297234 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 297854 46894
rect 297234 46574 297854 46658
rect 297234 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 297854 46574
rect 297234 10894 297854 46338
rect 297234 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 297854 10894
rect 297234 10574 297854 10658
rect 297234 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 297854 10574
rect 297234 -4186 297854 10338
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 300954 374614 301574 398000
rect 303478 396813 303538 399470
rect 305870 396813 305930 399470
rect 303475 396812 303541 396813
rect 303475 396748 303476 396812
rect 303540 396748 303541 396812
rect 303475 396747 303541 396748
rect 305867 396812 305933 396813
rect 305867 396748 305868 396812
rect 305932 396748 305933 396812
rect 305867 396747 305933 396748
rect 300954 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 301574 374614
rect 300954 374294 301574 374378
rect 300954 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 301574 374294
rect 300954 338614 301574 374058
rect 300954 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 301574 338614
rect 300954 338294 301574 338378
rect 300954 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 301574 338294
rect 300954 302614 301574 338058
rect 300954 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 301574 302614
rect 300954 302294 301574 302378
rect 300954 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 301574 302294
rect 300954 266614 301574 302058
rect 300954 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 301574 266614
rect 300954 266294 301574 266378
rect 300954 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 301574 266294
rect 300954 230614 301574 266058
rect 300954 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 301574 230614
rect 300954 230294 301574 230378
rect 300954 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 301574 230294
rect 300954 194614 301574 230058
rect 300954 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 301574 194614
rect 300954 194294 301574 194378
rect 300954 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 301574 194294
rect 300954 158614 301574 194058
rect 300954 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 301574 158614
rect 300954 158294 301574 158378
rect 300954 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 301574 158294
rect 300954 122614 301574 158058
rect 300954 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 301574 122614
rect 300954 122294 301574 122378
rect 300954 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 301574 122294
rect 300954 86614 301574 122058
rect 300954 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 301574 86614
rect 300954 86294 301574 86378
rect 300954 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 301574 86294
rect 300954 50614 301574 86058
rect 300954 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 301574 50614
rect 300954 50294 301574 50378
rect 300954 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 301574 50294
rect 300954 14614 301574 50058
rect 300954 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 301574 14614
rect 300954 14294 301574 14378
rect 300954 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 301574 14294
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 14058
rect 307794 381454 308414 398000
rect 308630 397357 308690 399470
rect 311022 397357 311082 399470
rect 313414 399470 313500 399530
rect 315806 399470 315948 399530
rect 318382 399470 318532 399530
rect 320920 399530 320980 400106
rect 323368 399530 323428 400106
rect 325952 399530 326012 400106
rect 343224 399530 343284 400106
rect 320920 399470 321018 399530
rect 308627 397356 308693 397357
rect 308627 397292 308628 397356
rect 308692 397292 308693 397356
rect 308627 397291 308693 397292
rect 311019 397356 311085 397357
rect 311019 397292 311020 397356
rect 311084 397292 311085 397356
rect 311019 397291 311085 397292
rect 307794 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 308414 381454
rect 307794 381134 308414 381218
rect 307794 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 308414 381134
rect 307794 345454 308414 380898
rect 307794 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 308414 345454
rect 307794 345134 308414 345218
rect 307794 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 308414 345134
rect 307794 309454 308414 344898
rect 307794 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 308414 309454
rect 307794 309134 308414 309218
rect 307794 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 308414 309134
rect 307794 273454 308414 308898
rect 307794 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 308414 273454
rect 307794 273134 308414 273218
rect 307794 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 308414 273134
rect 307794 237454 308414 272898
rect 307794 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 308414 237454
rect 307794 237134 308414 237218
rect 307794 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 308414 237134
rect 307794 201454 308414 236898
rect 307794 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 308414 201454
rect 307794 201134 308414 201218
rect 307794 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 308414 201134
rect 307794 165454 308414 200898
rect 307794 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 308414 165454
rect 307794 165134 308414 165218
rect 307794 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 308414 165134
rect 307794 129454 308414 164898
rect 307794 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 308414 129454
rect 307794 129134 308414 129218
rect 307794 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 308414 129134
rect 307794 93454 308414 128898
rect 307794 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 308414 93454
rect 307794 93134 308414 93218
rect 307794 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 308414 93134
rect 307794 57454 308414 92898
rect 307794 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 308414 57454
rect 307794 57134 308414 57218
rect 307794 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 308414 57134
rect 307794 21454 308414 56898
rect 307794 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 308414 21454
rect 307794 21134 308414 21218
rect 307794 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 308414 21134
rect 307794 -1306 308414 20898
rect 307794 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 308414 -1306
rect 307794 -1626 308414 -1542
rect 307794 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 308414 -1626
rect 307794 -1894 308414 -1862
rect 311514 385174 312134 398000
rect 313414 397357 313474 399470
rect 315806 398173 315866 399470
rect 315803 398172 315869 398173
rect 315803 398108 315804 398172
rect 315868 398108 315869 398172
rect 315803 398107 315869 398108
rect 313411 397356 313477 397357
rect 313411 397292 313412 397356
rect 313476 397292 313477 397356
rect 313411 397291 313477 397292
rect 311514 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 312134 385174
rect 311514 384854 312134 384938
rect 311514 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 312134 384854
rect 311514 349174 312134 384618
rect 311514 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 312134 349174
rect 311514 348854 312134 348938
rect 311514 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 312134 348854
rect 311514 313174 312134 348618
rect 311514 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 312134 313174
rect 311514 312854 312134 312938
rect 311514 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 312134 312854
rect 311514 277174 312134 312618
rect 311514 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 312134 277174
rect 311514 276854 312134 276938
rect 311514 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 312134 276854
rect 311514 241174 312134 276618
rect 311514 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 312134 241174
rect 311514 240854 312134 240938
rect 311514 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 312134 240854
rect 311514 205174 312134 240618
rect 311514 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 312134 205174
rect 311514 204854 312134 204938
rect 311514 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 312134 204854
rect 311514 169174 312134 204618
rect 311514 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 312134 169174
rect 311514 168854 312134 168938
rect 311514 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 312134 168854
rect 311514 133174 312134 168618
rect 311514 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 312134 133174
rect 311514 132854 312134 132938
rect 311514 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 312134 132854
rect 311514 97174 312134 132618
rect 311514 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 312134 97174
rect 311514 96854 312134 96938
rect 311514 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 312134 96854
rect 311514 61174 312134 96618
rect 311514 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 312134 61174
rect 311514 60854 312134 60938
rect 311514 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 312134 60854
rect 311514 25174 312134 60618
rect 311514 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 312134 25174
rect 311514 24854 312134 24938
rect 311514 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 312134 24854
rect 311514 -3226 312134 24618
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 388894 315854 398000
rect 318382 396813 318442 399470
rect 318379 396812 318445 396813
rect 318379 396748 318380 396812
rect 318444 396748 318445 396812
rect 318379 396747 318445 396748
rect 315234 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 315854 388894
rect 315234 388574 315854 388658
rect 315234 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 315854 388574
rect 315234 352894 315854 388338
rect 315234 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 315854 352894
rect 315234 352574 315854 352658
rect 315234 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 315854 352574
rect 315234 316894 315854 352338
rect 315234 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 315854 316894
rect 315234 316574 315854 316658
rect 315234 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 315854 316574
rect 315234 280894 315854 316338
rect 315234 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 315854 280894
rect 315234 280574 315854 280658
rect 315234 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 315854 280574
rect 315234 244894 315854 280338
rect 315234 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 315854 244894
rect 315234 244574 315854 244658
rect 315234 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 315854 244574
rect 315234 208894 315854 244338
rect 315234 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 315854 208894
rect 315234 208574 315854 208658
rect 315234 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 315854 208574
rect 315234 172894 315854 208338
rect 315234 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 315854 172894
rect 315234 172574 315854 172658
rect 315234 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 315854 172574
rect 315234 136894 315854 172338
rect 315234 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 315854 136894
rect 315234 136574 315854 136658
rect 315234 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 315854 136574
rect 315234 100894 315854 136338
rect 315234 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 315854 100894
rect 315234 100574 315854 100658
rect 315234 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 315854 100574
rect 315234 64894 315854 100338
rect 315234 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 315854 64894
rect 315234 64574 315854 64658
rect 315234 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 315854 64574
rect 315234 28894 315854 64338
rect 315234 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 315854 28894
rect 315234 28574 315854 28658
rect 315234 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 315854 28574
rect 315234 -5146 315854 28338
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 318954 392614 319574 398000
rect 320958 396813 321018 399470
rect 323350 399470 323428 399530
rect 325926 399470 326012 399530
rect 343222 399470 343284 399530
rect 343360 399530 343420 400106
rect 343360 399470 343466 399530
rect 323350 396813 323410 399470
rect 325926 398173 325986 399470
rect 325923 398172 325989 398173
rect 325923 398108 325924 398172
rect 325988 398108 325989 398172
rect 325923 398107 325989 398108
rect 320955 396812 321021 396813
rect 320955 396748 320956 396812
rect 321020 396748 321021 396812
rect 320955 396747 321021 396748
rect 323347 396812 323413 396813
rect 323347 396748 323348 396812
rect 323412 396748 323413 396812
rect 323347 396747 323413 396748
rect 318954 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 319574 392614
rect 318954 392294 319574 392378
rect 318954 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 319574 392294
rect 318954 356614 319574 392058
rect 318954 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 319574 356614
rect 318954 356294 319574 356378
rect 318954 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 319574 356294
rect 318954 320614 319574 356058
rect 318954 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 319574 320614
rect 318954 320294 319574 320378
rect 318954 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 319574 320294
rect 318954 284614 319574 320058
rect 318954 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 319574 284614
rect 318954 284294 319574 284378
rect 318954 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 319574 284294
rect 318954 248614 319574 284058
rect 318954 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 319574 248614
rect 318954 248294 319574 248378
rect 318954 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 319574 248294
rect 318954 212614 319574 248058
rect 318954 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 319574 212614
rect 318954 212294 319574 212378
rect 318954 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 319574 212294
rect 318954 176614 319574 212058
rect 318954 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 319574 176614
rect 318954 176294 319574 176378
rect 318954 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 319574 176294
rect 318954 140614 319574 176058
rect 318954 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 319574 140614
rect 318954 140294 319574 140378
rect 318954 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 319574 140294
rect 318954 104614 319574 140058
rect 318954 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 319574 104614
rect 318954 104294 319574 104378
rect 318954 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 319574 104294
rect 318954 68614 319574 104058
rect 318954 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 319574 68614
rect 318954 68294 319574 68378
rect 318954 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 319574 68294
rect 318954 32614 319574 68058
rect 318954 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 319574 32614
rect 318954 32294 319574 32378
rect 318954 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 319574 32294
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 32058
rect 325794 363454 326414 398000
rect 325794 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 326414 363454
rect 325794 363134 326414 363218
rect 325794 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 326414 363134
rect 325794 327454 326414 362898
rect 325794 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 326414 327454
rect 325794 327134 326414 327218
rect 325794 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 326414 327134
rect 325794 291454 326414 326898
rect 325794 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 326414 291454
rect 325794 291134 326414 291218
rect 325794 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 326414 291134
rect 325794 255454 326414 290898
rect 325794 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 326414 255454
rect 325794 255134 326414 255218
rect 325794 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 326414 255134
rect 325794 219454 326414 254898
rect 325794 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 326414 219454
rect 325794 219134 326414 219218
rect 325794 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 326414 219134
rect 325794 183454 326414 218898
rect 325794 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 326414 183454
rect 325794 183134 326414 183218
rect 325794 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 326414 183134
rect 325794 147454 326414 182898
rect 325794 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 326414 147454
rect 325794 147134 326414 147218
rect 325794 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 326414 147134
rect 325794 111454 326414 146898
rect 325794 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 326414 111454
rect 325794 111134 326414 111218
rect 325794 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 326414 111134
rect 325794 75454 326414 110898
rect 325794 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 326414 75454
rect 325794 75134 326414 75218
rect 325794 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 326414 75134
rect 325794 39454 326414 74898
rect 325794 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 326414 39454
rect 325794 39134 326414 39218
rect 325794 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 326414 39134
rect 325794 3454 326414 38898
rect 325794 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 326414 3454
rect 325794 3134 326414 3218
rect 325794 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 326414 3134
rect 325794 -346 326414 2898
rect 325794 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 326414 -346
rect 325794 -666 326414 -582
rect 325794 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 326414 -666
rect 325794 -1894 326414 -902
rect 329514 367174 330134 398000
rect 329514 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 330134 367174
rect 329514 366854 330134 366938
rect 329514 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 330134 366854
rect 329514 331174 330134 366618
rect 329514 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 330134 331174
rect 329514 330854 330134 330938
rect 329514 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 330134 330854
rect 329514 295174 330134 330618
rect 329514 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 330134 295174
rect 329514 294854 330134 294938
rect 329514 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 330134 294854
rect 329514 259174 330134 294618
rect 329514 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 330134 259174
rect 329514 258854 330134 258938
rect 329514 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 330134 258854
rect 329514 223174 330134 258618
rect 329514 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 330134 223174
rect 329514 222854 330134 222938
rect 329514 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 330134 222854
rect 329514 187174 330134 222618
rect 329514 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 330134 187174
rect 329514 186854 330134 186938
rect 329514 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 330134 186854
rect 329514 151174 330134 186618
rect 329514 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 330134 151174
rect 329514 150854 330134 150938
rect 329514 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 330134 150854
rect 329514 115174 330134 150618
rect 329514 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 330134 115174
rect 329514 114854 330134 114938
rect 329514 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 330134 114854
rect 329514 79174 330134 114618
rect 329514 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 330134 79174
rect 329514 78854 330134 78938
rect 329514 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 330134 78854
rect 329514 43174 330134 78618
rect 329514 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 330134 43174
rect 329514 42854 330134 42938
rect 329514 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 330134 42854
rect 329514 7174 330134 42618
rect 329514 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 330134 7174
rect 329514 6854 330134 6938
rect 329514 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 330134 6854
rect 329514 -2266 330134 6618
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 370894 333854 398000
rect 333234 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 333854 370894
rect 333234 370574 333854 370658
rect 333234 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 333854 370574
rect 333234 334894 333854 370338
rect 333234 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 333854 334894
rect 333234 334574 333854 334658
rect 333234 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 333854 334574
rect 333234 298894 333854 334338
rect 333234 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 333854 298894
rect 333234 298574 333854 298658
rect 333234 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 333854 298574
rect 333234 262894 333854 298338
rect 333234 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 333854 262894
rect 333234 262574 333854 262658
rect 333234 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 333854 262574
rect 333234 226894 333854 262338
rect 333234 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 333854 226894
rect 333234 226574 333854 226658
rect 333234 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 333854 226574
rect 333234 190894 333854 226338
rect 333234 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 333854 190894
rect 333234 190574 333854 190658
rect 333234 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 333854 190574
rect 333234 154894 333854 190338
rect 333234 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 333854 154894
rect 333234 154574 333854 154658
rect 333234 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 333854 154574
rect 333234 118894 333854 154338
rect 333234 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 333854 118894
rect 333234 118574 333854 118658
rect 333234 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 333854 118574
rect 333234 82894 333854 118338
rect 333234 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 333854 82894
rect 333234 82574 333854 82658
rect 333234 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 333854 82574
rect 333234 46894 333854 82338
rect 333234 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 333854 46894
rect 333234 46574 333854 46658
rect 333234 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 333854 46574
rect 333234 10894 333854 46338
rect 333234 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 333854 10894
rect 333234 10574 333854 10658
rect 333234 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 333854 10574
rect 333234 -4186 333854 10338
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 336954 374614 337574 398000
rect 343222 397357 343282 399470
rect 343219 397356 343285 397357
rect 343219 397292 343220 397356
rect 343284 397292 343285 397356
rect 343219 397291 343285 397292
rect 343406 396813 343466 399470
rect 361794 399454 362414 434898
rect 361794 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 362414 399454
rect 361794 399134 362414 399218
rect 361794 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 362414 399134
rect 343403 396812 343469 396813
rect 343403 396748 343404 396812
rect 343468 396748 343469 396812
rect 343403 396747 343469 396748
rect 336954 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 337574 374614
rect 336954 374294 337574 374378
rect 336954 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 337574 374294
rect 336954 338614 337574 374058
rect 336954 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 337574 338614
rect 336954 338294 337574 338378
rect 336954 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 337574 338294
rect 336954 302614 337574 338058
rect 336954 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 337574 302614
rect 336954 302294 337574 302378
rect 336954 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 337574 302294
rect 336954 266614 337574 302058
rect 336954 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 337574 266614
rect 336954 266294 337574 266378
rect 336954 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 337574 266294
rect 336954 230614 337574 266058
rect 336954 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 337574 230614
rect 336954 230294 337574 230378
rect 336954 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 337574 230294
rect 336954 194614 337574 230058
rect 336954 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 337574 194614
rect 336954 194294 337574 194378
rect 336954 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 337574 194294
rect 336954 158614 337574 194058
rect 336954 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 337574 158614
rect 336954 158294 337574 158378
rect 336954 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 337574 158294
rect 336954 122614 337574 158058
rect 336954 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 337574 122614
rect 336954 122294 337574 122378
rect 336954 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 337574 122294
rect 336954 86614 337574 122058
rect 336954 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 337574 86614
rect 336954 86294 337574 86378
rect 336954 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 337574 86294
rect 336954 50614 337574 86058
rect 336954 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 337574 50614
rect 336954 50294 337574 50378
rect 336954 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 337574 50294
rect 336954 14614 337574 50058
rect 336954 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 337574 14614
rect 336954 14294 337574 14378
rect 336954 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 337574 14294
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 14058
rect 343794 381454 344414 398000
rect 343794 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 344414 381454
rect 343794 381134 344414 381218
rect 343794 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 344414 381134
rect 343794 345454 344414 380898
rect 343794 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 344414 345454
rect 343794 345134 344414 345218
rect 343794 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 344414 345134
rect 343794 309454 344414 344898
rect 343794 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 344414 309454
rect 343794 309134 344414 309218
rect 343794 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 344414 309134
rect 343794 273454 344414 308898
rect 343794 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 344414 273454
rect 343794 273134 344414 273218
rect 343794 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 344414 273134
rect 343794 237454 344414 272898
rect 343794 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 344414 237454
rect 343794 237134 344414 237218
rect 343794 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 344414 237134
rect 343794 201454 344414 236898
rect 343794 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 344414 201454
rect 343794 201134 344414 201218
rect 343794 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 344414 201134
rect 343794 165454 344414 200898
rect 343794 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 344414 165454
rect 343794 165134 344414 165218
rect 343794 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 344414 165134
rect 343794 129454 344414 164898
rect 343794 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 344414 129454
rect 343794 129134 344414 129218
rect 343794 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 344414 129134
rect 343794 93454 344414 128898
rect 343794 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 344414 93454
rect 343794 93134 344414 93218
rect 343794 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 344414 93134
rect 343794 57454 344414 92898
rect 343794 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 344414 57454
rect 343794 57134 344414 57218
rect 343794 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 344414 57134
rect 343794 21454 344414 56898
rect 343794 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 344414 21454
rect 343794 21134 344414 21218
rect 343794 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 344414 21134
rect 343794 -1306 344414 20898
rect 343794 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 344414 -1306
rect 343794 -1626 344414 -1542
rect 343794 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 344414 -1626
rect 343794 -1894 344414 -1862
rect 347514 385174 348134 398000
rect 347514 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 348134 385174
rect 347514 384854 348134 384938
rect 347514 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 348134 384854
rect 347514 349174 348134 384618
rect 347514 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 348134 349174
rect 347514 348854 348134 348938
rect 347514 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 348134 348854
rect 347514 313174 348134 348618
rect 347514 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 348134 313174
rect 347514 312854 348134 312938
rect 347514 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 348134 312854
rect 347514 277174 348134 312618
rect 347514 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 348134 277174
rect 347514 276854 348134 276938
rect 347514 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 348134 276854
rect 347514 241174 348134 276618
rect 347514 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 348134 241174
rect 347514 240854 348134 240938
rect 347514 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 348134 240854
rect 347514 205174 348134 240618
rect 347514 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 348134 205174
rect 347514 204854 348134 204938
rect 347514 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 348134 204854
rect 347514 169174 348134 204618
rect 347514 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 348134 169174
rect 347514 168854 348134 168938
rect 347514 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 348134 168854
rect 347514 133174 348134 168618
rect 347514 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 348134 133174
rect 347514 132854 348134 132938
rect 347514 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 348134 132854
rect 347514 97174 348134 132618
rect 347514 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 348134 97174
rect 347514 96854 348134 96938
rect 347514 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 348134 96854
rect 347514 61174 348134 96618
rect 347514 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 348134 61174
rect 347514 60854 348134 60938
rect 347514 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 348134 60854
rect 347514 25174 348134 60618
rect 347514 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 348134 25174
rect 347514 24854 348134 24938
rect 347514 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 348134 24854
rect 347514 -3226 348134 24618
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 388894 351854 398000
rect 351234 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 351854 388894
rect 351234 388574 351854 388658
rect 351234 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 351854 388574
rect 351234 352894 351854 388338
rect 351234 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 351854 352894
rect 351234 352574 351854 352658
rect 351234 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 351854 352574
rect 351234 316894 351854 352338
rect 351234 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 351854 316894
rect 351234 316574 351854 316658
rect 351234 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 351854 316574
rect 351234 280894 351854 316338
rect 351234 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 351854 280894
rect 351234 280574 351854 280658
rect 351234 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 351854 280574
rect 351234 244894 351854 280338
rect 351234 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 351854 244894
rect 351234 244574 351854 244658
rect 351234 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 351854 244574
rect 351234 208894 351854 244338
rect 351234 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 351854 208894
rect 351234 208574 351854 208658
rect 351234 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 351854 208574
rect 351234 172894 351854 208338
rect 351234 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 351854 172894
rect 351234 172574 351854 172658
rect 351234 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 351854 172574
rect 351234 136894 351854 172338
rect 351234 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 351854 136894
rect 351234 136574 351854 136658
rect 351234 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 351854 136574
rect 351234 100894 351854 136338
rect 351234 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 351854 100894
rect 351234 100574 351854 100658
rect 351234 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 351854 100574
rect 351234 64894 351854 100338
rect 351234 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 351854 64894
rect 351234 64574 351854 64658
rect 351234 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 351854 64574
rect 351234 28894 351854 64338
rect 351234 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 351854 28894
rect 351234 28574 351854 28658
rect 351234 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 351854 28574
rect 351234 -5146 351854 28338
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 354954 392614 355574 398000
rect 354954 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 355574 392614
rect 354954 392294 355574 392378
rect 354954 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 355574 392294
rect 354954 356614 355574 392058
rect 354954 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 355574 356614
rect 354954 356294 355574 356378
rect 354954 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 355574 356294
rect 354954 320614 355574 356058
rect 354954 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 355574 320614
rect 354954 320294 355574 320378
rect 354954 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 355574 320294
rect 354954 284614 355574 320058
rect 354954 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 355574 284614
rect 354954 284294 355574 284378
rect 354954 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 355574 284294
rect 354954 248614 355574 284058
rect 354954 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 355574 248614
rect 354954 248294 355574 248378
rect 354954 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 355574 248294
rect 354954 212614 355574 248058
rect 354954 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 355574 212614
rect 354954 212294 355574 212378
rect 354954 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 355574 212294
rect 354954 176614 355574 212058
rect 354954 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 355574 176614
rect 354954 176294 355574 176378
rect 354954 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 355574 176294
rect 354954 140614 355574 176058
rect 354954 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 355574 140614
rect 354954 140294 355574 140378
rect 354954 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 355574 140294
rect 354954 104614 355574 140058
rect 354954 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 355574 104614
rect 354954 104294 355574 104378
rect 354954 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 355574 104294
rect 354954 68614 355574 104058
rect 354954 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 355574 68614
rect 354954 68294 355574 68378
rect 354954 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 355574 68294
rect 354954 32614 355574 68058
rect 354954 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 355574 32614
rect 354954 32294 355574 32378
rect 354954 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 355574 32294
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 32058
rect 361794 363454 362414 398898
rect 361794 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 362414 363454
rect 361794 363134 362414 363218
rect 361794 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 362414 363134
rect 361794 327454 362414 362898
rect 361794 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 362414 327454
rect 361794 327134 362414 327218
rect 361794 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 362414 327134
rect 361794 291454 362414 326898
rect 361794 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 362414 291454
rect 361794 291134 362414 291218
rect 361794 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 362414 291134
rect 361794 255454 362414 290898
rect 361794 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 362414 255454
rect 361794 255134 362414 255218
rect 361794 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 362414 255134
rect 361794 219454 362414 254898
rect 361794 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 362414 219454
rect 361794 219134 362414 219218
rect 361794 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 362414 219134
rect 361794 183454 362414 218898
rect 361794 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 362414 183454
rect 361794 183134 362414 183218
rect 361794 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 362414 183134
rect 361794 147454 362414 182898
rect 361794 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 362414 147454
rect 361794 147134 362414 147218
rect 361794 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 362414 147134
rect 361794 111454 362414 146898
rect 361794 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 362414 111454
rect 361794 111134 362414 111218
rect 361794 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 362414 111134
rect 361794 75454 362414 110898
rect 361794 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 362414 75454
rect 361794 75134 362414 75218
rect 361794 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 362414 75134
rect 361794 39454 362414 74898
rect 361794 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 362414 39454
rect 361794 39134 362414 39218
rect 361794 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 362414 39134
rect 361794 3454 362414 38898
rect 361794 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 362414 3454
rect 361794 3134 362414 3218
rect 361794 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 362414 3134
rect 361794 -346 362414 2898
rect 361794 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 362414 -346
rect 361794 -666 362414 -582
rect 361794 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 362414 -666
rect 361794 -1894 362414 -902
rect 365514 691174 366134 706202
rect 365514 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 366134 691174
rect 365514 690854 366134 690938
rect 365514 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 366134 690854
rect 365514 655174 366134 690618
rect 365514 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 366134 655174
rect 365514 654854 366134 654938
rect 365514 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 366134 654854
rect 365514 619174 366134 654618
rect 365514 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 366134 619174
rect 365514 618854 366134 618938
rect 365514 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 366134 618854
rect 365514 583174 366134 618618
rect 365514 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 366134 583174
rect 365514 582854 366134 582938
rect 365514 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 366134 582854
rect 365514 547174 366134 582618
rect 365514 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 366134 547174
rect 365514 546854 366134 546938
rect 365514 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 366134 546854
rect 365514 511174 366134 546618
rect 365514 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 366134 511174
rect 365514 510854 366134 510938
rect 365514 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 366134 510854
rect 365514 475174 366134 510618
rect 365514 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 366134 475174
rect 365514 474854 366134 474938
rect 365514 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 366134 474854
rect 365514 439174 366134 474618
rect 365514 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 366134 439174
rect 365514 438854 366134 438938
rect 365514 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 366134 438854
rect 365514 403174 366134 438618
rect 365514 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 366134 403174
rect 365514 402854 366134 402938
rect 365514 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 366134 402854
rect 365514 367174 366134 402618
rect 365514 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 366134 367174
rect 365514 366854 366134 366938
rect 365514 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 366134 366854
rect 365514 331174 366134 366618
rect 365514 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 366134 331174
rect 365514 330854 366134 330938
rect 365514 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 366134 330854
rect 365514 295174 366134 330618
rect 365514 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 366134 295174
rect 365514 294854 366134 294938
rect 365514 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 366134 294854
rect 365514 259174 366134 294618
rect 365514 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 366134 259174
rect 365514 258854 366134 258938
rect 365514 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 366134 258854
rect 365514 223174 366134 258618
rect 365514 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 366134 223174
rect 365514 222854 366134 222938
rect 365514 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 366134 222854
rect 365514 187174 366134 222618
rect 365514 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 366134 187174
rect 365514 186854 366134 186938
rect 365514 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 366134 186854
rect 365514 151174 366134 186618
rect 365514 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 366134 151174
rect 365514 150854 366134 150938
rect 365514 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 366134 150854
rect 365514 115174 366134 150618
rect 365514 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 366134 115174
rect 365514 114854 366134 114938
rect 365514 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 366134 114854
rect 365514 79174 366134 114618
rect 365514 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 366134 79174
rect 365514 78854 366134 78938
rect 365514 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 366134 78854
rect 365514 43174 366134 78618
rect 365514 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 366134 43174
rect 365514 42854 366134 42938
rect 365514 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 366134 42854
rect 365514 7174 366134 42618
rect 365514 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 366134 7174
rect 365514 6854 366134 6938
rect 365514 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 366134 6854
rect 365514 -2266 366134 6618
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 694894 369854 708122
rect 369234 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 369854 694894
rect 369234 694574 369854 694658
rect 369234 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 369854 694574
rect 369234 658894 369854 694338
rect 369234 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 369854 658894
rect 369234 658574 369854 658658
rect 369234 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 369854 658574
rect 369234 622894 369854 658338
rect 369234 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 369854 622894
rect 369234 622574 369854 622658
rect 369234 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 369854 622574
rect 369234 586894 369854 622338
rect 369234 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 369854 586894
rect 369234 586574 369854 586658
rect 369234 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 369854 586574
rect 369234 550894 369854 586338
rect 369234 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 369854 550894
rect 369234 550574 369854 550658
rect 369234 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 369854 550574
rect 369234 514894 369854 550338
rect 369234 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 369854 514894
rect 369234 514574 369854 514658
rect 369234 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 369854 514574
rect 369234 478894 369854 514338
rect 369234 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 369854 478894
rect 369234 478574 369854 478658
rect 369234 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 369854 478574
rect 369234 442894 369854 478338
rect 369234 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 369854 442894
rect 369234 442574 369854 442658
rect 369234 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 369854 442574
rect 369234 406894 369854 442338
rect 369234 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 369854 406894
rect 369234 406574 369854 406658
rect 369234 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 369854 406574
rect 369234 370894 369854 406338
rect 369234 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 369854 370894
rect 369234 370574 369854 370658
rect 369234 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 369854 370574
rect 369234 334894 369854 370338
rect 369234 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 369854 334894
rect 369234 334574 369854 334658
rect 369234 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 369854 334574
rect 369234 298894 369854 334338
rect 369234 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 369854 298894
rect 369234 298574 369854 298658
rect 369234 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 369854 298574
rect 369234 262894 369854 298338
rect 369234 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 369854 262894
rect 369234 262574 369854 262658
rect 369234 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 369854 262574
rect 369234 226894 369854 262338
rect 369234 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 369854 226894
rect 369234 226574 369854 226658
rect 369234 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 369854 226574
rect 369234 190894 369854 226338
rect 369234 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 369854 190894
rect 369234 190574 369854 190658
rect 369234 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 369854 190574
rect 369234 154894 369854 190338
rect 369234 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 369854 154894
rect 369234 154574 369854 154658
rect 369234 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 369854 154574
rect 369234 118894 369854 154338
rect 369234 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 369854 118894
rect 369234 118574 369854 118658
rect 369234 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 369854 118574
rect 369234 82894 369854 118338
rect 369234 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 369854 82894
rect 369234 82574 369854 82658
rect 369234 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 369854 82574
rect 369234 46894 369854 82338
rect 369234 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 369854 46894
rect 369234 46574 369854 46658
rect 369234 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 369854 46574
rect 369234 10894 369854 46338
rect 369234 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 369854 10894
rect 369234 10574 369854 10658
rect 369234 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 369854 10574
rect 369234 -4186 369854 10338
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 372954 698614 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 372954 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 373574 698614
rect 372954 698294 373574 698378
rect 372954 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 373574 698294
rect 372954 662614 373574 698058
rect 372954 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 373574 662614
rect 372954 662294 373574 662378
rect 372954 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 373574 662294
rect 372954 626614 373574 662058
rect 372954 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 373574 626614
rect 372954 626294 373574 626378
rect 372954 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 373574 626294
rect 372954 590614 373574 626058
rect 372954 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 373574 590614
rect 372954 590294 373574 590378
rect 372954 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 373574 590294
rect 372954 554614 373574 590058
rect 372954 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 373574 554614
rect 372954 554294 373574 554378
rect 372954 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 373574 554294
rect 372954 518614 373574 554058
rect 372954 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 373574 518614
rect 372954 518294 373574 518378
rect 372954 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 373574 518294
rect 372954 482614 373574 518058
rect 372954 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 373574 482614
rect 372954 482294 373574 482378
rect 372954 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 373574 482294
rect 372954 446614 373574 482058
rect 372954 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 373574 446614
rect 372954 446294 373574 446378
rect 372954 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 373574 446294
rect 372954 410614 373574 446058
rect 372954 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 373574 410614
rect 372954 410294 373574 410378
rect 372954 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 373574 410294
rect 372954 374614 373574 410058
rect 372954 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 373574 374614
rect 372954 374294 373574 374378
rect 372954 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 373574 374294
rect 372954 338614 373574 374058
rect 372954 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 373574 338614
rect 372954 338294 373574 338378
rect 372954 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 373574 338294
rect 372954 302614 373574 338058
rect 372954 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 373574 302614
rect 372954 302294 373574 302378
rect 372954 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 373574 302294
rect 372954 266614 373574 302058
rect 372954 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 373574 266614
rect 372954 266294 373574 266378
rect 372954 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 373574 266294
rect 372954 230614 373574 266058
rect 372954 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 373574 230614
rect 372954 230294 373574 230378
rect 372954 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 373574 230294
rect 372954 194614 373574 230058
rect 372954 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 373574 194614
rect 372954 194294 373574 194378
rect 372954 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 373574 194294
rect 372954 158614 373574 194058
rect 372954 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 373574 158614
rect 372954 158294 373574 158378
rect 372954 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 373574 158294
rect 372954 122614 373574 158058
rect 372954 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 373574 122614
rect 372954 122294 373574 122378
rect 372954 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 373574 122294
rect 372954 86614 373574 122058
rect 372954 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 373574 86614
rect 372954 86294 373574 86378
rect 372954 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 373574 86294
rect 372954 50614 373574 86058
rect 372954 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 373574 50614
rect 372954 50294 373574 50378
rect 372954 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 373574 50294
rect 372954 14614 373574 50058
rect 372954 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 373574 14614
rect 372954 14294 373574 14378
rect 372954 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 373574 14294
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 14058
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 669454 380414 705242
rect 379794 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 380414 669454
rect 379794 669134 380414 669218
rect 379794 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 380414 669134
rect 379794 633454 380414 668898
rect 379794 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 380414 633454
rect 379794 633134 380414 633218
rect 379794 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 380414 633134
rect 379794 597454 380414 632898
rect 379794 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 380414 597454
rect 379794 597134 380414 597218
rect 379794 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 380414 597134
rect 379794 561454 380414 596898
rect 379794 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 380414 561454
rect 379794 561134 380414 561218
rect 379794 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 380414 561134
rect 379794 525454 380414 560898
rect 379794 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 380414 525454
rect 379794 525134 380414 525218
rect 379794 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 380414 525134
rect 379794 489454 380414 524898
rect 379794 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 380414 489454
rect 379794 489134 380414 489218
rect 379794 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 380414 489134
rect 379794 453454 380414 488898
rect 379794 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 380414 453454
rect 379794 453134 380414 453218
rect 379794 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 380414 453134
rect 379794 417454 380414 452898
rect 379794 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 380414 417454
rect 379794 417134 380414 417218
rect 379794 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 380414 417134
rect 379794 381454 380414 416898
rect 379794 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 380414 381454
rect 379794 381134 380414 381218
rect 379794 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 380414 381134
rect 379794 345454 380414 380898
rect 379794 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 380414 345454
rect 379794 345134 380414 345218
rect 379794 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 380414 345134
rect 379794 309454 380414 344898
rect 379794 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 380414 309454
rect 379794 309134 380414 309218
rect 379794 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 380414 309134
rect 379794 273454 380414 308898
rect 379794 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 380414 273454
rect 379794 273134 380414 273218
rect 379794 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 380414 273134
rect 379794 237454 380414 272898
rect 379794 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 380414 237454
rect 379794 237134 380414 237218
rect 379794 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 380414 237134
rect 379794 201454 380414 236898
rect 379794 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 380414 201454
rect 379794 201134 380414 201218
rect 379794 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 380414 201134
rect 379794 165454 380414 200898
rect 379794 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 380414 165454
rect 379794 165134 380414 165218
rect 379794 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 380414 165134
rect 379794 129454 380414 164898
rect 379794 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 380414 129454
rect 379794 129134 380414 129218
rect 379794 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 380414 129134
rect 379794 93454 380414 128898
rect 379794 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 380414 93454
rect 379794 93134 380414 93218
rect 379794 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 380414 93134
rect 379794 57454 380414 92898
rect 379794 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 380414 57454
rect 379794 57134 380414 57218
rect 379794 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 380414 57134
rect 379794 21454 380414 56898
rect 379794 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 380414 21454
rect 379794 21134 380414 21218
rect 379794 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 380414 21134
rect 379794 -1306 380414 20898
rect 379794 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 380414 -1306
rect 379794 -1626 380414 -1542
rect 379794 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 380414 -1626
rect 379794 -1894 380414 -1862
rect 383514 673174 384134 707162
rect 383514 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 384134 673174
rect 383514 672854 384134 672938
rect 383514 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 384134 672854
rect 383514 637174 384134 672618
rect 383514 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 384134 637174
rect 383514 636854 384134 636938
rect 383514 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 384134 636854
rect 383514 601174 384134 636618
rect 383514 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 384134 601174
rect 383514 600854 384134 600938
rect 383514 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 384134 600854
rect 383514 565174 384134 600618
rect 383514 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 384134 565174
rect 383514 564854 384134 564938
rect 383514 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 384134 564854
rect 383514 529174 384134 564618
rect 383514 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 384134 529174
rect 383514 528854 384134 528938
rect 383514 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 384134 528854
rect 383514 493174 384134 528618
rect 383514 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 384134 493174
rect 383514 492854 384134 492938
rect 383514 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 384134 492854
rect 383514 457174 384134 492618
rect 383514 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 384134 457174
rect 383514 456854 384134 456938
rect 383514 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 384134 456854
rect 383514 421174 384134 456618
rect 383514 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 384134 421174
rect 383514 420854 384134 420938
rect 383514 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 384134 420854
rect 383514 385174 384134 420618
rect 383514 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 384134 385174
rect 383514 384854 384134 384938
rect 383514 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 384134 384854
rect 383514 349174 384134 384618
rect 383514 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 384134 349174
rect 383514 348854 384134 348938
rect 383514 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 384134 348854
rect 383514 313174 384134 348618
rect 383514 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 384134 313174
rect 383514 312854 384134 312938
rect 383514 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 384134 312854
rect 383514 277174 384134 312618
rect 383514 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 384134 277174
rect 383514 276854 384134 276938
rect 383514 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 384134 276854
rect 383514 241174 384134 276618
rect 383514 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 384134 241174
rect 383514 240854 384134 240938
rect 383514 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 384134 240854
rect 383514 205174 384134 240618
rect 383514 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 384134 205174
rect 383514 204854 384134 204938
rect 383514 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 384134 204854
rect 383514 169174 384134 204618
rect 383514 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 384134 169174
rect 383514 168854 384134 168938
rect 383514 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 384134 168854
rect 383514 133174 384134 168618
rect 383514 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 384134 133174
rect 383514 132854 384134 132938
rect 383514 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 384134 132854
rect 383514 97174 384134 132618
rect 383514 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 384134 97174
rect 383514 96854 384134 96938
rect 383514 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 384134 96854
rect 383514 61174 384134 96618
rect 383514 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 384134 61174
rect 383514 60854 384134 60938
rect 383514 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 384134 60854
rect 383514 25174 384134 60618
rect 383514 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 384134 25174
rect 383514 24854 384134 24938
rect 383514 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 384134 24854
rect 383514 -3226 384134 24618
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 676894 387854 709082
rect 387234 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 387854 676894
rect 387234 676574 387854 676658
rect 387234 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 387854 676574
rect 387234 640894 387854 676338
rect 387234 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 387854 640894
rect 387234 640574 387854 640658
rect 387234 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 387854 640574
rect 387234 604894 387854 640338
rect 387234 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 387854 604894
rect 387234 604574 387854 604658
rect 387234 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 387854 604574
rect 387234 568894 387854 604338
rect 387234 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 387854 568894
rect 387234 568574 387854 568658
rect 387234 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 387854 568574
rect 387234 532894 387854 568338
rect 387234 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 387854 532894
rect 387234 532574 387854 532658
rect 387234 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 387854 532574
rect 387234 496894 387854 532338
rect 387234 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 387854 496894
rect 387234 496574 387854 496658
rect 387234 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 387854 496574
rect 387234 460894 387854 496338
rect 387234 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 387854 460894
rect 387234 460574 387854 460658
rect 387234 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 387854 460574
rect 387234 424894 387854 460338
rect 387234 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 387854 424894
rect 387234 424574 387854 424658
rect 387234 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 387854 424574
rect 387234 388894 387854 424338
rect 387234 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 387854 388894
rect 387234 388574 387854 388658
rect 387234 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 387854 388574
rect 387234 352894 387854 388338
rect 387234 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 387854 352894
rect 387234 352574 387854 352658
rect 387234 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 387854 352574
rect 387234 316894 387854 352338
rect 387234 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 387854 316894
rect 387234 316574 387854 316658
rect 387234 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 387854 316574
rect 387234 280894 387854 316338
rect 387234 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 387854 280894
rect 387234 280574 387854 280658
rect 387234 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 387854 280574
rect 387234 244894 387854 280338
rect 387234 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 387854 244894
rect 387234 244574 387854 244658
rect 387234 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 387854 244574
rect 387234 208894 387854 244338
rect 387234 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 387854 208894
rect 387234 208574 387854 208658
rect 387234 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 387854 208574
rect 387234 172894 387854 208338
rect 387234 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 387854 172894
rect 387234 172574 387854 172658
rect 387234 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 387854 172574
rect 387234 136894 387854 172338
rect 387234 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 387854 136894
rect 387234 136574 387854 136658
rect 387234 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 387854 136574
rect 387234 100894 387854 136338
rect 387234 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 387854 100894
rect 387234 100574 387854 100658
rect 387234 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 387854 100574
rect 387234 64894 387854 100338
rect 387234 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 387854 64894
rect 387234 64574 387854 64658
rect 387234 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 387854 64574
rect 387234 28894 387854 64338
rect 387234 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 387854 28894
rect 387234 28574 387854 28658
rect 387234 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 387854 28574
rect 387234 -5146 387854 28338
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 390954 680614 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 390954 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 391574 680614
rect 390954 680294 391574 680378
rect 390954 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 391574 680294
rect 390954 644614 391574 680058
rect 390954 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 391574 644614
rect 390954 644294 391574 644378
rect 390954 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 391574 644294
rect 390954 608614 391574 644058
rect 390954 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 391574 608614
rect 390954 608294 391574 608378
rect 390954 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 391574 608294
rect 390954 572614 391574 608058
rect 390954 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 391574 572614
rect 390954 572294 391574 572378
rect 390954 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 391574 572294
rect 390954 536614 391574 572058
rect 390954 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 391574 536614
rect 390954 536294 391574 536378
rect 390954 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 391574 536294
rect 390954 500614 391574 536058
rect 390954 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 391574 500614
rect 390954 500294 391574 500378
rect 390954 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 391574 500294
rect 390954 464614 391574 500058
rect 390954 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 391574 464614
rect 390954 464294 391574 464378
rect 390954 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 391574 464294
rect 390954 428614 391574 464058
rect 390954 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 391574 428614
rect 390954 428294 391574 428378
rect 390954 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 391574 428294
rect 390954 392614 391574 428058
rect 390954 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 391574 392614
rect 390954 392294 391574 392378
rect 390954 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 391574 392294
rect 390954 356614 391574 392058
rect 390954 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 391574 356614
rect 390954 356294 391574 356378
rect 390954 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 391574 356294
rect 390954 320614 391574 356058
rect 390954 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 391574 320614
rect 390954 320294 391574 320378
rect 390954 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 391574 320294
rect 390954 284614 391574 320058
rect 390954 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 391574 284614
rect 390954 284294 391574 284378
rect 390954 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 391574 284294
rect 390954 248614 391574 284058
rect 390954 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 391574 248614
rect 390954 248294 391574 248378
rect 390954 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 391574 248294
rect 390954 212614 391574 248058
rect 390954 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 391574 212614
rect 390954 212294 391574 212378
rect 390954 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 391574 212294
rect 390954 176614 391574 212058
rect 390954 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 391574 176614
rect 390954 176294 391574 176378
rect 390954 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 391574 176294
rect 390954 140614 391574 176058
rect 390954 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 391574 140614
rect 390954 140294 391574 140378
rect 390954 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 391574 140294
rect 390954 104614 391574 140058
rect 390954 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 391574 104614
rect 390954 104294 391574 104378
rect 390954 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 391574 104294
rect 390954 68614 391574 104058
rect 390954 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 391574 68614
rect 390954 68294 391574 68378
rect 390954 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 391574 68294
rect 390954 32614 391574 68058
rect 390954 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 391574 32614
rect 390954 32294 391574 32378
rect 390954 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 391574 32294
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 32058
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 687454 398414 704282
rect 397794 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 398414 687454
rect 397794 687134 398414 687218
rect 397794 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 398414 687134
rect 397794 651454 398414 686898
rect 397794 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 398414 651454
rect 397794 651134 398414 651218
rect 397794 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 398414 651134
rect 397794 615454 398414 650898
rect 397794 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 398414 615454
rect 397794 615134 398414 615218
rect 397794 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 398414 615134
rect 397794 579454 398414 614898
rect 397794 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 398414 579454
rect 397794 579134 398414 579218
rect 397794 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 398414 579134
rect 397794 543454 398414 578898
rect 397794 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 398414 543454
rect 397794 543134 398414 543218
rect 397794 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 398414 543134
rect 397794 507454 398414 542898
rect 397794 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 398414 507454
rect 397794 507134 398414 507218
rect 397794 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 398414 507134
rect 397794 471454 398414 506898
rect 397794 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 398414 471454
rect 397794 471134 398414 471218
rect 397794 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 398414 471134
rect 397794 435454 398414 470898
rect 397794 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 398414 435454
rect 397794 435134 398414 435218
rect 397794 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 398414 435134
rect 397794 399454 398414 434898
rect 397794 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 398414 399454
rect 397794 399134 398414 399218
rect 397794 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 398414 399134
rect 397794 363454 398414 398898
rect 397794 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 398414 363454
rect 397794 363134 398414 363218
rect 397794 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 398414 363134
rect 397794 327454 398414 362898
rect 397794 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 398414 327454
rect 397794 327134 398414 327218
rect 397794 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 398414 327134
rect 397794 291454 398414 326898
rect 397794 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 398414 291454
rect 397794 291134 398414 291218
rect 397794 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 398414 291134
rect 397794 255454 398414 290898
rect 397794 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 398414 255454
rect 397794 255134 398414 255218
rect 397794 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 398414 255134
rect 397794 219454 398414 254898
rect 397794 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 398414 219454
rect 397794 219134 398414 219218
rect 397794 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 398414 219134
rect 397794 183454 398414 218898
rect 397794 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 398414 183454
rect 397794 183134 398414 183218
rect 397794 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 398414 183134
rect 397794 147454 398414 182898
rect 397794 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 398414 147454
rect 397794 147134 398414 147218
rect 397794 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 398414 147134
rect 397794 111454 398414 146898
rect 397794 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 398414 111454
rect 397794 111134 398414 111218
rect 397794 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 398414 111134
rect 397794 75454 398414 110898
rect 397794 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 398414 75454
rect 397794 75134 398414 75218
rect 397794 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 398414 75134
rect 397794 39454 398414 74898
rect 397794 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 398414 39454
rect 397794 39134 398414 39218
rect 397794 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 398414 39134
rect 397794 3454 398414 38898
rect 397794 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 398414 3454
rect 397794 3134 398414 3218
rect 397794 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 398414 3134
rect 397794 -346 398414 2898
rect 397794 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 398414 -346
rect 397794 -666 398414 -582
rect 397794 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 398414 -666
rect 397794 -1894 398414 -902
rect 401514 691174 402134 706202
rect 401514 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 402134 691174
rect 401514 690854 402134 690938
rect 401514 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 402134 690854
rect 401514 655174 402134 690618
rect 401514 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 402134 655174
rect 401514 654854 402134 654938
rect 401514 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 402134 654854
rect 401514 619174 402134 654618
rect 401514 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 402134 619174
rect 401514 618854 402134 618938
rect 401514 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 402134 618854
rect 401514 583174 402134 618618
rect 401514 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 402134 583174
rect 401514 582854 402134 582938
rect 401514 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 402134 582854
rect 401514 547174 402134 582618
rect 401514 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 402134 547174
rect 401514 546854 402134 546938
rect 401514 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 402134 546854
rect 401514 511174 402134 546618
rect 401514 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 402134 511174
rect 401514 510854 402134 510938
rect 401514 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 402134 510854
rect 401514 475174 402134 510618
rect 401514 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 402134 475174
rect 401514 474854 402134 474938
rect 401514 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 402134 474854
rect 401514 439174 402134 474618
rect 401514 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 402134 439174
rect 401514 438854 402134 438938
rect 401514 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 402134 438854
rect 401514 403174 402134 438618
rect 401514 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 402134 403174
rect 401514 402854 402134 402938
rect 401514 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 402134 402854
rect 401514 367174 402134 402618
rect 401514 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 402134 367174
rect 401514 366854 402134 366938
rect 401514 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 402134 366854
rect 401514 331174 402134 366618
rect 401514 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 402134 331174
rect 401514 330854 402134 330938
rect 401514 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 402134 330854
rect 401514 295174 402134 330618
rect 401514 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 402134 295174
rect 401514 294854 402134 294938
rect 401514 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 402134 294854
rect 401514 259174 402134 294618
rect 401514 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 402134 259174
rect 401514 258854 402134 258938
rect 401514 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 402134 258854
rect 401514 223174 402134 258618
rect 401514 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 402134 223174
rect 401514 222854 402134 222938
rect 401514 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 402134 222854
rect 401514 187174 402134 222618
rect 401514 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 402134 187174
rect 401514 186854 402134 186938
rect 401514 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 402134 186854
rect 401514 151174 402134 186618
rect 401514 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 402134 151174
rect 401514 150854 402134 150938
rect 401514 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 402134 150854
rect 401514 115174 402134 150618
rect 401514 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 402134 115174
rect 401514 114854 402134 114938
rect 401514 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 402134 114854
rect 401514 79174 402134 114618
rect 401514 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 402134 79174
rect 401514 78854 402134 78938
rect 401514 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 402134 78854
rect 401514 43174 402134 78618
rect 401514 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 402134 43174
rect 401514 42854 402134 42938
rect 401514 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 402134 42854
rect 401514 7174 402134 42618
rect 401514 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 402134 7174
rect 401514 6854 402134 6938
rect 401514 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 402134 6854
rect 401514 -2266 402134 6618
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 694894 405854 708122
rect 405234 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 405854 694894
rect 405234 694574 405854 694658
rect 405234 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 405854 694574
rect 405234 658894 405854 694338
rect 405234 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 405854 658894
rect 405234 658574 405854 658658
rect 405234 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 405854 658574
rect 405234 622894 405854 658338
rect 405234 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 405854 622894
rect 405234 622574 405854 622658
rect 405234 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 405854 622574
rect 405234 586894 405854 622338
rect 405234 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 405854 586894
rect 405234 586574 405854 586658
rect 405234 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 405854 586574
rect 405234 550894 405854 586338
rect 405234 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 405854 550894
rect 405234 550574 405854 550658
rect 405234 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 405854 550574
rect 405234 514894 405854 550338
rect 405234 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 405854 514894
rect 405234 514574 405854 514658
rect 405234 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 405854 514574
rect 405234 478894 405854 514338
rect 405234 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 405854 478894
rect 405234 478574 405854 478658
rect 405234 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 405854 478574
rect 405234 442894 405854 478338
rect 405234 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 405854 442894
rect 405234 442574 405854 442658
rect 405234 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 405854 442574
rect 405234 406894 405854 442338
rect 405234 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 405854 406894
rect 405234 406574 405854 406658
rect 405234 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 405854 406574
rect 405234 370894 405854 406338
rect 405234 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 405854 370894
rect 405234 370574 405854 370658
rect 405234 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 405854 370574
rect 405234 334894 405854 370338
rect 405234 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 405854 334894
rect 405234 334574 405854 334658
rect 405234 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 405854 334574
rect 405234 298894 405854 334338
rect 405234 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 405854 298894
rect 405234 298574 405854 298658
rect 405234 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 405854 298574
rect 405234 262894 405854 298338
rect 405234 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 405854 262894
rect 405234 262574 405854 262658
rect 405234 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 405854 262574
rect 405234 226894 405854 262338
rect 405234 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 405854 226894
rect 405234 226574 405854 226658
rect 405234 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 405854 226574
rect 405234 190894 405854 226338
rect 405234 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 405854 190894
rect 405234 190574 405854 190658
rect 405234 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 405854 190574
rect 405234 154894 405854 190338
rect 405234 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 405854 154894
rect 405234 154574 405854 154658
rect 405234 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 405854 154574
rect 405234 118894 405854 154338
rect 405234 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 405854 118894
rect 405234 118574 405854 118658
rect 405234 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 405854 118574
rect 405234 82894 405854 118338
rect 405234 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 405854 82894
rect 405234 82574 405854 82658
rect 405234 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 405854 82574
rect 405234 46894 405854 82338
rect 405234 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 405854 46894
rect 405234 46574 405854 46658
rect 405234 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 405854 46574
rect 405234 10894 405854 46338
rect 405234 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 405854 10894
rect 405234 10574 405854 10658
rect 405234 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 405854 10574
rect 405234 -4186 405854 10338
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 408954 698614 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 408954 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 409574 698614
rect 408954 698294 409574 698378
rect 408954 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 409574 698294
rect 408954 662614 409574 698058
rect 408954 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 409574 662614
rect 408954 662294 409574 662378
rect 408954 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 409574 662294
rect 408954 626614 409574 662058
rect 408954 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 409574 626614
rect 408954 626294 409574 626378
rect 408954 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 409574 626294
rect 408954 590614 409574 626058
rect 408954 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 409574 590614
rect 408954 590294 409574 590378
rect 408954 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 409574 590294
rect 408954 554614 409574 590058
rect 408954 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 409574 554614
rect 408954 554294 409574 554378
rect 408954 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 409574 554294
rect 408954 518614 409574 554058
rect 408954 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 409574 518614
rect 408954 518294 409574 518378
rect 408954 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 409574 518294
rect 408954 482614 409574 518058
rect 408954 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 409574 482614
rect 408954 482294 409574 482378
rect 408954 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 409574 482294
rect 408954 446614 409574 482058
rect 408954 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 409574 446614
rect 408954 446294 409574 446378
rect 408954 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 409574 446294
rect 408954 410614 409574 446058
rect 408954 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 409574 410614
rect 408954 410294 409574 410378
rect 408954 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 409574 410294
rect 408954 374614 409574 410058
rect 408954 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 409574 374614
rect 408954 374294 409574 374378
rect 408954 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 409574 374294
rect 408954 338614 409574 374058
rect 408954 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 409574 338614
rect 408954 338294 409574 338378
rect 408954 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 409574 338294
rect 408954 302614 409574 338058
rect 408954 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 409574 302614
rect 408954 302294 409574 302378
rect 408954 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 409574 302294
rect 408954 266614 409574 302058
rect 408954 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 409574 266614
rect 408954 266294 409574 266378
rect 408954 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 409574 266294
rect 408954 230614 409574 266058
rect 408954 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 409574 230614
rect 408954 230294 409574 230378
rect 408954 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 409574 230294
rect 408954 194614 409574 230058
rect 408954 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 409574 194614
rect 408954 194294 409574 194378
rect 408954 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 409574 194294
rect 408954 158614 409574 194058
rect 408954 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 409574 158614
rect 408954 158294 409574 158378
rect 408954 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 409574 158294
rect 408954 122614 409574 158058
rect 408954 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 409574 122614
rect 408954 122294 409574 122378
rect 408954 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 409574 122294
rect 408954 86614 409574 122058
rect 408954 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 409574 86614
rect 408954 86294 409574 86378
rect 408954 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 409574 86294
rect 408954 50614 409574 86058
rect 408954 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 409574 50614
rect 408954 50294 409574 50378
rect 408954 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 409574 50294
rect 408954 14614 409574 50058
rect 408954 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 409574 14614
rect 408954 14294 409574 14378
rect 408954 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 409574 14294
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 14058
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 669454 416414 705242
rect 415794 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 416414 669454
rect 415794 669134 416414 669218
rect 415794 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 416414 669134
rect 415794 633454 416414 668898
rect 415794 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 416414 633454
rect 415794 633134 416414 633218
rect 415794 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 416414 633134
rect 415794 597454 416414 632898
rect 415794 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 416414 597454
rect 415794 597134 416414 597218
rect 415794 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 416414 597134
rect 415794 561454 416414 596898
rect 415794 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 416414 561454
rect 415794 561134 416414 561218
rect 415794 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 416414 561134
rect 415794 525454 416414 560898
rect 415794 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 416414 525454
rect 415794 525134 416414 525218
rect 415794 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 416414 525134
rect 415794 489454 416414 524898
rect 415794 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 416414 489454
rect 415794 489134 416414 489218
rect 415794 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 416414 489134
rect 415794 453454 416414 488898
rect 415794 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 416414 453454
rect 415794 453134 416414 453218
rect 415794 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 416414 453134
rect 415794 417454 416414 452898
rect 415794 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 416414 417454
rect 415794 417134 416414 417218
rect 415794 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 416414 417134
rect 415794 381454 416414 416898
rect 415794 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 416414 381454
rect 415794 381134 416414 381218
rect 415794 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 416414 381134
rect 415794 345454 416414 380898
rect 415794 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 416414 345454
rect 415794 345134 416414 345218
rect 415794 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 416414 345134
rect 415794 309454 416414 344898
rect 415794 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 416414 309454
rect 415794 309134 416414 309218
rect 415794 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 416414 309134
rect 415794 273454 416414 308898
rect 415794 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 416414 273454
rect 415794 273134 416414 273218
rect 415794 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 416414 273134
rect 415794 237454 416414 272898
rect 415794 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 416414 237454
rect 415794 237134 416414 237218
rect 415794 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 416414 237134
rect 415794 201454 416414 236898
rect 415794 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 416414 201454
rect 415794 201134 416414 201218
rect 415794 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 416414 201134
rect 415794 165454 416414 200898
rect 415794 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 416414 165454
rect 415794 165134 416414 165218
rect 415794 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 416414 165134
rect 415794 129454 416414 164898
rect 415794 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 416414 129454
rect 415794 129134 416414 129218
rect 415794 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 416414 129134
rect 415794 93454 416414 128898
rect 415794 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 416414 93454
rect 415794 93134 416414 93218
rect 415794 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 416414 93134
rect 415794 57454 416414 92898
rect 415794 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 416414 57454
rect 415794 57134 416414 57218
rect 415794 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 416414 57134
rect 415794 21454 416414 56898
rect 415794 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 416414 21454
rect 415794 21134 416414 21218
rect 415794 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 416414 21134
rect 415794 -1306 416414 20898
rect 415794 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 416414 -1306
rect 415794 -1626 416414 -1542
rect 415794 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 416414 -1626
rect 415794 -1894 416414 -1862
rect 419514 673174 420134 707162
rect 419514 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 420134 673174
rect 419514 672854 420134 672938
rect 419514 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 420134 672854
rect 419514 637174 420134 672618
rect 419514 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 420134 637174
rect 419514 636854 420134 636938
rect 419514 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 420134 636854
rect 419514 601174 420134 636618
rect 419514 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 420134 601174
rect 419514 600854 420134 600938
rect 419514 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 420134 600854
rect 419514 565174 420134 600618
rect 419514 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 420134 565174
rect 419514 564854 420134 564938
rect 419514 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 420134 564854
rect 419514 529174 420134 564618
rect 419514 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 420134 529174
rect 419514 528854 420134 528938
rect 419514 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 420134 528854
rect 419514 493174 420134 528618
rect 419514 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 420134 493174
rect 419514 492854 420134 492938
rect 419514 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 420134 492854
rect 419514 457174 420134 492618
rect 419514 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 420134 457174
rect 419514 456854 420134 456938
rect 419514 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 420134 456854
rect 419514 421174 420134 456618
rect 419514 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 420134 421174
rect 419514 420854 420134 420938
rect 419514 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 420134 420854
rect 419514 385174 420134 420618
rect 419514 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 420134 385174
rect 419514 384854 420134 384938
rect 419514 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 420134 384854
rect 419514 349174 420134 384618
rect 419514 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 420134 349174
rect 419514 348854 420134 348938
rect 419514 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 420134 348854
rect 419514 313174 420134 348618
rect 419514 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 420134 313174
rect 419514 312854 420134 312938
rect 419514 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 420134 312854
rect 419514 277174 420134 312618
rect 419514 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 420134 277174
rect 419514 276854 420134 276938
rect 419514 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 420134 276854
rect 419514 241174 420134 276618
rect 419514 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 420134 241174
rect 419514 240854 420134 240938
rect 419514 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 420134 240854
rect 419514 205174 420134 240618
rect 419514 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 420134 205174
rect 419514 204854 420134 204938
rect 419514 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 420134 204854
rect 419514 169174 420134 204618
rect 419514 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 420134 169174
rect 419514 168854 420134 168938
rect 419514 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 420134 168854
rect 419514 133174 420134 168618
rect 419514 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 420134 133174
rect 419514 132854 420134 132938
rect 419514 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 420134 132854
rect 419514 97174 420134 132618
rect 419514 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 420134 97174
rect 419514 96854 420134 96938
rect 419514 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 420134 96854
rect 419514 61174 420134 96618
rect 419514 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 420134 61174
rect 419514 60854 420134 60938
rect 419514 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 420134 60854
rect 419514 25174 420134 60618
rect 419514 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 420134 25174
rect 419514 24854 420134 24938
rect 419514 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 420134 24854
rect 419514 -3226 420134 24618
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 676894 423854 709082
rect 423234 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 423854 676894
rect 423234 676574 423854 676658
rect 423234 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 423854 676574
rect 423234 640894 423854 676338
rect 423234 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 423854 640894
rect 423234 640574 423854 640658
rect 423234 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 423854 640574
rect 423234 604894 423854 640338
rect 423234 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 423854 604894
rect 423234 604574 423854 604658
rect 423234 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 423854 604574
rect 423234 568894 423854 604338
rect 423234 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 423854 568894
rect 423234 568574 423854 568658
rect 423234 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 423854 568574
rect 423234 532894 423854 568338
rect 423234 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 423854 532894
rect 423234 532574 423854 532658
rect 423234 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 423854 532574
rect 423234 496894 423854 532338
rect 423234 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 423854 496894
rect 423234 496574 423854 496658
rect 423234 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 423854 496574
rect 423234 460894 423854 496338
rect 423234 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 423854 460894
rect 423234 460574 423854 460658
rect 423234 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 423854 460574
rect 423234 424894 423854 460338
rect 423234 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 423854 424894
rect 423234 424574 423854 424658
rect 423234 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 423854 424574
rect 423234 388894 423854 424338
rect 423234 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 423854 388894
rect 423234 388574 423854 388658
rect 423234 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 423854 388574
rect 423234 352894 423854 388338
rect 423234 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 423854 352894
rect 423234 352574 423854 352658
rect 423234 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 423854 352574
rect 423234 316894 423854 352338
rect 423234 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 423854 316894
rect 423234 316574 423854 316658
rect 423234 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 423854 316574
rect 423234 280894 423854 316338
rect 423234 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 423854 280894
rect 423234 280574 423854 280658
rect 423234 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 423854 280574
rect 423234 244894 423854 280338
rect 423234 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 423854 244894
rect 423234 244574 423854 244658
rect 423234 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 423854 244574
rect 423234 208894 423854 244338
rect 423234 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 423854 208894
rect 423234 208574 423854 208658
rect 423234 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 423854 208574
rect 423234 172894 423854 208338
rect 423234 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 423854 172894
rect 423234 172574 423854 172658
rect 423234 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 423854 172574
rect 423234 136894 423854 172338
rect 423234 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 423854 136894
rect 423234 136574 423854 136658
rect 423234 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 423854 136574
rect 423234 100894 423854 136338
rect 423234 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 423854 100894
rect 423234 100574 423854 100658
rect 423234 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 423854 100574
rect 423234 64894 423854 100338
rect 423234 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 423854 64894
rect 423234 64574 423854 64658
rect 423234 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 423854 64574
rect 423234 28894 423854 64338
rect 423234 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 423854 28894
rect 423234 28574 423854 28658
rect 423234 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 423854 28574
rect 423234 -5146 423854 28338
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 426954 680614 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 426954 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 427574 680614
rect 426954 680294 427574 680378
rect 426954 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 427574 680294
rect 426954 644614 427574 680058
rect 426954 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 427574 644614
rect 426954 644294 427574 644378
rect 426954 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 427574 644294
rect 426954 608614 427574 644058
rect 426954 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 427574 608614
rect 426954 608294 427574 608378
rect 426954 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 427574 608294
rect 426954 572614 427574 608058
rect 426954 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 427574 572614
rect 426954 572294 427574 572378
rect 426954 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 427574 572294
rect 426954 536614 427574 572058
rect 426954 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 427574 536614
rect 426954 536294 427574 536378
rect 426954 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 427574 536294
rect 426954 500614 427574 536058
rect 426954 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 427574 500614
rect 426954 500294 427574 500378
rect 426954 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 427574 500294
rect 426954 464614 427574 500058
rect 426954 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 427574 464614
rect 426954 464294 427574 464378
rect 426954 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 427574 464294
rect 426954 428614 427574 464058
rect 426954 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 427574 428614
rect 426954 428294 427574 428378
rect 426954 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 427574 428294
rect 426954 392614 427574 428058
rect 426954 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 427574 392614
rect 426954 392294 427574 392378
rect 426954 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 427574 392294
rect 426954 356614 427574 392058
rect 426954 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 427574 356614
rect 426954 356294 427574 356378
rect 426954 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 427574 356294
rect 426954 320614 427574 356058
rect 426954 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 427574 320614
rect 426954 320294 427574 320378
rect 426954 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 427574 320294
rect 426954 284614 427574 320058
rect 426954 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 427574 284614
rect 426954 284294 427574 284378
rect 426954 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 427574 284294
rect 426954 248614 427574 284058
rect 426954 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 427574 248614
rect 426954 248294 427574 248378
rect 426954 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 427574 248294
rect 426954 212614 427574 248058
rect 426954 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 427574 212614
rect 426954 212294 427574 212378
rect 426954 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 427574 212294
rect 426954 176614 427574 212058
rect 426954 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 427574 176614
rect 426954 176294 427574 176378
rect 426954 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 427574 176294
rect 426954 140614 427574 176058
rect 426954 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 427574 140614
rect 426954 140294 427574 140378
rect 426954 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 427574 140294
rect 426954 104614 427574 140058
rect 426954 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 427574 104614
rect 426954 104294 427574 104378
rect 426954 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 427574 104294
rect 426954 68614 427574 104058
rect 426954 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 427574 68614
rect 426954 68294 427574 68378
rect 426954 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 427574 68294
rect 426954 32614 427574 68058
rect 426954 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 427574 32614
rect 426954 32294 427574 32378
rect 426954 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 427574 32294
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 32058
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 687454 434414 704282
rect 433794 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 434414 687454
rect 433794 687134 434414 687218
rect 433794 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 434414 687134
rect 433794 651454 434414 686898
rect 433794 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 434414 651454
rect 433794 651134 434414 651218
rect 433794 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 434414 651134
rect 433794 615454 434414 650898
rect 433794 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 434414 615454
rect 433794 615134 434414 615218
rect 433794 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 434414 615134
rect 433794 579454 434414 614898
rect 433794 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 434414 579454
rect 433794 579134 434414 579218
rect 433794 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 434414 579134
rect 433794 543454 434414 578898
rect 433794 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 434414 543454
rect 433794 543134 434414 543218
rect 433794 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 434414 543134
rect 433794 507454 434414 542898
rect 433794 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 434414 507454
rect 433794 507134 434414 507218
rect 433794 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 434414 507134
rect 433794 471454 434414 506898
rect 433794 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 434414 471454
rect 433794 471134 434414 471218
rect 433794 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 434414 471134
rect 433794 435454 434414 470898
rect 433794 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 434414 435454
rect 433794 435134 434414 435218
rect 433794 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 434414 435134
rect 433794 399454 434414 434898
rect 433794 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 434414 399454
rect 433794 399134 434414 399218
rect 433794 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 434414 399134
rect 433794 363454 434414 398898
rect 433794 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 434414 363454
rect 433794 363134 434414 363218
rect 433794 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 434414 363134
rect 433794 327454 434414 362898
rect 433794 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 434414 327454
rect 433794 327134 434414 327218
rect 433794 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 434414 327134
rect 433794 291454 434414 326898
rect 433794 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 434414 291454
rect 433794 291134 434414 291218
rect 433794 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 434414 291134
rect 433794 255454 434414 290898
rect 433794 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 434414 255454
rect 433794 255134 434414 255218
rect 433794 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 434414 255134
rect 433794 219454 434414 254898
rect 433794 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 434414 219454
rect 433794 219134 434414 219218
rect 433794 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 434414 219134
rect 433794 183454 434414 218898
rect 433794 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 434414 183454
rect 433794 183134 434414 183218
rect 433794 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 434414 183134
rect 433794 147454 434414 182898
rect 433794 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 434414 147454
rect 433794 147134 434414 147218
rect 433794 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 434414 147134
rect 433794 111454 434414 146898
rect 433794 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 434414 111454
rect 433794 111134 434414 111218
rect 433794 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 434414 111134
rect 433794 75454 434414 110898
rect 433794 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 434414 75454
rect 433794 75134 434414 75218
rect 433794 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 434414 75134
rect 433794 39454 434414 74898
rect 433794 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 434414 39454
rect 433794 39134 434414 39218
rect 433794 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 434414 39134
rect 433794 3454 434414 38898
rect 433794 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 434414 3454
rect 433794 3134 434414 3218
rect 433794 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 434414 3134
rect 433794 -346 434414 2898
rect 433794 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 434414 -346
rect 433794 -666 434414 -582
rect 433794 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 434414 -666
rect 433794 -1894 434414 -902
rect 437514 691174 438134 706202
rect 437514 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 438134 691174
rect 437514 690854 438134 690938
rect 437514 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 438134 690854
rect 437514 655174 438134 690618
rect 437514 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 438134 655174
rect 437514 654854 438134 654938
rect 437514 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 438134 654854
rect 437514 619174 438134 654618
rect 437514 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 438134 619174
rect 437514 618854 438134 618938
rect 437514 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 438134 618854
rect 437514 583174 438134 618618
rect 437514 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 438134 583174
rect 437514 582854 438134 582938
rect 437514 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 438134 582854
rect 437514 547174 438134 582618
rect 437514 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 438134 547174
rect 437514 546854 438134 546938
rect 437514 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 438134 546854
rect 437514 511174 438134 546618
rect 437514 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 438134 511174
rect 437514 510854 438134 510938
rect 437514 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 438134 510854
rect 437514 475174 438134 510618
rect 437514 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 438134 475174
rect 437514 474854 438134 474938
rect 437514 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 438134 474854
rect 437514 439174 438134 474618
rect 437514 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 438134 439174
rect 437514 438854 438134 438938
rect 437514 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 438134 438854
rect 437514 403174 438134 438618
rect 437514 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 438134 403174
rect 437514 402854 438134 402938
rect 437514 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 438134 402854
rect 437514 367174 438134 402618
rect 437514 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 438134 367174
rect 437514 366854 438134 366938
rect 437514 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 438134 366854
rect 437514 331174 438134 366618
rect 437514 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 438134 331174
rect 437514 330854 438134 330938
rect 437514 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 438134 330854
rect 437514 295174 438134 330618
rect 437514 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 438134 295174
rect 437514 294854 438134 294938
rect 437514 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 438134 294854
rect 437514 259174 438134 294618
rect 437514 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 438134 259174
rect 437514 258854 438134 258938
rect 437514 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 438134 258854
rect 437514 223174 438134 258618
rect 437514 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 438134 223174
rect 437514 222854 438134 222938
rect 437514 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 438134 222854
rect 437514 187174 438134 222618
rect 437514 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 438134 187174
rect 437514 186854 438134 186938
rect 437514 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 438134 186854
rect 437514 151174 438134 186618
rect 437514 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 438134 151174
rect 437514 150854 438134 150938
rect 437514 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 438134 150854
rect 437514 115174 438134 150618
rect 437514 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 438134 115174
rect 437514 114854 438134 114938
rect 437514 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 438134 114854
rect 437514 79174 438134 114618
rect 437514 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 438134 79174
rect 437514 78854 438134 78938
rect 437514 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 438134 78854
rect 437514 43174 438134 78618
rect 437514 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 438134 43174
rect 437514 42854 438134 42938
rect 437514 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 438134 42854
rect 437514 7174 438134 42618
rect 437514 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 438134 7174
rect 437514 6854 438134 6938
rect 437514 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 438134 6854
rect 437514 -2266 438134 6618
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 694894 441854 708122
rect 441234 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 441854 694894
rect 441234 694574 441854 694658
rect 441234 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 441854 694574
rect 441234 658894 441854 694338
rect 441234 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 441854 658894
rect 441234 658574 441854 658658
rect 441234 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 441854 658574
rect 441234 622894 441854 658338
rect 441234 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 441854 622894
rect 441234 622574 441854 622658
rect 441234 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 441854 622574
rect 441234 586894 441854 622338
rect 441234 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 441854 586894
rect 441234 586574 441854 586658
rect 441234 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 441854 586574
rect 441234 550894 441854 586338
rect 441234 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 441854 550894
rect 441234 550574 441854 550658
rect 441234 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 441854 550574
rect 441234 514894 441854 550338
rect 441234 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 441854 514894
rect 441234 514574 441854 514658
rect 441234 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 441854 514574
rect 441234 478894 441854 514338
rect 441234 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 441854 478894
rect 441234 478574 441854 478658
rect 441234 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 441854 478574
rect 441234 442894 441854 478338
rect 441234 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 441854 442894
rect 441234 442574 441854 442658
rect 441234 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 441854 442574
rect 441234 406894 441854 442338
rect 441234 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 441854 406894
rect 441234 406574 441854 406658
rect 441234 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 441854 406574
rect 441234 370894 441854 406338
rect 441234 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 441854 370894
rect 441234 370574 441854 370658
rect 441234 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 441854 370574
rect 441234 334894 441854 370338
rect 441234 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 441854 334894
rect 441234 334574 441854 334658
rect 441234 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 441854 334574
rect 441234 298894 441854 334338
rect 441234 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 441854 298894
rect 441234 298574 441854 298658
rect 441234 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 441854 298574
rect 441234 262894 441854 298338
rect 441234 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 441854 262894
rect 441234 262574 441854 262658
rect 441234 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 441854 262574
rect 441234 226894 441854 262338
rect 441234 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 441854 226894
rect 441234 226574 441854 226658
rect 441234 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 441854 226574
rect 441234 190894 441854 226338
rect 441234 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 441854 190894
rect 441234 190574 441854 190658
rect 441234 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 441854 190574
rect 441234 154894 441854 190338
rect 441234 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 441854 154894
rect 441234 154574 441854 154658
rect 441234 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 441854 154574
rect 441234 118894 441854 154338
rect 441234 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 441854 118894
rect 441234 118574 441854 118658
rect 441234 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 441854 118574
rect 441234 82894 441854 118338
rect 441234 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 441854 82894
rect 441234 82574 441854 82658
rect 441234 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 441854 82574
rect 441234 46894 441854 82338
rect 441234 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 441854 46894
rect 441234 46574 441854 46658
rect 441234 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 441854 46574
rect 441234 10894 441854 46338
rect 441234 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 441854 10894
rect 441234 10574 441854 10658
rect 441234 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 441854 10574
rect 441234 -4186 441854 10338
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 444954 698614 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 444954 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 445574 698614
rect 444954 698294 445574 698378
rect 444954 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 445574 698294
rect 444954 662614 445574 698058
rect 444954 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 445574 662614
rect 444954 662294 445574 662378
rect 444954 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 445574 662294
rect 444954 626614 445574 662058
rect 444954 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 445574 626614
rect 444954 626294 445574 626378
rect 444954 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 445574 626294
rect 444954 590614 445574 626058
rect 444954 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 445574 590614
rect 444954 590294 445574 590378
rect 444954 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 445574 590294
rect 444954 554614 445574 590058
rect 444954 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 445574 554614
rect 444954 554294 445574 554378
rect 444954 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 445574 554294
rect 444954 518614 445574 554058
rect 444954 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 445574 518614
rect 444954 518294 445574 518378
rect 444954 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 445574 518294
rect 444954 482614 445574 518058
rect 444954 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 445574 482614
rect 444954 482294 445574 482378
rect 444954 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 445574 482294
rect 444954 446614 445574 482058
rect 444954 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 445574 446614
rect 444954 446294 445574 446378
rect 444954 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 445574 446294
rect 444954 410614 445574 446058
rect 444954 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 445574 410614
rect 444954 410294 445574 410378
rect 444954 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 445574 410294
rect 444954 374614 445574 410058
rect 444954 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 445574 374614
rect 444954 374294 445574 374378
rect 444954 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 445574 374294
rect 444954 338614 445574 374058
rect 444954 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 445574 338614
rect 444954 338294 445574 338378
rect 444954 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 445574 338294
rect 444954 302614 445574 338058
rect 444954 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 445574 302614
rect 444954 302294 445574 302378
rect 444954 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 445574 302294
rect 444954 266614 445574 302058
rect 444954 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 445574 266614
rect 444954 266294 445574 266378
rect 444954 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 445574 266294
rect 444954 230614 445574 266058
rect 444954 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 445574 230614
rect 444954 230294 445574 230378
rect 444954 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 445574 230294
rect 444954 194614 445574 230058
rect 444954 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 445574 194614
rect 444954 194294 445574 194378
rect 444954 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 445574 194294
rect 444954 158614 445574 194058
rect 444954 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 445574 158614
rect 444954 158294 445574 158378
rect 444954 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 445574 158294
rect 444954 122614 445574 158058
rect 444954 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 445574 122614
rect 444954 122294 445574 122378
rect 444954 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 445574 122294
rect 444954 86614 445574 122058
rect 444954 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 445574 86614
rect 444954 86294 445574 86378
rect 444954 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 445574 86294
rect 444954 50614 445574 86058
rect 444954 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 445574 50614
rect 444954 50294 445574 50378
rect 444954 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 445574 50294
rect 444954 14614 445574 50058
rect 444954 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 445574 14614
rect 444954 14294 445574 14378
rect 444954 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 445574 14294
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 14058
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 669454 452414 705242
rect 451794 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 452414 669454
rect 451794 669134 452414 669218
rect 451794 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 452414 669134
rect 451794 633454 452414 668898
rect 451794 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 452414 633454
rect 451794 633134 452414 633218
rect 451794 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 452414 633134
rect 451794 597454 452414 632898
rect 451794 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 452414 597454
rect 451794 597134 452414 597218
rect 451794 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 452414 597134
rect 451794 561454 452414 596898
rect 451794 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 452414 561454
rect 451794 561134 452414 561218
rect 451794 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 452414 561134
rect 451794 525454 452414 560898
rect 451794 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 452414 525454
rect 451794 525134 452414 525218
rect 451794 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 452414 525134
rect 451794 489454 452414 524898
rect 451794 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 452414 489454
rect 451794 489134 452414 489218
rect 451794 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 452414 489134
rect 451794 453454 452414 488898
rect 451794 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 452414 453454
rect 451794 453134 452414 453218
rect 451794 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 452414 453134
rect 451794 417454 452414 452898
rect 451794 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 452414 417454
rect 451794 417134 452414 417218
rect 451794 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 452414 417134
rect 451794 381454 452414 416898
rect 451794 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 452414 381454
rect 451794 381134 452414 381218
rect 451794 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 452414 381134
rect 451794 345454 452414 380898
rect 451794 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 452414 345454
rect 451794 345134 452414 345218
rect 451794 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 452414 345134
rect 451794 309454 452414 344898
rect 451794 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 452414 309454
rect 451794 309134 452414 309218
rect 451794 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 452414 309134
rect 451794 273454 452414 308898
rect 451794 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 452414 273454
rect 451794 273134 452414 273218
rect 451794 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 452414 273134
rect 451794 237454 452414 272898
rect 451794 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 452414 237454
rect 451794 237134 452414 237218
rect 451794 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 452414 237134
rect 451794 201454 452414 236898
rect 451794 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 452414 201454
rect 451794 201134 452414 201218
rect 451794 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 452414 201134
rect 451794 165454 452414 200898
rect 451794 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 452414 165454
rect 451794 165134 452414 165218
rect 451794 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 452414 165134
rect 451794 129454 452414 164898
rect 451794 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 452414 129454
rect 451794 129134 452414 129218
rect 451794 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 452414 129134
rect 451794 93454 452414 128898
rect 451794 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 452414 93454
rect 451794 93134 452414 93218
rect 451794 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 452414 93134
rect 451794 57454 452414 92898
rect 451794 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 452414 57454
rect 451794 57134 452414 57218
rect 451794 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 452414 57134
rect 451794 21454 452414 56898
rect 451794 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 452414 21454
rect 451794 21134 452414 21218
rect 451794 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 452414 21134
rect 451794 -1306 452414 20898
rect 451794 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 452414 -1306
rect 451794 -1626 452414 -1542
rect 451794 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 452414 -1626
rect 451794 -1894 452414 -1862
rect 455514 673174 456134 707162
rect 455514 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 456134 673174
rect 455514 672854 456134 672938
rect 455514 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 456134 672854
rect 455514 637174 456134 672618
rect 455514 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 456134 637174
rect 455514 636854 456134 636938
rect 455514 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 456134 636854
rect 455514 601174 456134 636618
rect 455514 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 456134 601174
rect 455514 600854 456134 600938
rect 455514 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 456134 600854
rect 455514 565174 456134 600618
rect 455514 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 456134 565174
rect 455514 564854 456134 564938
rect 455514 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 456134 564854
rect 455514 529174 456134 564618
rect 455514 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 456134 529174
rect 455514 528854 456134 528938
rect 455514 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 456134 528854
rect 455514 493174 456134 528618
rect 455514 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 456134 493174
rect 455514 492854 456134 492938
rect 455514 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 456134 492854
rect 455514 457174 456134 492618
rect 455514 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 456134 457174
rect 455514 456854 456134 456938
rect 455514 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 456134 456854
rect 455514 421174 456134 456618
rect 455514 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 456134 421174
rect 455514 420854 456134 420938
rect 455514 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 456134 420854
rect 455514 385174 456134 420618
rect 455514 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 456134 385174
rect 455514 384854 456134 384938
rect 455514 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 456134 384854
rect 455514 349174 456134 384618
rect 455514 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 456134 349174
rect 455514 348854 456134 348938
rect 455514 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 456134 348854
rect 455514 313174 456134 348618
rect 455514 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 456134 313174
rect 455514 312854 456134 312938
rect 455514 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 456134 312854
rect 455514 277174 456134 312618
rect 455514 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 456134 277174
rect 455514 276854 456134 276938
rect 455514 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 456134 276854
rect 455514 241174 456134 276618
rect 455514 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 456134 241174
rect 455514 240854 456134 240938
rect 455514 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 456134 240854
rect 455514 205174 456134 240618
rect 455514 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 456134 205174
rect 455514 204854 456134 204938
rect 455514 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 456134 204854
rect 455514 169174 456134 204618
rect 455514 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 456134 169174
rect 455514 168854 456134 168938
rect 455514 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 456134 168854
rect 455514 133174 456134 168618
rect 455514 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 456134 133174
rect 455514 132854 456134 132938
rect 455514 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 456134 132854
rect 455514 97174 456134 132618
rect 455514 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 456134 97174
rect 455514 96854 456134 96938
rect 455514 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 456134 96854
rect 455514 61174 456134 96618
rect 455514 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 456134 61174
rect 455514 60854 456134 60938
rect 455514 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 456134 60854
rect 455514 25174 456134 60618
rect 455514 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 456134 25174
rect 455514 24854 456134 24938
rect 455514 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 456134 24854
rect 455514 -3226 456134 24618
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 676894 459854 709082
rect 459234 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 459854 676894
rect 459234 676574 459854 676658
rect 459234 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 459854 676574
rect 459234 640894 459854 676338
rect 459234 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 459854 640894
rect 459234 640574 459854 640658
rect 459234 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 459854 640574
rect 459234 604894 459854 640338
rect 459234 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 459854 604894
rect 459234 604574 459854 604658
rect 459234 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 459854 604574
rect 459234 568894 459854 604338
rect 459234 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 459854 568894
rect 459234 568574 459854 568658
rect 459234 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 459854 568574
rect 459234 532894 459854 568338
rect 459234 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 459854 532894
rect 459234 532574 459854 532658
rect 459234 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 459854 532574
rect 459234 496894 459854 532338
rect 459234 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 459854 496894
rect 459234 496574 459854 496658
rect 459234 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 459854 496574
rect 459234 460894 459854 496338
rect 459234 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 459854 460894
rect 459234 460574 459854 460658
rect 459234 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 459854 460574
rect 459234 424894 459854 460338
rect 459234 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 459854 424894
rect 459234 424574 459854 424658
rect 459234 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 459854 424574
rect 459234 388894 459854 424338
rect 459234 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 459854 388894
rect 459234 388574 459854 388658
rect 459234 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 459854 388574
rect 459234 352894 459854 388338
rect 459234 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 459854 352894
rect 459234 352574 459854 352658
rect 459234 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 459854 352574
rect 459234 316894 459854 352338
rect 459234 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 459854 316894
rect 459234 316574 459854 316658
rect 459234 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 459854 316574
rect 459234 280894 459854 316338
rect 459234 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 459854 280894
rect 459234 280574 459854 280658
rect 459234 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 459854 280574
rect 459234 244894 459854 280338
rect 459234 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 459854 244894
rect 459234 244574 459854 244658
rect 459234 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 459854 244574
rect 459234 208894 459854 244338
rect 459234 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 459854 208894
rect 459234 208574 459854 208658
rect 459234 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 459854 208574
rect 459234 172894 459854 208338
rect 459234 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 459854 172894
rect 459234 172574 459854 172658
rect 459234 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 459854 172574
rect 459234 136894 459854 172338
rect 459234 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 459854 136894
rect 459234 136574 459854 136658
rect 459234 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 459854 136574
rect 459234 100894 459854 136338
rect 459234 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 459854 100894
rect 459234 100574 459854 100658
rect 459234 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 459854 100574
rect 459234 64894 459854 100338
rect 459234 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 459854 64894
rect 459234 64574 459854 64658
rect 459234 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 459854 64574
rect 459234 28894 459854 64338
rect 459234 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 459854 28894
rect 459234 28574 459854 28658
rect 459234 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 459854 28574
rect 459234 -5146 459854 28338
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 462954 680614 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 462954 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 463574 680614
rect 462954 680294 463574 680378
rect 462954 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 463574 680294
rect 462954 644614 463574 680058
rect 462954 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 463574 644614
rect 462954 644294 463574 644378
rect 462954 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 463574 644294
rect 462954 608614 463574 644058
rect 462954 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 463574 608614
rect 462954 608294 463574 608378
rect 462954 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 463574 608294
rect 462954 572614 463574 608058
rect 462954 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 463574 572614
rect 462954 572294 463574 572378
rect 462954 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 463574 572294
rect 462954 536614 463574 572058
rect 462954 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 463574 536614
rect 462954 536294 463574 536378
rect 462954 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 463574 536294
rect 462954 500614 463574 536058
rect 462954 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 463574 500614
rect 462954 500294 463574 500378
rect 462954 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 463574 500294
rect 462954 464614 463574 500058
rect 462954 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 463574 464614
rect 462954 464294 463574 464378
rect 462954 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 463574 464294
rect 462954 428614 463574 464058
rect 462954 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 463574 428614
rect 462954 428294 463574 428378
rect 462954 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 463574 428294
rect 462954 392614 463574 428058
rect 462954 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 463574 392614
rect 462954 392294 463574 392378
rect 462954 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 463574 392294
rect 462954 356614 463574 392058
rect 462954 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 463574 356614
rect 462954 356294 463574 356378
rect 462954 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 463574 356294
rect 462954 320614 463574 356058
rect 462954 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 463574 320614
rect 462954 320294 463574 320378
rect 462954 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 463574 320294
rect 462954 284614 463574 320058
rect 462954 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 463574 284614
rect 462954 284294 463574 284378
rect 462954 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 463574 284294
rect 462954 248614 463574 284058
rect 462954 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 463574 248614
rect 462954 248294 463574 248378
rect 462954 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 463574 248294
rect 462954 212614 463574 248058
rect 462954 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 463574 212614
rect 462954 212294 463574 212378
rect 462954 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 463574 212294
rect 462954 176614 463574 212058
rect 462954 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 463574 176614
rect 462954 176294 463574 176378
rect 462954 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 463574 176294
rect 462954 140614 463574 176058
rect 462954 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 463574 140614
rect 462954 140294 463574 140378
rect 462954 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 463574 140294
rect 462954 104614 463574 140058
rect 462954 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 463574 104614
rect 462954 104294 463574 104378
rect 462954 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 463574 104294
rect 462954 68614 463574 104058
rect 462954 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 463574 68614
rect 462954 68294 463574 68378
rect 462954 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 463574 68294
rect 462954 32614 463574 68058
rect 462954 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 463574 32614
rect 462954 32294 463574 32378
rect 462954 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 463574 32294
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 32058
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 687454 470414 704282
rect 469794 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 470414 687454
rect 469794 687134 470414 687218
rect 469794 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 470414 687134
rect 469794 651454 470414 686898
rect 469794 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 470414 651454
rect 469794 651134 470414 651218
rect 469794 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 470414 651134
rect 469794 615454 470414 650898
rect 469794 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 470414 615454
rect 469794 615134 470414 615218
rect 469794 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 470414 615134
rect 469794 579454 470414 614898
rect 469794 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 470414 579454
rect 469794 579134 470414 579218
rect 469794 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 470414 579134
rect 469794 543454 470414 578898
rect 469794 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 470414 543454
rect 469794 543134 470414 543218
rect 469794 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 470414 543134
rect 469794 507454 470414 542898
rect 469794 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 470414 507454
rect 469794 507134 470414 507218
rect 469794 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 470414 507134
rect 469794 471454 470414 506898
rect 469794 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 470414 471454
rect 469794 471134 470414 471218
rect 469794 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 470414 471134
rect 469794 435454 470414 470898
rect 469794 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 470414 435454
rect 469794 435134 470414 435218
rect 469794 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 470414 435134
rect 469794 399454 470414 434898
rect 469794 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 470414 399454
rect 469794 399134 470414 399218
rect 469794 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 470414 399134
rect 469794 363454 470414 398898
rect 469794 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 470414 363454
rect 469794 363134 470414 363218
rect 469794 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 470414 363134
rect 469794 327454 470414 362898
rect 469794 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 470414 327454
rect 469794 327134 470414 327218
rect 469794 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 470414 327134
rect 469794 291454 470414 326898
rect 469794 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 470414 291454
rect 469794 291134 470414 291218
rect 469794 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 470414 291134
rect 469794 255454 470414 290898
rect 469794 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 470414 255454
rect 469794 255134 470414 255218
rect 469794 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 470414 255134
rect 469794 219454 470414 254898
rect 469794 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 470414 219454
rect 469794 219134 470414 219218
rect 469794 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 470414 219134
rect 469794 183454 470414 218898
rect 469794 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 470414 183454
rect 469794 183134 470414 183218
rect 469794 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 470414 183134
rect 469794 147454 470414 182898
rect 469794 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 470414 147454
rect 469794 147134 470414 147218
rect 469794 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 470414 147134
rect 469794 111454 470414 146898
rect 469794 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 470414 111454
rect 469794 111134 470414 111218
rect 469794 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 470414 111134
rect 469794 75454 470414 110898
rect 469794 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 470414 75454
rect 469794 75134 470414 75218
rect 469794 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 470414 75134
rect 469794 39454 470414 74898
rect 469794 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 470414 39454
rect 469794 39134 470414 39218
rect 469794 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 470414 39134
rect 469794 3454 470414 38898
rect 469794 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 470414 3454
rect 469794 3134 470414 3218
rect 469794 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 470414 3134
rect 469794 -346 470414 2898
rect 469794 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 470414 -346
rect 469794 -666 470414 -582
rect 469794 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 470414 -666
rect 469794 -1894 470414 -902
rect 473514 691174 474134 706202
rect 473514 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 474134 691174
rect 473514 690854 474134 690938
rect 473514 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 474134 690854
rect 473514 655174 474134 690618
rect 473514 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 474134 655174
rect 473514 654854 474134 654938
rect 473514 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 474134 654854
rect 473514 619174 474134 654618
rect 473514 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 474134 619174
rect 473514 618854 474134 618938
rect 473514 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 474134 618854
rect 473514 583174 474134 618618
rect 473514 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 474134 583174
rect 473514 582854 474134 582938
rect 473514 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 474134 582854
rect 473514 547174 474134 582618
rect 473514 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 474134 547174
rect 473514 546854 474134 546938
rect 473514 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 474134 546854
rect 473514 511174 474134 546618
rect 473514 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 474134 511174
rect 473514 510854 474134 510938
rect 473514 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 474134 510854
rect 473514 475174 474134 510618
rect 473514 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 474134 475174
rect 473514 474854 474134 474938
rect 473514 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 474134 474854
rect 473514 439174 474134 474618
rect 473514 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 474134 439174
rect 473514 438854 474134 438938
rect 473514 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 474134 438854
rect 473514 403174 474134 438618
rect 473514 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 474134 403174
rect 473514 402854 474134 402938
rect 473514 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 474134 402854
rect 473514 367174 474134 402618
rect 473514 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 474134 367174
rect 473514 366854 474134 366938
rect 473514 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 474134 366854
rect 473514 331174 474134 366618
rect 473514 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 474134 331174
rect 473514 330854 474134 330938
rect 473514 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 474134 330854
rect 473514 295174 474134 330618
rect 473514 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 474134 295174
rect 473514 294854 474134 294938
rect 473514 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 474134 294854
rect 473514 259174 474134 294618
rect 473514 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 474134 259174
rect 473514 258854 474134 258938
rect 473514 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 474134 258854
rect 473514 223174 474134 258618
rect 473514 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 474134 223174
rect 473514 222854 474134 222938
rect 473514 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 474134 222854
rect 473514 187174 474134 222618
rect 473514 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 474134 187174
rect 473514 186854 474134 186938
rect 473514 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 474134 186854
rect 473514 151174 474134 186618
rect 473514 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 474134 151174
rect 473514 150854 474134 150938
rect 473514 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 474134 150854
rect 473514 115174 474134 150618
rect 473514 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 474134 115174
rect 473514 114854 474134 114938
rect 473514 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 474134 114854
rect 473514 79174 474134 114618
rect 473514 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 474134 79174
rect 473514 78854 474134 78938
rect 473514 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 474134 78854
rect 473514 43174 474134 78618
rect 473514 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 474134 43174
rect 473514 42854 474134 42938
rect 473514 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 474134 42854
rect 473514 7174 474134 42618
rect 473514 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 474134 7174
rect 473514 6854 474134 6938
rect 473514 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 474134 6854
rect 473514 -2266 474134 6618
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 694894 477854 708122
rect 477234 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 477854 694894
rect 477234 694574 477854 694658
rect 477234 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 477854 694574
rect 477234 658894 477854 694338
rect 477234 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 477854 658894
rect 477234 658574 477854 658658
rect 477234 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 477854 658574
rect 477234 622894 477854 658338
rect 477234 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 477854 622894
rect 477234 622574 477854 622658
rect 477234 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 477854 622574
rect 477234 586894 477854 622338
rect 477234 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 477854 586894
rect 477234 586574 477854 586658
rect 477234 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 477854 586574
rect 477234 550894 477854 586338
rect 477234 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 477854 550894
rect 477234 550574 477854 550658
rect 477234 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 477854 550574
rect 477234 514894 477854 550338
rect 477234 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 477854 514894
rect 477234 514574 477854 514658
rect 477234 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 477854 514574
rect 477234 478894 477854 514338
rect 477234 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 477854 478894
rect 477234 478574 477854 478658
rect 477234 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 477854 478574
rect 477234 442894 477854 478338
rect 477234 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 477854 442894
rect 477234 442574 477854 442658
rect 477234 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 477854 442574
rect 477234 406894 477854 442338
rect 477234 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 477854 406894
rect 477234 406574 477854 406658
rect 477234 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 477854 406574
rect 477234 370894 477854 406338
rect 477234 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 477854 370894
rect 477234 370574 477854 370658
rect 477234 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 477854 370574
rect 477234 334894 477854 370338
rect 477234 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 477854 334894
rect 477234 334574 477854 334658
rect 477234 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 477854 334574
rect 477234 298894 477854 334338
rect 477234 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 477854 298894
rect 477234 298574 477854 298658
rect 477234 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 477854 298574
rect 477234 262894 477854 298338
rect 477234 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 477854 262894
rect 477234 262574 477854 262658
rect 477234 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 477854 262574
rect 477234 226894 477854 262338
rect 477234 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 477854 226894
rect 477234 226574 477854 226658
rect 477234 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 477854 226574
rect 477234 190894 477854 226338
rect 477234 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 477854 190894
rect 477234 190574 477854 190658
rect 477234 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 477854 190574
rect 477234 154894 477854 190338
rect 477234 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 477854 154894
rect 477234 154574 477854 154658
rect 477234 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 477854 154574
rect 477234 118894 477854 154338
rect 477234 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 477854 118894
rect 477234 118574 477854 118658
rect 477234 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 477854 118574
rect 477234 82894 477854 118338
rect 477234 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 477854 82894
rect 477234 82574 477854 82658
rect 477234 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 477854 82574
rect 477234 46894 477854 82338
rect 477234 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 477854 46894
rect 477234 46574 477854 46658
rect 477234 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 477854 46574
rect 477234 10894 477854 46338
rect 477234 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 477854 10894
rect 477234 10574 477854 10658
rect 477234 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 477854 10574
rect 477234 -4186 477854 10338
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 480954 698614 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 480954 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 481574 698614
rect 480954 698294 481574 698378
rect 480954 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 481574 698294
rect 480954 662614 481574 698058
rect 480954 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 481574 662614
rect 480954 662294 481574 662378
rect 480954 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 481574 662294
rect 480954 626614 481574 662058
rect 480954 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 481574 626614
rect 480954 626294 481574 626378
rect 480954 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 481574 626294
rect 480954 590614 481574 626058
rect 480954 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 481574 590614
rect 480954 590294 481574 590378
rect 480954 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 481574 590294
rect 480954 554614 481574 590058
rect 480954 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 481574 554614
rect 480954 554294 481574 554378
rect 480954 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 481574 554294
rect 480954 518614 481574 554058
rect 480954 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 481574 518614
rect 480954 518294 481574 518378
rect 480954 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 481574 518294
rect 480954 482614 481574 518058
rect 480954 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 481574 482614
rect 480954 482294 481574 482378
rect 480954 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 481574 482294
rect 480954 446614 481574 482058
rect 480954 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 481574 446614
rect 480954 446294 481574 446378
rect 480954 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 481574 446294
rect 480954 410614 481574 446058
rect 480954 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 481574 410614
rect 480954 410294 481574 410378
rect 480954 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 481574 410294
rect 480954 374614 481574 410058
rect 480954 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 481574 374614
rect 480954 374294 481574 374378
rect 480954 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 481574 374294
rect 480954 338614 481574 374058
rect 480954 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 481574 338614
rect 480954 338294 481574 338378
rect 480954 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 481574 338294
rect 480954 302614 481574 338058
rect 480954 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 481574 302614
rect 480954 302294 481574 302378
rect 480954 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 481574 302294
rect 480954 266614 481574 302058
rect 480954 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 481574 266614
rect 480954 266294 481574 266378
rect 480954 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 481574 266294
rect 480954 230614 481574 266058
rect 480954 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 481574 230614
rect 480954 230294 481574 230378
rect 480954 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 481574 230294
rect 480954 194614 481574 230058
rect 480954 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 481574 194614
rect 480954 194294 481574 194378
rect 480954 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 481574 194294
rect 480954 158614 481574 194058
rect 480954 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 481574 158614
rect 480954 158294 481574 158378
rect 480954 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 481574 158294
rect 480954 122614 481574 158058
rect 480954 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 481574 122614
rect 480954 122294 481574 122378
rect 480954 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 481574 122294
rect 480954 86614 481574 122058
rect 480954 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 481574 86614
rect 480954 86294 481574 86378
rect 480954 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 481574 86294
rect 480954 50614 481574 86058
rect 480954 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 481574 50614
rect 480954 50294 481574 50378
rect 480954 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 481574 50294
rect 480954 14614 481574 50058
rect 480954 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 481574 14614
rect 480954 14294 481574 14378
rect 480954 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 481574 14294
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 14058
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 669454 488414 705242
rect 487794 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 488414 669454
rect 487794 669134 488414 669218
rect 487794 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 488414 669134
rect 487794 633454 488414 668898
rect 487794 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 488414 633454
rect 487794 633134 488414 633218
rect 487794 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 488414 633134
rect 487794 597454 488414 632898
rect 487794 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 488414 597454
rect 487794 597134 488414 597218
rect 487794 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 488414 597134
rect 487794 561454 488414 596898
rect 487794 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 488414 561454
rect 487794 561134 488414 561218
rect 487794 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 488414 561134
rect 487794 525454 488414 560898
rect 487794 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 488414 525454
rect 487794 525134 488414 525218
rect 487794 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 488414 525134
rect 487794 489454 488414 524898
rect 487794 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 488414 489454
rect 487794 489134 488414 489218
rect 487794 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 488414 489134
rect 487794 453454 488414 488898
rect 487794 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 488414 453454
rect 487794 453134 488414 453218
rect 487794 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 488414 453134
rect 487794 417454 488414 452898
rect 487794 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 488414 417454
rect 487794 417134 488414 417218
rect 487794 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 488414 417134
rect 487794 381454 488414 416898
rect 487794 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 488414 381454
rect 487794 381134 488414 381218
rect 487794 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 488414 381134
rect 487794 345454 488414 380898
rect 487794 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 488414 345454
rect 487794 345134 488414 345218
rect 487794 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 488414 345134
rect 487794 309454 488414 344898
rect 487794 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 488414 309454
rect 487794 309134 488414 309218
rect 487794 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 488414 309134
rect 487794 273454 488414 308898
rect 487794 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 488414 273454
rect 487794 273134 488414 273218
rect 487794 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 488414 273134
rect 487794 237454 488414 272898
rect 487794 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 488414 237454
rect 487794 237134 488414 237218
rect 487794 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 488414 237134
rect 487794 201454 488414 236898
rect 487794 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 488414 201454
rect 487794 201134 488414 201218
rect 487794 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 488414 201134
rect 487794 165454 488414 200898
rect 487794 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 488414 165454
rect 487794 165134 488414 165218
rect 487794 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 488414 165134
rect 487794 129454 488414 164898
rect 487794 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 488414 129454
rect 487794 129134 488414 129218
rect 487794 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 488414 129134
rect 487794 93454 488414 128898
rect 487794 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 488414 93454
rect 487794 93134 488414 93218
rect 487794 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 488414 93134
rect 487794 57454 488414 92898
rect 487794 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 488414 57454
rect 487794 57134 488414 57218
rect 487794 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 488414 57134
rect 487794 21454 488414 56898
rect 487794 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 488414 21454
rect 487794 21134 488414 21218
rect 487794 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 488414 21134
rect 487794 -1306 488414 20898
rect 487794 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 488414 -1306
rect 487794 -1626 488414 -1542
rect 487794 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 488414 -1626
rect 487794 -1894 488414 -1862
rect 491514 673174 492134 707162
rect 491514 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 492134 673174
rect 491514 672854 492134 672938
rect 491514 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 492134 672854
rect 491514 637174 492134 672618
rect 491514 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 492134 637174
rect 491514 636854 492134 636938
rect 491514 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 492134 636854
rect 491514 601174 492134 636618
rect 491514 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 492134 601174
rect 491514 600854 492134 600938
rect 491514 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 492134 600854
rect 491514 565174 492134 600618
rect 491514 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 492134 565174
rect 491514 564854 492134 564938
rect 491514 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 492134 564854
rect 491514 529174 492134 564618
rect 491514 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 492134 529174
rect 491514 528854 492134 528938
rect 491514 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 492134 528854
rect 491514 493174 492134 528618
rect 491514 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 492134 493174
rect 491514 492854 492134 492938
rect 491514 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 492134 492854
rect 491514 457174 492134 492618
rect 491514 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 492134 457174
rect 491514 456854 492134 456938
rect 491514 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 492134 456854
rect 491514 421174 492134 456618
rect 491514 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 492134 421174
rect 491514 420854 492134 420938
rect 491514 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 492134 420854
rect 491514 385174 492134 420618
rect 491514 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 492134 385174
rect 491514 384854 492134 384938
rect 491514 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 492134 384854
rect 491514 349174 492134 384618
rect 491514 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 492134 349174
rect 491514 348854 492134 348938
rect 491514 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 492134 348854
rect 491514 313174 492134 348618
rect 491514 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 492134 313174
rect 491514 312854 492134 312938
rect 491514 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 492134 312854
rect 491514 277174 492134 312618
rect 491514 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 492134 277174
rect 491514 276854 492134 276938
rect 491514 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 492134 276854
rect 491514 241174 492134 276618
rect 491514 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 492134 241174
rect 491514 240854 492134 240938
rect 491514 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 492134 240854
rect 491514 205174 492134 240618
rect 491514 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 492134 205174
rect 491514 204854 492134 204938
rect 491514 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 492134 204854
rect 491514 169174 492134 204618
rect 491514 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 492134 169174
rect 491514 168854 492134 168938
rect 491514 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 492134 168854
rect 491514 133174 492134 168618
rect 491514 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 492134 133174
rect 491514 132854 492134 132938
rect 491514 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 492134 132854
rect 491514 97174 492134 132618
rect 491514 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 492134 97174
rect 491514 96854 492134 96938
rect 491514 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 492134 96854
rect 491514 61174 492134 96618
rect 491514 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 492134 61174
rect 491514 60854 492134 60938
rect 491514 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 492134 60854
rect 491514 25174 492134 60618
rect 491514 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 492134 25174
rect 491514 24854 492134 24938
rect 491514 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 492134 24854
rect 491514 -3226 492134 24618
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 676894 495854 709082
rect 495234 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 495854 676894
rect 495234 676574 495854 676658
rect 495234 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 495854 676574
rect 495234 640894 495854 676338
rect 495234 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 495854 640894
rect 495234 640574 495854 640658
rect 495234 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 495854 640574
rect 495234 604894 495854 640338
rect 495234 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 495854 604894
rect 495234 604574 495854 604658
rect 495234 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 495854 604574
rect 495234 568894 495854 604338
rect 495234 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 495854 568894
rect 495234 568574 495854 568658
rect 495234 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 495854 568574
rect 495234 532894 495854 568338
rect 495234 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 495854 532894
rect 495234 532574 495854 532658
rect 495234 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 495854 532574
rect 495234 496894 495854 532338
rect 495234 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 495854 496894
rect 495234 496574 495854 496658
rect 495234 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 495854 496574
rect 495234 460894 495854 496338
rect 495234 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 495854 460894
rect 495234 460574 495854 460658
rect 495234 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 495854 460574
rect 495234 424894 495854 460338
rect 495234 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 495854 424894
rect 495234 424574 495854 424658
rect 495234 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 495854 424574
rect 495234 388894 495854 424338
rect 495234 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 495854 388894
rect 495234 388574 495854 388658
rect 495234 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 495854 388574
rect 495234 352894 495854 388338
rect 495234 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 495854 352894
rect 495234 352574 495854 352658
rect 495234 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 495854 352574
rect 495234 316894 495854 352338
rect 495234 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 495854 316894
rect 495234 316574 495854 316658
rect 495234 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 495854 316574
rect 495234 280894 495854 316338
rect 495234 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 495854 280894
rect 495234 280574 495854 280658
rect 495234 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 495854 280574
rect 495234 244894 495854 280338
rect 495234 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 495854 244894
rect 495234 244574 495854 244658
rect 495234 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 495854 244574
rect 495234 208894 495854 244338
rect 495234 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 495854 208894
rect 495234 208574 495854 208658
rect 495234 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 495854 208574
rect 495234 172894 495854 208338
rect 495234 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 495854 172894
rect 495234 172574 495854 172658
rect 495234 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 495854 172574
rect 495234 136894 495854 172338
rect 495234 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 495854 136894
rect 495234 136574 495854 136658
rect 495234 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 495854 136574
rect 495234 100894 495854 136338
rect 495234 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 495854 100894
rect 495234 100574 495854 100658
rect 495234 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 495854 100574
rect 495234 64894 495854 100338
rect 495234 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 495854 64894
rect 495234 64574 495854 64658
rect 495234 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 495854 64574
rect 495234 28894 495854 64338
rect 495234 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 495854 28894
rect 495234 28574 495854 28658
rect 495234 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 495854 28574
rect 495234 -5146 495854 28338
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 498954 680614 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 498954 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 499574 680614
rect 498954 680294 499574 680378
rect 498954 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 499574 680294
rect 498954 644614 499574 680058
rect 498954 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 499574 644614
rect 498954 644294 499574 644378
rect 498954 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 499574 644294
rect 498954 608614 499574 644058
rect 498954 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 499574 608614
rect 498954 608294 499574 608378
rect 498954 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 499574 608294
rect 498954 572614 499574 608058
rect 498954 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 499574 572614
rect 498954 572294 499574 572378
rect 498954 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 499574 572294
rect 498954 536614 499574 572058
rect 498954 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 499574 536614
rect 498954 536294 499574 536378
rect 498954 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 499574 536294
rect 498954 500614 499574 536058
rect 498954 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 499574 500614
rect 498954 500294 499574 500378
rect 498954 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 499574 500294
rect 498954 464614 499574 500058
rect 498954 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 499574 464614
rect 498954 464294 499574 464378
rect 498954 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 499574 464294
rect 498954 428614 499574 464058
rect 498954 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 499574 428614
rect 498954 428294 499574 428378
rect 498954 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 499574 428294
rect 498954 392614 499574 428058
rect 498954 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 499574 392614
rect 498954 392294 499574 392378
rect 498954 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 499574 392294
rect 498954 356614 499574 392058
rect 498954 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 499574 356614
rect 498954 356294 499574 356378
rect 498954 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 499574 356294
rect 498954 320614 499574 356058
rect 498954 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 499574 320614
rect 498954 320294 499574 320378
rect 498954 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 499574 320294
rect 498954 284614 499574 320058
rect 498954 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 499574 284614
rect 498954 284294 499574 284378
rect 498954 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 499574 284294
rect 498954 248614 499574 284058
rect 498954 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 499574 248614
rect 498954 248294 499574 248378
rect 498954 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 499574 248294
rect 498954 212614 499574 248058
rect 498954 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 499574 212614
rect 498954 212294 499574 212378
rect 498954 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 499574 212294
rect 498954 176614 499574 212058
rect 498954 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 499574 176614
rect 498954 176294 499574 176378
rect 498954 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 499574 176294
rect 498954 140614 499574 176058
rect 498954 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 499574 140614
rect 498954 140294 499574 140378
rect 498954 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 499574 140294
rect 498954 104614 499574 140058
rect 498954 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 499574 104614
rect 498954 104294 499574 104378
rect 498954 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 499574 104294
rect 498954 68614 499574 104058
rect 498954 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 499574 68614
rect 498954 68294 499574 68378
rect 498954 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 499574 68294
rect 498954 32614 499574 68058
rect 498954 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 499574 32614
rect 498954 32294 499574 32378
rect 498954 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 499574 32294
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 32058
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 687454 506414 704282
rect 505794 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 506414 687454
rect 505794 687134 506414 687218
rect 505794 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 506414 687134
rect 505794 651454 506414 686898
rect 505794 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 506414 651454
rect 505794 651134 506414 651218
rect 505794 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 506414 651134
rect 505794 615454 506414 650898
rect 505794 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 506414 615454
rect 505794 615134 506414 615218
rect 505794 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 506414 615134
rect 505794 579454 506414 614898
rect 505794 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 506414 579454
rect 505794 579134 506414 579218
rect 505794 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 506414 579134
rect 505794 543454 506414 578898
rect 505794 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 506414 543454
rect 505794 543134 506414 543218
rect 505794 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 506414 543134
rect 505794 507454 506414 542898
rect 505794 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 506414 507454
rect 505794 507134 506414 507218
rect 505794 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 506414 507134
rect 505794 471454 506414 506898
rect 505794 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 506414 471454
rect 505794 471134 506414 471218
rect 505794 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 506414 471134
rect 505794 435454 506414 470898
rect 505794 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 506414 435454
rect 505794 435134 506414 435218
rect 505794 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 506414 435134
rect 505794 399454 506414 434898
rect 505794 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 506414 399454
rect 505794 399134 506414 399218
rect 505794 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 506414 399134
rect 505794 363454 506414 398898
rect 505794 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 506414 363454
rect 505794 363134 506414 363218
rect 505794 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 506414 363134
rect 505794 327454 506414 362898
rect 505794 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 506414 327454
rect 505794 327134 506414 327218
rect 505794 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 506414 327134
rect 505794 291454 506414 326898
rect 505794 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 506414 291454
rect 505794 291134 506414 291218
rect 505794 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 506414 291134
rect 505794 255454 506414 290898
rect 505794 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 506414 255454
rect 505794 255134 506414 255218
rect 505794 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 506414 255134
rect 505794 219454 506414 254898
rect 505794 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 506414 219454
rect 505794 219134 506414 219218
rect 505794 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 506414 219134
rect 505794 183454 506414 218898
rect 505794 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 506414 183454
rect 505794 183134 506414 183218
rect 505794 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 506414 183134
rect 505794 147454 506414 182898
rect 505794 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 506414 147454
rect 505794 147134 506414 147218
rect 505794 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 506414 147134
rect 505794 111454 506414 146898
rect 505794 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 506414 111454
rect 505794 111134 506414 111218
rect 505794 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 506414 111134
rect 505794 75454 506414 110898
rect 505794 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 506414 75454
rect 505794 75134 506414 75218
rect 505794 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 506414 75134
rect 505794 39454 506414 74898
rect 505794 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 506414 39454
rect 505794 39134 506414 39218
rect 505794 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 506414 39134
rect 505794 3454 506414 38898
rect 505794 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 506414 3454
rect 505794 3134 506414 3218
rect 505794 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 506414 3134
rect 505794 -346 506414 2898
rect 505794 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 506414 -346
rect 505794 -666 506414 -582
rect 505794 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 506414 -666
rect 505794 -1894 506414 -902
rect 509514 691174 510134 706202
rect 509514 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 510134 691174
rect 509514 690854 510134 690938
rect 509514 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 510134 690854
rect 509514 655174 510134 690618
rect 509514 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 510134 655174
rect 509514 654854 510134 654938
rect 509514 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 510134 654854
rect 509514 619174 510134 654618
rect 509514 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 510134 619174
rect 509514 618854 510134 618938
rect 509514 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 510134 618854
rect 509514 583174 510134 618618
rect 509514 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 510134 583174
rect 509514 582854 510134 582938
rect 509514 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 510134 582854
rect 509514 547174 510134 582618
rect 509514 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 510134 547174
rect 509514 546854 510134 546938
rect 509514 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 510134 546854
rect 509514 511174 510134 546618
rect 509514 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 510134 511174
rect 509514 510854 510134 510938
rect 509514 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 510134 510854
rect 509514 475174 510134 510618
rect 509514 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 510134 475174
rect 509514 474854 510134 474938
rect 509514 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 510134 474854
rect 509514 439174 510134 474618
rect 509514 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 510134 439174
rect 509514 438854 510134 438938
rect 509514 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 510134 438854
rect 509514 403174 510134 438618
rect 509514 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 510134 403174
rect 509514 402854 510134 402938
rect 509514 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 510134 402854
rect 509514 367174 510134 402618
rect 509514 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 510134 367174
rect 509514 366854 510134 366938
rect 509514 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 510134 366854
rect 509514 331174 510134 366618
rect 509514 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 510134 331174
rect 509514 330854 510134 330938
rect 509514 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 510134 330854
rect 509514 295174 510134 330618
rect 509514 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 510134 295174
rect 509514 294854 510134 294938
rect 509514 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 510134 294854
rect 509514 259174 510134 294618
rect 509514 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 510134 259174
rect 509514 258854 510134 258938
rect 509514 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 510134 258854
rect 509514 223174 510134 258618
rect 509514 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 510134 223174
rect 509514 222854 510134 222938
rect 509514 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 510134 222854
rect 509514 187174 510134 222618
rect 509514 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 510134 187174
rect 509514 186854 510134 186938
rect 509514 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 510134 186854
rect 509514 151174 510134 186618
rect 509514 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 510134 151174
rect 509514 150854 510134 150938
rect 509514 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 510134 150854
rect 509514 115174 510134 150618
rect 509514 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 510134 115174
rect 509514 114854 510134 114938
rect 509514 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 510134 114854
rect 509514 79174 510134 114618
rect 509514 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 510134 79174
rect 509514 78854 510134 78938
rect 509514 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 510134 78854
rect 509514 43174 510134 78618
rect 509514 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 510134 43174
rect 509514 42854 510134 42938
rect 509514 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 510134 42854
rect 509514 7174 510134 42618
rect 509514 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 510134 7174
rect 509514 6854 510134 6938
rect 509514 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 510134 6854
rect 509514 -2266 510134 6618
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 694894 513854 708122
rect 513234 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 513854 694894
rect 513234 694574 513854 694658
rect 513234 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 513854 694574
rect 513234 658894 513854 694338
rect 513234 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 513854 658894
rect 513234 658574 513854 658658
rect 513234 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 513854 658574
rect 513234 622894 513854 658338
rect 513234 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 513854 622894
rect 513234 622574 513854 622658
rect 513234 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 513854 622574
rect 513234 586894 513854 622338
rect 513234 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 513854 586894
rect 513234 586574 513854 586658
rect 513234 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 513854 586574
rect 513234 550894 513854 586338
rect 513234 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 513854 550894
rect 513234 550574 513854 550658
rect 513234 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 513854 550574
rect 513234 514894 513854 550338
rect 513234 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 513854 514894
rect 513234 514574 513854 514658
rect 513234 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 513854 514574
rect 513234 478894 513854 514338
rect 513234 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 513854 478894
rect 513234 478574 513854 478658
rect 513234 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 513854 478574
rect 513234 442894 513854 478338
rect 513234 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 513854 442894
rect 513234 442574 513854 442658
rect 513234 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 513854 442574
rect 513234 406894 513854 442338
rect 513234 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 513854 406894
rect 513234 406574 513854 406658
rect 513234 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 513854 406574
rect 513234 370894 513854 406338
rect 513234 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 513854 370894
rect 513234 370574 513854 370658
rect 513234 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 513854 370574
rect 513234 334894 513854 370338
rect 513234 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 513854 334894
rect 513234 334574 513854 334658
rect 513234 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 513854 334574
rect 513234 298894 513854 334338
rect 513234 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 513854 298894
rect 513234 298574 513854 298658
rect 513234 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 513854 298574
rect 513234 262894 513854 298338
rect 513234 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 513854 262894
rect 513234 262574 513854 262658
rect 513234 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 513854 262574
rect 513234 226894 513854 262338
rect 513234 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 513854 226894
rect 513234 226574 513854 226658
rect 513234 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 513854 226574
rect 513234 190894 513854 226338
rect 513234 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 513854 190894
rect 513234 190574 513854 190658
rect 513234 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 513854 190574
rect 513234 154894 513854 190338
rect 513234 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 513854 154894
rect 513234 154574 513854 154658
rect 513234 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 513854 154574
rect 513234 118894 513854 154338
rect 513234 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 513854 118894
rect 513234 118574 513854 118658
rect 513234 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 513854 118574
rect 513234 82894 513854 118338
rect 513234 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 513854 82894
rect 513234 82574 513854 82658
rect 513234 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 513854 82574
rect 513234 46894 513854 82338
rect 513234 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 513854 46894
rect 513234 46574 513854 46658
rect 513234 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 513854 46574
rect 513234 10894 513854 46338
rect 513234 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 513854 10894
rect 513234 10574 513854 10658
rect 513234 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 513854 10574
rect 513234 -4186 513854 10338
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 516954 698614 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 516954 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 517574 698614
rect 516954 698294 517574 698378
rect 516954 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 517574 698294
rect 516954 662614 517574 698058
rect 516954 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 517574 662614
rect 516954 662294 517574 662378
rect 516954 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 517574 662294
rect 516954 626614 517574 662058
rect 516954 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 517574 626614
rect 516954 626294 517574 626378
rect 516954 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 517574 626294
rect 516954 590614 517574 626058
rect 516954 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 517574 590614
rect 516954 590294 517574 590378
rect 516954 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 517574 590294
rect 516954 554614 517574 590058
rect 516954 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 517574 554614
rect 516954 554294 517574 554378
rect 516954 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 517574 554294
rect 516954 518614 517574 554058
rect 516954 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 517574 518614
rect 516954 518294 517574 518378
rect 516954 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 517574 518294
rect 516954 482614 517574 518058
rect 516954 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 517574 482614
rect 516954 482294 517574 482378
rect 516954 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 517574 482294
rect 516954 446614 517574 482058
rect 516954 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 517574 446614
rect 516954 446294 517574 446378
rect 516954 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 517574 446294
rect 516954 410614 517574 446058
rect 516954 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 517574 410614
rect 516954 410294 517574 410378
rect 516954 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 517574 410294
rect 516954 374614 517574 410058
rect 516954 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 517574 374614
rect 516954 374294 517574 374378
rect 516954 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 517574 374294
rect 516954 338614 517574 374058
rect 516954 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 517574 338614
rect 516954 338294 517574 338378
rect 516954 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 517574 338294
rect 516954 302614 517574 338058
rect 516954 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 517574 302614
rect 516954 302294 517574 302378
rect 516954 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 517574 302294
rect 516954 266614 517574 302058
rect 516954 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 517574 266614
rect 516954 266294 517574 266378
rect 516954 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 517574 266294
rect 516954 230614 517574 266058
rect 516954 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 517574 230614
rect 516954 230294 517574 230378
rect 516954 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 517574 230294
rect 516954 194614 517574 230058
rect 516954 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 517574 194614
rect 516954 194294 517574 194378
rect 516954 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 517574 194294
rect 516954 158614 517574 194058
rect 516954 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 517574 158614
rect 516954 158294 517574 158378
rect 516954 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 517574 158294
rect 516954 122614 517574 158058
rect 516954 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 517574 122614
rect 516954 122294 517574 122378
rect 516954 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 517574 122294
rect 516954 86614 517574 122058
rect 516954 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 517574 86614
rect 516954 86294 517574 86378
rect 516954 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 517574 86294
rect 516954 50614 517574 86058
rect 516954 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 517574 50614
rect 516954 50294 517574 50378
rect 516954 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 517574 50294
rect 516954 14614 517574 50058
rect 516954 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 517574 14614
rect 516954 14294 517574 14378
rect 516954 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 517574 14294
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 14058
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 669454 524414 705242
rect 523794 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 524414 669454
rect 523794 669134 524414 669218
rect 523794 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 524414 669134
rect 523794 633454 524414 668898
rect 523794 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 524414 633454
rect 523794 633134 524414 633218
rect 523794 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 524414 633134
rect 523794 597454 524414 632898
rect 523794 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 524414 597454
rect 523794 597134 524414 597218
rect 523794 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 524414 597134
rect 523794 561454 524414 596898
rect 523794 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 524414 561454
rect 523794 561134 524414 561218
rect 523794 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 524414 561134
rect 523794 525454 524414 560898
rect 523794 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 524414 525454
rect 523794 525134 524414 525218
rect 523794 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 524414 525134
rect 523794 489454 524414 524898
rect 523794 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 524414 489454
rect 523794 489134 524414 489218
rect 523794 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 524414 489134
rect 523794 453454 524414 488898
rect 523794 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 524414 453454
rect 523794 453134 524414 453218
rect 523794 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 524414 453134
rect 523794 417454 524414 452898
rect 523794 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 524414 417454
rect 523794 417134 524414 417218
rect 523794 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 524414 417134
rect 523794 381454 524414 416898
rect 523794 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 524414 381454
rect 523794 381134 524414 381218
rect 523794 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 524414 381134
rect 523794 345454 524414 380898
rect 523794 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 524414 345454
rect 523794 345134 524414 345218
rect 523794 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 524414 345134
rect 523794 309454 524414 344898
rect 523794 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 524414 309454
rect 523794 309134 524414 309218
rect 523794 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 524414 309134
rect 523794 273454 524414 308898
rect 523794 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 524414 273454
rect 523794 273134 524414 273218
rect 523794 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 524414 273134
rect 523794 237454 524414 272898
rect 523794 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 524414 237454
rect 523794 237134 524414 237218
rect 523794 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 524414 237134
rect 523794 201454 524414 236898
rect 523794 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 524414 201454
rect 523794 201134 524414 201218
rect 523794 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 524414 201134
rect 523794 165454 524414 200898
rect 523794 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 524414 165454
rect 523794 165134 524414 165218
rect 523794 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 524414 165134
rect 523794 129454 524414 164898
rect 523794 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 524414 129454
rect 523794 129134 524414 129218
rect 523794 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 524414 129134
rect 523794 93454 524414 128898
rect 523794 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 524414 93454
rect 523794 93134 524414 93218
rect 523794 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 524414 93134
rect 523794 57454 524414 92898
rect 523794 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 524414 57454
rect 523794 57134 524414 57218
rect 523794 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 524414 57134
rect 523794 21454 524414 56898
rect 523794 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 524414 21454
rect 523794 21134 524414 21218
rect 523794 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 524414 21134
rect 523794 -1306 524414 20898
rect 523794 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 524414 -1306
rect 523794 -1626 524414 -1542
rect 523794 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 524414 -1626
rect 523794 -1894 524414 -1862
rect 527514 673174 528134 707162
rect 527514 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 528134 673174
rect 527514 672854 528134 672938
rect 527514 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 528134 672854
rect 527514 637174 528134 672618
rect 527514 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 528134 637174
rect 527514 636854 528134 636938
rect 527514 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 528134 636854
rect 527514 601174 528134 636618
rect 527514 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 528134 601174
rect 527514 600854 528134 600938
rect 527514 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 528134 600854
rect 527514 565174 528134 600618
rect 527514 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 528134 565174
rect 527514 564854 528134 564938
rect 527514 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 528134 564854
rect 527514 529174 528134 564618
rect 527514 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 528134 529174
rect 527514 528854 528134 528938
rect 527514 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 528134 528854
rect 527514 493174 528134 528618
rect 527514 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 528134 493174
rect 527514 492854 528134 492938
rect 527514 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 528134 492854
rect 527514 457174 528134 492618
rect 527514 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 528134 457174
rect 527514 456854 528134 456938
rect 527514 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 528134 456854
rect 527514 421174 528134 456618
rect 527514 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 528134 421174
rect 527514 420854 528134 420938
rect 527514 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 528134 420854
rect 527514 385174 528134 420618
rect 527514 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 528134 385174
rect 527514 384854 528134 384938
rect 527514 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 528134 384854
rect 527514 349174 528134 384618
rect 527514 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 528134 349174
rect 527514 348854 528134 348938
rect 527514 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 528134 348854
rect 527514 313174 528134 348618
rect 527514 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 528134 313174
rect 527514 312854 528134 312938
rect 527514 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 528134 312854
rect 527514 277174 528134 312618
rect 527514 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 528134 277174
rect 527514 276854 528134 276938
rect 527514 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 528134 276854
rect 527514 241174 528134 276618
rect 527514 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 528134 241174
rect 527514 240854 528134 240938
rect 527514 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 528134 240854
rect 527514 205174 528134 240618
rect 527514 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 528134 205174
rect 527514 204854 528134 204938
rect 527514 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 528134 204854
rect 527514 169174 528134 204618
rect 527514 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 528134 169174
rect 527514 168854 528134 168938
rect 527514 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 528134 168854
rect 527514 133174 528134 168618
rect 527514 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 528134 133174
rect 527514 132854 528134 132938
rect 527514 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 528134 132854
rect 527514 97174 528134 132618
rect 527514 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 528134 97174
rect 527514 96854 528134 96938
rect 527514 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 528134 96854
rect 527514 61174 528134 96618
rect 527514 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 528134 61174
rect 527514 60854 528134 60938
rect 527514 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 528134 60854
rect 527514 25174 528134 60618
rect 527514 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 528134 25174
rect 527514 24854 528134 24938
rect 527514 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 528134 24854
rect 527514 -3226 528134 24618
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 676894 531854 709082
rect 531234 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 531854 676894
rect 531234 676574 531854 676658
rect 531234 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 531854 676574
rect 531234 640894 531854 676338
rect 531234 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 531854 640894
rect 531234 640574 531854 640658
rect 531234 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 531854 640574
rect 531234 604894 531854 640338
rect 531234 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 531854 604894
rect 531234 604574 531854 604658
rect 531234 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 531854 604574
rect 531234 568894 531854 604338
rect 531234 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 531854 568894
rect 531234 568574 531854 568658
rect 531234 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 531854 568574
rect 531234 532894 531854 568338
rect 531234 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 531854 532894
rect 531234 532574 531854 532658
rect 531234 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 531854 532574
rect 531234 496894 531854 532338
rect 531234 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 531854 496894
rect 531234 496574 531854 496658
rect 531234 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 531854 496574
rect 531234 460894 531854 496338
rect 531234 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 531854 460894
rect 531234 460574 531854 460658
rect 531234 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 531854 460574
rect 531234 424894 531854 460338
rect 531234 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 531854 424894
rect 531234 424574 531854 424658
rect 531234 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 531854 424574
rect 531234 388894 531854 424338
rect 531234 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 531854 388894
rect 531234 388574 531854 388658
rect 531234 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 531854 388574
rect 531234 352894 531854 388338
rect 531234 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 531854 352894
rect 531234 352574 531854 352658
rect 531234 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 531854 352574
rect 531234 316894 531854 352338
rect 531234 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 531854 316894
rect 531234 316574 531854 316658
rect 531234 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 531854 316574
rect 531234 280894 531854 316338
rect 531234 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 531854 280894
rect 531234 280574 531854 280658
rect 531234 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 531854 280574
rect 531234 244894 531854 280338
rect 531234 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 531854 244894
rect 531234 244574 531854 244658
rect 531234 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 531854 244574
rect 531234 208894 531854 244338
rect 531234 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 531854 208894
rect 531234 208574 531854 208658
rect 531234 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 531854 208574
rect 531234 172894 531854 208338
rect 531234 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 531854 172894
rect 531234 172574 531854 172658
rect 531234 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 531854 172574
rect 531234 136894 531854 172338
rect 531234 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 531854 136894
rect 531234 136574 531854 136658
rect 531234 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 531854 136574
rect 531234 100894 531854 136338
rect 531234 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 531854 100894
rect 531234 100574 531854 100658
rect 531234 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 531854 100574
rect 531234 64894 531854 100338
rect 531234 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 531854 64894
rect 531234 64574 531854 64658
rect 531234 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 531854 64574
rect 531234 28894 531854 64338
rect 531234 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 531854 28894
rect 531234 28574 531854 28658
rect 531234 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 531854 28574
rect 531234 -5146 531854 28338
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 534954 680614 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 534954 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 535574 680614
rect 534954 680294 535574 680378
rect 534954 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 535574 680294
rect 534954 644614 535574 680058
rect 534954 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 535574 644614
rect 534954 644294 535574 644378
rect 534954 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 535574 644294
rect 534954 608614 535574 644058
rect 534954 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 535574 608614
rect 534954 608294 535574 608378
rect 534954 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 535574 608294
rect 534954 572614 535574 608058
rect 534954 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 535574 572614
rect 534954 572294 535574 572378
rect 534954 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 535574 572294
rect 534954 536614 535574 572058
rect 534954 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 535574 536614
rect 534954 536294 535574 536378
rect 534954 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 535574 536294
rect 534954 500614 535574 536058
rect 534954 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 535574 500614
rect 534954 500294 535574 500378
rect 534954 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 535574 500294
rect 534954 464614 535574 500058
rect 534954 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 535574 464614
rect 534954 464294 535574 464378
rect 534954 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 535574 464294
rect 534954 428614 535574 464058
rect 534954 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 535574 428614
rect 534954 428294 535574 428378
rect 534954 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 535574 428294
rect 534954 392614 535574 428058
rect 534954 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 535574 392614
rect 534954 392294 535574 392378
rect 534954 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 535574 392294
rect 534954 356614 535574 392058
rect 534954 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 535574 356614
rect 534954 356294 535574 356378
rect 534954 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 535574 356294
rect 534954 320614 535574 356058
rect 534954 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 535574 320614
rect 534954 320294 535574 320378
rect 534954 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 535574 320294
rect 534954 284614 535574 320058
rect 534954 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 535574 284614
rect 534954 284294 535574 284378
rect 534954 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 535574 284294
rect 534954 248614 535574 284058
rect 534954 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 535574 248614
rect 534954 248294 535574 248378
rect 534954 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 535574 248294
rect 534954 212614 535574 248058
rect 534954 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 535574 212614
rect 534954 212294 535574 212378
rect 534954 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 535574 212294
rect 534954 176614 535574 212058
rect 534954 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 535574 176614
rect 534954 176294 535574 176378
rect 534954 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 535574 176294
rect 534954 140614 535574 176058
rect 534954 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 535574 140614
rect 534954 140294 535574 140378
rect 534954 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 535574 140294
rect 534954 104614 535574 140058
rect 534954 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 535574 104614
rect 534954 104294 535574 104378
rect 534954 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 535574 104294
rect 534954 68614 535574 104058
rect 534954 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 535574 68614
rect 534954 68294 535574 68378
rect 534954 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 535574 68294
rect 534954 32614 535574 68058
rect 534954 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 535574 32614
rect 534954 32294 535574 32378
rect 534954 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 535574 32294
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 32058
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 687454 542414 704282
rect 541794 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 542414 687454
rect 541794 687134 542414 687218
rect 541794 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 542414 687134
rect 541794 651454 542414 686898
rect 541794 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 542414 651454
rect 541794 651134 542414 651218
rect 541794 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 542414 651134
rect 541794 615454 542414 650898
rect 541794 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 542414 615454
rect 541794 615134 542414 615218
rect 541794 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 542414 615134
rect 541794 579454 542414 614898
rect 541794 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 542414 579454
rect 541794 579134 542414 579218
rect 541794 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 542414 579134
rect 541794 543454 542414 578898
rect 541794 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 542414 543454
rect 541794 543134 542414 543218
rect 541794 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 542414 543134
rect 541794 507454 542414 542898
rect 541794 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 542414 507454
rect 541794 507134 542414 507218
rect 541794 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 542414 507134
rect 541794 471454 542414 506898
rect 541794 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 542414 471454
rect 541794 471134 542414 471218
rect 541794 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 542414 471134
rect 541794 435454 542414 470898
rect 541794 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 542414 435454
rect 541794 435134 542414 435218
rect 541794 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 542414 435134
rect 541794 399454 542414 434898
rect 541794 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 542414 399454
rect 541794 399134 542414 399218
rect 541794 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 542414 399134
rect 541794 363454 542414 398898
rect 541794 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 542414 363454
rect 541794 363134 542414 363218
rect 541794 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 542414 363134
rect 541794 327454 542414 362898
rect 541794 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 542414 327454
rect 541794 327134 542414 327218
rect 541794 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 542414 327134
rect 541794 291454 542414 326898
rect 541794 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 542414 291454
rect 541794 291134 542414 291218
rect 541794 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 542414 291134
rect 541794 255454 542414 290898
rect 541794 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 542414 255454
rect 541794 255134 542414 255218
rect 541794 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 542414 255134
rect 541794 219454 542414 254898
rect 541794 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 542414 219454
rect 541794 219134 542414 219218
rect 541794 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 542414 219134
rect 541794 183454 542414 218898
rect 541794 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 542414 183454
rect 541794 183134 542414 183218
rect 541794 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 542414 183134
rect 541794 147454 542414 182898
rect 541794 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 542414 147454
rect 541794 147134 542414 147218
rect 541794 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 542414 147134
rect 541794 111454 542414 146898
rect 541794 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 542414 111454
rect 541794 111134 542414 111218
rect 541794 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 542414 111134
rect 541794 75454 542414 110898
rect 541794 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 542414 75454
rect 541794 75134 542414 75218
rect 541794 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 542414 75134
rect 541794 39454 542414 74898
rect 541794 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 542414 39454
rect 541794 39134 542414 39218
rect 541794 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 542414 39134
rect 541794 3454 542414 38898
rect 541794 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 542414 3454
rect 541794 3134 542414 3218
rect 541794 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 542414 3134
rect 541794 -346 542414 2898
rect 541794 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 542414 -346
rect 541794 -666 542414 -582
rect 541794 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 542414 -666
rect 541794 -1894 542414 -902
rect 545514 691174 546134 706202
rect 545514 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 546134 691174
rect 545514 690854 546134 690938
rect 545514 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 546134 690854
rect 545514 655174 546134 690618
rect 545514 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 546134 655174
rect 545514 654854 546134 654938
rect 545514 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 546134 654854
rect 545514 619174 546134 654618
rect 545514 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 546134 619174
rect 545514 618854 546134 618938
rect 545514 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 546134 618854
rect 545514 583174 546134 618618
rect 545514 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 546134 583174
rect 545514 582854 546134 582938
rect 545514 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 546134 582854
rect 545514 547174 546134 582618
rect 545514 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 546134 547174
rect 545514 546854 546134 546938
rect 545514 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 546134 546854
rect 545514 511174 546134 546618
rect 545514 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 546134 511174
rect 545514 510854 546134 510938
rect 545514 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 546134 510854
rect 545514 475174 546134 510618
rect 545514 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 546134 475174
rect 545514 474854 546134 474938
rect 545514 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 546134 474854
rect 545514 439174 546134 474618
rect 545514 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 546134 439174
rect 545514 438854 546134 438938
rect 545514 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 546134 438854
rect 545514 403174 546134 438618
rect 545514 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 546134 403174
rect 545514 402854 546134 402938
rect 545514 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 546134 402854
rect 545514 367174 546134 402618
rect 545514 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 546134 367174
rect 545514 366854 546134 366938
rect 545514 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 546134 366854
rect 545514 331174 546134 366618
rect 545514 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 546134 331174
rect 545514 330854 546134 330938
rect 545514 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 546134 330854
rect 545514 295174 546134 330618
rect 545514 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 546134 295174
rect 545514 294854 546134 294938
rect 545514 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 546134 294854
rect 545514 259174 546134 294618
rect 545514 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 546134 259174
rect 545514 258854 546134 258938
rect 545514 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 546134 258854
rect 545514 223174 546134 258618
rect 545514 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 546134 223174
rect 545514 222854 546134 222938
rect 545514 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 546134 222854
rect 545514 187174 546134 222618
rect 545514 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 546134 187174
rect 545514 186854 546134 186938
rect 545514 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 546134 186854
rect 545514 151174 546134 186618
rect 545514 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 546134 151174
rect 545514 150854 546134 150938
rect 545514 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 546134 150854
rect 545514 115174 546134 150618
rect 545514 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 546134 115174
rect 545514 114854 546134 114938
rect 545514 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 546134 114854
rect 545514 79174 546134 114618
rect 545514 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 546134 79174
rect 545514 78854 546134 78938
rect 545514 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 546134 78854
rect 545514 43174 546134 78618
rect 545514 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 546134 43174
rect 545514 42854 546134 42938
rect 545514 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 546134 42854
rect 545514 7174 546134 42618
rect 545514 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 546134 7174
rect 545514 6854 546134 6938
rect 545514 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 546134 6854
rect 545514 -2266 546134 6618
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 694894 549854 708122
rect 549234 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 549854 694894
rect 549234 694574 549854 694658
rect 549234 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 549854 694574
rect 549234 658894 549854 694338
rect 549234 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 549854 658894
rect 549234 658574 549854 658658
rect 549234 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 549854 658574
rect 549234 622894 549854 658338
rect 549234 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 549854 622894
rect 549234 622574 549854 622658
rect 549234 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 549854 622574
rect 549234 586894 549854 622338
rect 549234 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 549854 586894
rect 549234 586574 549854 586658
rect 549234 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 549854 586574
rect 549234 550894 549854 586338
rect 549234 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 549854 550894
rect 549234 550574 549854 550658
rect 549234 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 549854 550574
rect 549234 514894 549854 550338
rect 549234 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 549854 514894
rect 549234 514574 549854 514658
rect 549234 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 549854 514574
rect 549234 478894 549854 514338
rect 549234 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 549854 478894
rect 549234 478574 549854 478658
rect 549234 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 549854 478574
rect 549234 442894 549854 478338
rect 549234 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 549854 442894
rect 549234 442574 549854 442658
rect 549234 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 549854 442574
rect 549234 406894 549854 442338
rect 549234 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 549854 406894
rect 549234 406574 549854 406658
rect 549234 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 549854 406574
rect 549234 370894 549854 406338
rect 549234 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 549854 370894
rect 549234 370574 549854 370658
rect 549234 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 549854 370574
rect 549234 334894 549854 370338
rect 549234 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 549854 334894
rect 549234 334574 549854 334658
rect 549234 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 549854 334574
rect 549234 298894 549854 334338
rect 549234 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 549854 298894
rect 549234 298574 549854 298658
rect 549234 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 549854 298574
rect 549234 262894 549854 298338
rect 549234 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 549854 262894
rect 549234 262574 549854 262658
rect 549234 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 549854 262574
rect 549234 226894 549854 262338
rect 549234 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 549854 226894
rect 549234 226574 549854 226658
rect 549234 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 549854 226574
rect 549234 190894 549854 226338
rect 549234 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 549854 190894
rect 549234 190574 549854 190658
rect 549234 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 549854 190574
rect 549234 154894 549854 190338
rect 549234 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 549854 154894
rect 549234 154574 549854 154658
rect 549234 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 549854 154574
rect 549234 118894 549854 154338
rect 549234 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 549854 118894
rect 549234 118574 549854 118658
rect 549234 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 549854 118574
rect 549234 82894 549854 118338
rect 549234 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 549854 82894
rect 549234 82574 549854 82658
rect 549234 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 549854 82574
rect 549234 46894 549854 82338
rect 549234 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 549854 46894
rect 549234 46574 549854 46658
rect 549234 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 549854 46574
rect 549234 10894 549854 46338
rect 549234 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 549854 10894
rect 549234 10574 549854 10658
rect 549234 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 549854 10574
rect 549234 -4186 549854 10338
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 552954 698614 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 552954 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 553574 698614
rect 552954 698294 553574 698378
rect 552954 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 553574 698294
rect 552954 662614 553574 698058
rect 552954 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 553574 662614
rect 552954 662294 553574 662378
rect 552954 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 553574 662294
rect 552954 626614 553574 662058
rect 552954 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 553574 626614
rect 552954 626294 553574 626378
rect 552954 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 553574 626294
rect 552954 590614 553574 626058
rect 552954 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 553574 590614
rect 552954 590294 553574 590378
rect 552954 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 553574 590294
rect 552954 554614 553574 590058
rect 552954 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 553574 554614
rect 552954 554294 553574 554378
rect 552954 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 553574 554294
rect 552954 518614 553574 554058
rect 552954 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 553574 518614
rect 552954 518294 553574 518378
rect 552954 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 553574 518294
rect 552954 482614 553574 518058
rect 552954 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 553574 482614
rect 552954 482294 553574 482378
rect 552954 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 553574 482294
rect 552954 446614 553574 482058
rect 552954 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 553574 446614
rect 552954 446294 553574 446378
rect 552954 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 553574 446294
rect 552954 410614 553574 446058
rect 552954 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 553574 410614
rect 552954 410294 553574 410378
rect 552954 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 553574 410294
rect 552954 374614 553574 410058
rect 552954 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 553574 374614
rect 552954 374294 553574 374378
rect 552954 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 553574 374294
rect 552954 338614 553574 374058
rect 552954 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 553574 338614
rect 552954 338294 553574 338378
rect 552954 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 553574 338294
rect 552954 302614 553574 338058
rect 552954 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 553574 302614
rect 552954 302294 553574 302378
rect 552954 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 553574 302294
rect 552954 266614 553574 302058
rect 552954 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 553574 266614
rect 552954 266294 553574 266378
rect 552954 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 553574 266294
rect 552954 230614 553574 266058
rect 552954 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 553574 230614
rect 552954 230294 553574 230378
rect 552954 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 553574 230294
rect 552954 194614 553574 230058
rect 552954 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 553574 194614
rect 552954 194294 553574 194378
rect 552954 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 553574 194294
rect 552954 158614 553574 194058
rect 552954 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 553574 158614
rect 552954 158294 553574 158378
rect 552954 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 553574 158294
rect 552954 122614 553574 158058
rect 552954 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 553574 122614
rect 552954 122294 553574 122378
rect 552954 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 553574 122294
rect 552954 86614 553574 122058
rect 552954 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 553574 86614
rect 552954 86294 553574 86378
rect 552954 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 553574 86294
rect 552954 50614 553574 86058
rect 552954 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 553574 50614
rect 552954 50294 553574 50378
rect 552954 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 553574 50294
rect 552954 14614 553574 50058
rect 552954 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 553574 14614
rect 552954 14294 553574 14378
rect 552954 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 553574 14294
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 14058
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 669454 560414 705242
rect 559794 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 560414 669454
rect 559794 669134 560414 669218
rect 559794 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 560414 669134
rect 559794 633454 560414 668898
rect 559794 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 560414 633454
rect 559794 633134 560414 633218
rect 559794 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 560414 633134
rect 559794 597454 560414 632898
rect 559794 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 560414 597454
rect 559794 597134 560414 597218
rect 559794 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 560414 597134
rect 559794 561454 560414 596898
rect 559794 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 560414 561454
rect 559794 561134 560414 561218
rect 559794 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 560414 561134
rect 559794 525454 560414 560898
rect 559794 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 560414 525454
rect 559794 525134 560414 525218
rect 559794 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 560414 525134
rect 559794 489454 560414 524898
rect 559794 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 560414 489454
rect 559794 489134 560414 489218
rect 559794 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 560414 489134
rect 559794 453454 560414 488898
rect 559794 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 560414 453454
rect 559794 453134 560414 453218
rect 559794 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 560414 453134
rect 559794 417454 560414 452898
rect 559794 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 560414 417454
rect 559794 417134 560414 417218
rect 559794 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 560414 417134
rect 559794 381454 560414 416898
rect 559794 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 560414 381454
rect 559794 381134 560414 381218
rect 559794 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 560414 381134
rect 559794 345454 560414 380898
rect 559794 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 560414 345454
rect 559794 345134 560414 345218
rect 559794 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 560414 345134
rect 559794 309454 560414 344898
rect 559794 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 560414 309454
rect 559794 309134 560414 309218
rect 559794 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 560414 309134
rect 559794 273454 560414 308898
rect 559794 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 560414 273454
rect 559794 273134 560414 273218
rect 559794 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 560414 273134
rect 559794 237454 560414 272898
rect 559794 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 560414 237454
rect 559794 237134 560414 237218
rect 559794 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 560414 237134
rect 559794 201454 560414 236898
rect 559794 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 560414 201454
rect 559794 201134 560414 201218
rect 559794 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 560414 201134
rect 559794 165454 560414 200898
rect 559794 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 560414 165454
rect 559794 165134 560414 165218
rect 559794 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 560414 165134
rect 559794 129454 560414 164898
rect 559794 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 560414 129454
rect 559794 129134 560414 129218
rect 559794 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 560414 129134
rect 559794 93454 560414 128898
rect 559794 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 560414 93454
rect 559794 93134 560414 93218
rect 559794 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 560414 93134
rect 559794 57454 560414 92898
rect 559794 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 560414 57454
rect 559794 57134 560414 57218
rect 559794 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 560414 57134
rect 559794 21454 560414 56898
rect 559794 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 560414 21454
rect 559794 21134 560414 21218
rect 559794 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 560414 21134
rect 559794 -1306 560414 20898
rect 559794 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 560414 -1306
rect 559794 -1626 560414 -1542
rect 559794 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 560414 -1626
rect 559794 -1894 560414 -1862
rect 563514 673174 564134 707162
rect 563514 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 564134 673174
rect 563514 672854 564134 672938
rect 563514 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 564134 672854
rect 563514 637174 564134 672618
rect 563514 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 564134 637174
rect 563514 636854 564134 636938
rect 563514 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 564134 636854
rect 563514 601174 564134 636618
rect 563514 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 564134 601174
rect 563514 600854 564134 600938
rect 563514 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 564134 600854
rect 563514 565174 564134 600618
rect 563514 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 564134 565174
rect 563514 564854 564134 564938
rect 563514 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 564134 564854
rect 563514 529174 564134 564618
rect 563514 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 564134 529174
rect 563514 528854 564134 528938
rect 563514 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 564134 528854
rect 563514 493174 564134 528618
rect 563514 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 564134 493174
rect 563514 492854 564134 492938
rect 563514 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 564134 492854
rect 563514 457174 564134 492618
rect 563514 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 564134 457174
rect 563514 456854 564134 456938
rect 563514 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 564134 456854
rect 563514 421174 564134 456618
rect 563514 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 564134 421174
rect 563514 420854 564134 420938
rect 563514 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 564134 420854
rect 563514 385174 564134 420618
rect 563514 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 564134 385174
rect 563514 384854 564134 384938
rect 563514 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 564134 384854
rect 563514 349174 564134 384618
rect 563514 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 564134 349174
rect 563514 348854 564134 348938
rect 563514 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 564134 348854
rect 563514 313174 564134 348618
rect 563514 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 564134 313174
rect 563514 312854 564134 312938
rect 563514 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 564134 312854
rect 563514 277174 564134 312618
rect 563514 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 564134 277174
rect 563514 276854 564134 276938
rect 563514 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 564134 276854
rect 563514 241174 564134 276618
rect 563514 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 564134 241174
rect 563514 240854 564134 240938
rect 563514 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 564134 240854
rect 563514 205174 564134 240618
rect 563514 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 564134 205174
rect 563514 204854 564134 204938
rect 563514 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 564134 204854
rect 563514 169174 564134 204618
rect 563514 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 564134 169174
rect 563514 168854 564134 168938
rect 563514 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 564134 168854
rect 563514 133174 564134 168618
rect 563514 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 564134 133174
rect 563514 132854 564134 132938
rect 563514 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 564134 132854
rect 563514 97174 564134 132618
rect 563514 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 564134 97174
rect 563514 96854 564134 96938
rect 563514 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 564134 96854
rect 563514 61174 564134 96618
rect 563514 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 564134 61174
rect 563514 60854 564134 60938
rect 563514 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 564134 60854
rect 563514 25174 564134 60618
rect 563514 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 564134 25174
rect 563514 24854 564134 24938
rect 563514 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 564134 24854
rect 563514 -3226 564134 24618
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 1826 687218 2062 687454
rect 2146 687218 2382 687454
rect 1826 686898 2062 687134
rect 2146 686898 2382 687134
rect 1826 651218 2062 651454
rect 2146 651218 2382 651454
rect 1826 650898 2062 651134
rect 2146 650898 2382 651134
rect 1826 615218 2062 615454
rect 2146 615218 2382 615454
rect 1826 614898 2062 615134
rect 2146 614898 2382 615134
rect 1826 579218 2062 579454
rect 2146 579218 2382 579454
rect 1826 578898 2062 579134
rect 2146 578898 2382 579134
rect 1826 543218 2062 543454
rect 2146 543218 2382 543454
rect 1826 542898 2062 543134
rect 2146 542898 2382 543134
rect 1826 507218 2062 507454
rect 2146 507218 2382 507454
rect 1826 506898 2062 507134
rect 2146 506898 2382 507134
rect 1826 471218 2062 471454
rect 2146 471218 2382 471454
rect 1826 470898 2062 471134
rect 2146 470898 2382 471134
rect 1826 435218 2062 435454
rect 2146 435218 2382 435454
rect 1826 434898 2062 435134
rect 2146 434898 2382 435134
rect 1826 399218 2062 399454
rect 2146 399218 2382 399454
rect 1826 398898 2062 399134
rect 2146 398898 2382 399134
rect 1826 363218 2062 363454
rect 2146 363218 2382 363454
rect 1826 362898 2062 363134
rect 2146 362898 2382 363134
rect 1826 327218 2062 327454
rect 2146 327218 2382 327454
rect 1826 326898 2062 327134
rect 2146 326898 2382 327134
rect 1826 291218 2062 291454
rect 2146 291218 2382 291454
rect 1826 290898 2062 291134
rect 2146 290898 2382 291134
rect 1826 255218 2062 255454
rect 2146 255218 2382 255454
rect 1826 254898 2062 255134
rect 2146 254898 2382 255134
rect 1826 219218 2062 219454
rect 2146 219218 2382 219454
rect 1826 218898 2062 219134
rect 2146 218898 2382 219134
rect 1826 183218 2062 183454
rect 2146 183218 2382 183454
rect 1826 182898 2062 183134
rect 2146 182898 2382 183134
rect 1826 147218 2062 147454
rect 2146 147218 2382 147454
rect 1826 146898 2062 147134
rect 2146 146898 2382 147134
rect 1826 111218 2062 111454
rect 2146 111218 2382 111454
rect 1826 110898 2062 111134
rect 2146 110898 2382 111134
rect 1826 75218 2062 75454
rect 2146 75218 2382 75454
rect 1826 74898 2062 75134
rect 2146 74898 2382 75134
rect 1826 39218 2062 39454
rect 2146 39218 2382 39454
rect 1826 38898 2062 39134
rect 2146 38898 2382 39134
rect 1826 3218 2062 3454
rect 2146 3218 2382 3454
rect 1826 2898 2062 3134
rect 2146 2898 2382 3134
rect 1826 -582 2062 -346
rect 2146 -582 2382 -346
rect 1826 -902 2062 -666
rect 2146 -902 2382 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect 5546 690938 5782 691174
rect 5866 690938 6102 691174
rect 5546 690618 5782 690854
rect 5866 690618 6102 690854
rect 5546 654938 5782 655174
rect 5866 654938 6102 655174
rect 5546 654618 5782 654854
rect 5866 654618 6102 654854
rect 5546 618938 5782 619174
rect 5866 618938 6102 619174
rect 5546 618618 5782 618854
rect 5866 618618 6102 618854
rect 5546 582938 5782 583174
rect 5866 582938 6102 583174
rect 5546 582618 5782 582854
rect 5866 582618 6102 582854
rect 5546 546938 5782 547174
rect 5866 546938 6102 547174
rect 5546 546618 5782 546854
rect 5866 546618 6102 546854
rect 5546 510938 5782 511174
rect 5866 510938 6102 511174
rect 5546 510618 5782 510854
rect 5866 510618 6102 510854
rect 5546 474938 5782 475174
rect 5866 474938 6102 475174
rect 5546 474618 5782 474854
rect 5866 474618 6102 474854
rect 5546 438938 5782 439174
rect 5866 438938 6102 439174
rect 5546 438618 5782 438854
rect 5866 438618 6102 438854
rect 5546 402938 5782 403174
rect 5866 402938 6102 403174
rect 5546 402618 5782 402854
rect 5866 402618 6102 402854
rect 5546 366938 5782 367174
rect 5866 366938 6102 367174
rect 5546 366618 5782 366854
rect 5866 366618 6102 366854
rect 5546 330938 5782 331174
rect 5866 330938 6102 331174
rect 5546 330618 5782 330854
rect 5866 330618 6102 330854
rect 5546 294938 5782 295174
rect 5866 294938 6102 295174
rect 5546 294618 5782 294854
rect 5866 294618 6102 294854
rect 5546 258938 5782 259174
rect 5866 258938 6102 259174
rect 5546 258618 5782 258854
rect 5866 258618 6102 258854
rect 5546 222938 5782 223174
rect 5866 222938 6102 223174
rect 5546 222618 5782 222854
rect 5866 222618 6102 222854
rect 5546 186938 5782 187174
rect 5866 186938 6102 187174
rect 5546 186618 5782 186854
rect 5866 186618 6102 186854
rect 5546 150938 5782 151174
rect 5866 150938 6102 151174
rect 5546 150618 5782 150854
rect 5866 150618 6102 150854
rect 5546 114938 5782 115174
rect 5866 114938 6102 115174
rect 5546 114618 5782 114854
rect 5866 114618 6102 114854
rect 5546 78938 5782 79174
rect 5866 78938 6102 79174
rect 5546 78618 5782 78854
rect 5866 78618 6102 78854
rect 5546 42938 5782 43174
rect 5866 42938 6102 43174
rect 5546 42618 5782 42854
rect 5866 42618 6102 42854
rect 5546 6938 5782 7174
rect 5866 6938 6102 7174
rect 5546 6618 5782 6854
rect 5866 6618 6102 6854
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect 9266 694658 9502 694894
rect 9586 694658 9822 694894
rect 9266 694338 9502 694574
rect 9586 694338 9822 694574
rect 9266 658658 9502 658894
rect 9586 658658 9822 658894
rect 9266 658338 9502 658574
rect 9586 658338 9822 658574
rect 9266 622658 9502 622894
rect 9586 622658 9822 622894
rect 9266 622338 9502 622574
rect 9586 622338 9822 622574
rect 9266 586658 9502 586894
rect 9586 586658 9822 586894
rect 9266 586338 9502 586574
rect 9586 586338 9822 586574
rect 9266 550658 9502 550894
rect 9586 550658 9822 550894
rect 9266 550338 9502 550574
rect 9586 550338 9822 550574
rect 9266 514658 9502 514894
rect 9586 514658 9822 514894
rect 9266 514338 9502 514574
rect 9586 514338 9822 514574
rect 9266 478658 9502 478894
rect 9586 478658 9822 478894
rect 9266 478338 9502 478574
rect 9586 478338 9822 478574
rect 9266 442658 9502 442894
rect 9586 442658 9822 442894
rect 9266 442338 9502 442574
rect 9586 442338 9822 442574
rect 9266 406658 9502 406894
rect 9586 406658 9822 406894
rect 9266 406338 9502 406574
rect 9586 406338 9822 406574
rect 9266 370658 9502 370894
rect 9586 370658 9822 370894
rect 9266 370338 9502 370574
rect 9586 370338 9822 370574
rect 9266 334658 9502 334894
rect 9586 334658 9822 334894
rect 9266 334338 9502 334574
rect 9586 334338 9822 334574
rect 9266 298658 9502 298894
rect 9586 298658 9822 298894
rect 9266 298338 9502 298574
rect 9586 298338 9822 298574
rect 9266 262658 9502 262894
rect 9586 262658 9822 262894
rect 9266 262338 9502 262574
rect 9586 262338 9822 262574
rect 9266 226658 9502 226894
rect 9586 226658 9822 226894
rect 9266 226338 9502 226574
rect 9586 226338 9822 226574
rect 9266 190658 9502 190894
rect 9586 190658 9822 190894
rect 9266 190338 9502 190574
rect 9586 190338 9822 190574
rect 9266 154658 9502 154894
rect 9586 154658 9822 154894
rect 9266 154338 9502 154574
rect 9586 154338 9822 154574
rect 9266 118658 9502 118894
rect 9586 118658 9822 118894
rect 9266 118338 9502 118574
rect 9586 118338 9822 118574
rect 9266 82658 9502 82894
rect 9586 82658 9822 82894
rect 9266 82338 9502 82574
rect 9586 82338 9822 82574
rect 9266 46658 9502 46894
rect 9586 46658 9822 46894
rect 9266 46338 9502 46574
rect 9586 46338 9822 46574
rect 9266 10658 9502 10894
rect 9586 10658 9822 10894
rect 9266 10338 9502 10574
rect 9586 10338 9822 10574
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 12986 698378 13222 698614
rect 13306 698378 13542 698614
rect 12986 698058 13222 698294
rect 13306 698058 13542 698294
rect 12986 662378 13222 662614
rect 13306 662378 13542 662614
rect 12986 662058 13222 662294
rect 13306 662058 13542 662294
rect 12986 626378 13222 626614
rect 13306 626378 13542 626614
rect 12986 626058 13222 626294
rect 13306 626058 13542 626294
rect 12986 590378 13222 590614
rect 13306 590378 13542 590614
rect 12986 590058 13222 590294
rect 13306 590058 13542 590294
rect 12986 554378 13222 554614
rect 13306 554378 13542 554614
rect 12986 554058 13222 554294
rect 13306 554058 13542 554294
rect 12986 518378 13222 518614
rect 13306 518378 13542 518614
rect 12986 518058 13222 518294
rect 13306 518058 13542 518294
rect 12986 482378 13222 482614
rect 13306 482378 13542 482614
rect 12986 482058 13222 482294
rect 13306 482058 13542 482294
rect 12986 446378 13222 446614
rect 13306 446378 13542 446614
rect 12986 446058 13222 446294
rect 13306 446058 13542 446294
rect 12986 410378 13222 410614
rect 13306 410378 13542 410614
rect 12986 410058 13222 410294
rect 13306 410058 13542 410294
rect 12986 374378 13222 374614
rect 13306 374378 13542 374614
rect 12986 374058 13222 374294
rect 13306 374058 13542 374294
rect 12986 338378 13222 338614
rect 13306 338378 13542 338614
rect 12986 338058 13222 338294
rect 13306 338058 13542 338294
rect 12986 302378 13222 302614
rect 13306 302378 13542 302614
rect 12986 302058 13222 302294
rect 13306 302058 13542 302294
rect 12986 266378 13222 266614
rect 13306 266378 13542 266614
rect 12986 266058 13222 266294
rect 13306 266058 13542 266294
rect 12986 230378 13222 230614
rect 13306 230378 13542 230614
rect 12986 230058 13222 230294
rect 13306 230058 13542 230294
rect 12986 194378 13222 194614
rect 13306 194378 13542 194614
rect 12986 194058 13222 194294
rect 13306 194058 13542 194294
rect 12986 158378 13222 158614
rect 13306 158378 13542 158614
rect 12986 158058 13222 158294
rect 13306 158058 13542 158294
rect 12986 122378 13222 122614
rect 13306 122378 13542 122614
rect 12986 122058 13222 122294
rect 13306 122058 13542 122294
rect 12986 86378 13222 86614
rect 13306 86378 13542 86614
rect 12986 86058 13222 86294
rect 13306 86058 13542 86294
rect 12986 50378 13222 50614
rect 13306 50378 13542 50614
rect 12986 50058 13222 50294
rect 13306 50058 13542 50294
rect 12986 14378 13222 14614
rect 13306 14378 13542 14614
rect 12986 14058 13222 14294
rect 13306 14058 13542 14294
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 19826 669218 20062 669454
rect 20146 669218 20382 669454
rect 19826 668898 20062 669134
rect 20146 668898 20382 669134
rect 19826 633218 20062 633454
rect 20146 633218 20382 633454
rect 19826 632898 20062 633134
rect 20146 632898 20382 633134
rect 19826 597218 20062 597454
rect 20146 597218 20382 597454
rect 19826 596898 20062 597134
rect 20146 596898 20382 597134
rect 19826 561218 20062 561454
rect 20146 561218 20382 561454
rect 19826 560898 20062 561134
rect 20146 560898 20382 561134
rect 19826 525218 20062 525454
rect 20146 525218 20382 525454
rect 19826 524898 20062 525134
rect 20146 524898 20382 525134
rect 19826 489218 20062 489454
rect 20146 489218 20382 489454
rect 19826 488898 20062 489134
rect 20146 488898 20382 489134
rect 19826 453218 20062 453454
rect 20146 453218 20382 453454
rect 19826 452898 20062 453134
rect 20146 452898 20382 453134
rect 19826 417218 20062 417454
rect 20146 417218 20382 417454
rect 19826 416898 20062 417134
rect 20146 416898 20382 417134
rect 19826 381218 20062 381454
rect 20146 381218 20382 381454
rect 19826 380898 20062 381134
rect 20146 380898 20382 381134
rect 19826 345218 20062 345454
rect 20146 345218 20382 345454
rect 19826 344898 20062 345134
rect 20146 344898 20382 345134
rect 19826 309218 20062 309454
rect 20146 309218 20382 309454
rect 19826 308898 20062 309134
rect 20146 308898 20382 309134
rect 19826 273218 20062 273454
rect 20146 273218 20382 273454
rect 19826 272898 20062 273134
rect 20146 272898 20382 273134
rect 19826 237218 20062 237454
rect 20146 237218 20382 237454
rect 19826 236898 20062 237134
rect 20146 236898 20382 237134
rect 19826 201218 20062 201454
rect 20146 201218 20382 201454
rect 19826 200898 20062 201134
rect 20146 200898 20382 201134
rect 19826 165218 20062 165454
rect 20146 165218 20382 165454
rect 19826 164898 20062 165134
rect 20146 164898 20382 165134
rect 19826 129218 20062 129454
rect 20146 129218 20382 129454
rect 19826 128898 20062 129134
rect 20146 128898 20382 129134
rect 19826 93218 20062 93454
rect 20146 93218 20382 93454
rect 19826 92898 20062 93134
rect 20146 92898 20382 93134
rect 19826 57218 20062 57454
rect 20146 57218 20382 57454
rect 19826 56898 20062 57134
rect 20146 56898 20382 57134
rect 19826 21218 20062 21454
rect 20146 21218 20382 21454
rect 19826 20898 20062 21134
rect 20146 20898 20382 21134
rect 19826 -1542 20062 -1306
rect 20146 -1542 20382 -1306
rect 19826 -1862 20062 -1626
rect 20146 -1862 20382 -1626
rect 23546 672938 23782 673174
rect 23866 672938 24102 673174
rect 23546 672618 23782 672854
rect 23866 672618 24102 672854
rect 23546 636938 23782 637174
rect 23866 636938 24102 637174
rect 23546 636618 23782 636854
rect 23866 636618 24102 636854
rect 23546 600938 23782 601174
rect 23866 600938 24102 601174
rect 23546 600618 23782 600854
rect 23866 600618 24102 600854
rect 23546 564938 23782 565174
rect 23866 564938 24102 565174
rect 23546 564618 23782 564854
rect 23866 564618 24102 564854
rect 23546 528938 23782 529174
rect 23866 528938 24102 529174
rect 23546 528618 23782 528854
rect 23866 528618 24102 528854
rect 23546 492938 23782 493174
rect 23866 492938 24102 493174
rect 23546 492618 23782 492854
rect 23866 492618 24102 492854
rect 23546 456938 23782 457174
rect 23866 456938 24102 457174
rect 23546 456618 23782 456854
rect 23866 456618 24102 456854
rect 23546 420938 23782 421174
rect 23866 420938 24102 421174
rect 23546 420618 23782 420854
rect 23866 420618 24102 420854
rect 23546 384938 23782 385174
rect 23866 384938 24102 385174
rect 23546 384618 23782 384854
rect 23866 384618 24102 384854
rect 23546 348938 23782 349174
rect 23866 348938 24102 349174
rect 23546 348618 23782 348854
rect 23866 348618 24102 348854
rect 23546 312938 23782 313174
rect 23866 312938 24102 313174
rect 23546 312618 23782 312854
rect 23866 312618 24102 312854
rect 23546 276938 23782 277174
rect 23866 276938 24102 277174
rect 23546 276618 23782 276854
rect 23866 276618 24102 276854
rect 23546 240938 23782 241174
rect 23866 240938 24102 241174
rect 23546 240618 23782 240854
rect 23866 240618 24102 240854
rect 23546 204938 23782 205174
rect 23866 204938 24102 205174
rect 23546 204618 23782 204854
rect 23866 204618 24102 204854
rect 23546 168938 23782 169174
rect 23866 168938 24102 169174
rect 23546 168618 23782 168854
rect 23866 168618 24102 168854
rect 23546 132938 23782 133174
rect 23866 132938 24102 133174
rect 23546 132618 23782 132854
rect 23866 132618 24102 132854
rect 23546 96938 23782 97174
rect 23866 96938 24102 97174
rect 23546 96618 23782 96854
rect 23866 96618 24102 96854
rect 23546 60938 23782 61174
rect 23866 60938 24102 61174
rect 23546 60618 23782 60854
rect 23866 60618 24102 60854
rect 23546 24938 23782 25174
rect 23866 24938 24102 25174
rect 23546 24618 23782 24854
rect 23866 24618 24102 24854
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 676658 27502 676894
rect 27586 676658 27822 676894
rect 27266 676338 27502 676574
rect 27586 676338 27822 676574
rect 27266 640658 27502 640894
rect 27586 640658 27822 640894
rect 27266 640338 27502 640574
rect 27586 640338 27822 640574
rect 27266 604658 27502 604894
rect 27586 604658 27822 604894
rect 27266 604338 27502 604574
rect 27586 604338 27822 604574
rect 27266 568658 27502 568894
rect 27586 568658 27822 568894
rect 27266 568338 27502 568574
rect 27586 568338 27822 568574
rect 27266 532658 27502 532894
rect 27586 532658 27822 532894
rect 27266 532338 27502 532574
rect 27586 532338 27822 532574
rect 27266 496658 27502 496894
rect 27586 496658 27822 496894
rect 27266 496338 27502 496574
rect 27586 496338 27822 496574
rect 27266 460658 27502 460894
rect 27586 460658 27822 460894
rect 27266 460338 27502 460574
rect 27586 460338 27822 460574
rect 27266 424658 27502 424894
rect 27586 424658 27822 424894
rect 27266 424338 27502 424574
rect 27586 424338 27822 424574
rect 27266 388658 27502 388894
rect 27586 388658 27822 388894
rect 27266 388338 27502 388574
rect 27586 388338 27822 388574
rect 27266 352658 27502 352894
rect 27586 352658 27822 352894
rect 27266 352338 27502 352574
rect 27586 352338 27822 352574
rect 27266 316658 27502 316894
rect 27586 316658 27822 316894
rect 27266 316338 27502 316574
rect 27586 316338 27822 316574
rect 27266 280658 27502 280894
rect 27586 280658 27822 280894
rect 27266 280338 27502 280574
rect 27586 280338 27822 280574
rect 27266 244658 27502 244894
rect 27586 244658 27822 244894
rect 27266 244338 27502 244574
rect 27586 244338 27822 244574
rect 27266 208658 27502 208894
rect 27586 208658 27822 208894
rect 27266 208338 27502 208574
rect 27586 208338 27822 208574
rect 27266 172658 27502 172894
rect 27586 172658 27822 172894
rect 27266 172338 27502 172574
rect 27586 172338 27822 172574
rect 27266 136658 27502 136894
rect 27586 136658 27822 136894
rect 27266 136338 27502 136574
rect 27586 136338 27822 136574
rect 27266 100658 27502 100894
rect 27586 100658 27822 100894
rect 27266 100338 27502 100574
rect 27586 100338 27822 100574
rect 27266 64658 27502 64894
rect 27586 64658 27822 64894
rect 27266 64338 27502 64574
rect 27586 64338 27822 64574
rect 27266 28658 27502 28894
rect 27586 28658 27822 28894
rect 27266 28338 27502 28574
rect 27586 28338 27822 28574
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 30986 680378 31222 680614
rect 31306 680378 31542 680614
rect 30986 680058 31222 680294
rect 31306 680058 31542 680294
rect 30986 644378 31222 644614
rect 31306 644378 31542 644614
rect 30986 644058 31222 644294
rect 31306 644058 31542 644294
rect 30986 608378 31222 608614
rect 31306 608378 31542 608614
rect 30986 608058 31222 608294
rect 31306 608058 31542 608294
rect 30986 572378 31222 572614
rect 31306 572378 31542 572614
rect 30986 572058 31222 572294
rect 31306 572058 31542 572294
rect 30986 536378 31222 536614
rect 31306 536378 31542 536614
rect 30986 536058 31222 536294
rect 31306 536058 31542 536294
rect 30986 500378 31222 500614
rect 31306 500378 31542 500614
rect 30986 500058 31222 500294
rect 31306 500058 31542 500294
rect 30986 464378 31222 464614
rect 31306 464378 31542 464614
rect 30986 464058 31222 464294
rect 31306 464058 31542 464294
rect 30986 428378 31222 428614
rect 31306 428378 31542 428614
rect 30986 428058 31222 428294
rect 31306 428058 31542 428294
rect 30986 392378 31222 392614
rect 31306 392378 31542 392614
rect 30986 392058 31222 392294
rect 31306 392058 31542 392294
rect 30986 356378 31222 356614
rect 31306 356378 31542 356614
rect 30986 356058 31222 356294
rect 31306 356058 31542 356294
rect 30986 320378 31222 320614
rect 31306 320378 31542 320614
rect 30986 320058 31222 320294
rect 31306 320058 31542 320294
rect 30986 284378 31222 284614
rect 31306 284378 31542 284614
rect 30986 284058 31222 284294
rect 31306 284058 31542 284294
rect 30986 248378 31222 248614
rect 31306 248378 31542 248614
rect 30986 248058 31222 248294
rect 31306 248058 31542 248294
rect 30986 212378 31222 212614
rect 31306 212378 31542 212614
rect 30986 212058 31222 212294
rect 31306 212058 31542 212294
rect 30986 176378 31222 176614
rect 31306 176378 31542 176614
rect 30986 176058 31222 176294
rect 31306 176058 31542 176294
rect 30986 140378 31222 140614
rect 31306 140378 31542 140614
rect 30986 140058 31222 140294
rect 31306 140058 31542 140294
rect 30986 104378 31222 104614
rect 31306 104378 31542 104614
rect 30986 104058 31222 104294
rect 31306 104058 31542 104294
rect 30986 68378 31222 68614
rect 31306 68378 31542 68614
rect 30986 68058 31222 68294
rect 31306 68058 31542 68294
rect 30986 32378 31222 32614
rect 31306 32378 31542 32614
rect 30986 32058 31222 32294
rect 31306 32058 31542 32294
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 37826 687218 38062 687454
rect 38146 687218 38382 687454
rect 37826 686898 38062 687134
rect 38146 686898 38382 687134
rect 37826 651218 38062 651454
rect 38146 651218 38382 651454
rect 37826 650898 38062 651134
rect 38146 650898 38382 651134
rect 37826 615218 38062 615454
rect 38146 615218 38382 615454
rect 37826 614898 38062 615134
rect 38146 614898 38382 615134
rect 37826 579218 38062 579454
rect 38146 579218 38382 579454
rect 37826 578898 38062 579134
rect 38146 578898 38382 579134
rect 37826 543218 38062 543454
rect 38146 543218 38382 543454
rect 37826 542898 38062 543134
rect 38146 542898 38382 543134
rect 37826 507218 38062 507454
rect 38146 507218 38382 507454
rect 37826 506898 38062 507134
rect 38146 506898 38382 507134
rect 37826 471218 38062 471454
rect 38146 471218 38382 471454
rect 37826 470898 38062 471134
rect 38146 470898 38382 471134
rect 37826 435218 38062 435454
rect 38146 435218 38382 435454
rect 37826 434898 38062 435134
rect 38146 434898 38382 435134
rect 37826 399218 38062 399454
rect 38146 399218 38382 399454
rect 37826 398898 38062 399134
rect 38146 398898 38382 399134
rect 37826 363218 38062 363454
rect 38146 363218 38382 363454
rect 37826 362898 38062 363134
rect 38146 362898 38382 363134
rect 37826 327218 38062 327454
rect 38146 327218 38382 327454
rect 37826 326898 38062 327134
rect 38146 326898 38382 327134
rect 37826 291218 38062 291454
rect 38146 291218 38382 291454
rect 37826 290898 38062 291134
rect 38146 290898 38382 291134
rect 37826 255218 38062 255454
rect 38146 255218 38382 255454
rect 37826 254898 38062 255134
rect 38146 254898 38382 255134
rect 37826 219218 38062 219454
rect 38146 219218 38382 219454
rect 37826 218898 38062 219134
rect 38146 218898 38382 219134
rect 37826 183218 38062 183454
rect 38146 183218 38382 183454
rect 37826 182898 38062 183134
rect 38146 182898 38382 183134
rect 37826 147218 38062 147454
rect 38146 147218 38382 147454
rect 37826 146898 38062 147134
rect 38146 146898 38382 147134
rect 37826 111218 38062 111454
rect 38146 111218 38382 111454
rect 37826 110898 38062 111134
rect 38146 110898 38382 111134
rect 37826 75218 38062 75454
rect 38146 75218 38382 75454
rect 37826 74898 38062 75134
rect 38146 74898 38382 75134
rect 37826 39218 38062 39454
rect 38146 39218 38382 39454
rect 37826 38898 38062 39134
rect 38146 38898 38382 39134
rect 37826 3218 38062 3454
rect 38146 3218 38382 3454
rect 37826 2898 38062 3134
rect 38146 2898 38382 3134
rect 37826 -582 38062 -346
rect 38146 -582 38382 -346
rect 37826 -902 38062 -666
rect 38146 -902 38382 -666
rect 41546 690938 41782 691174
rect 41866 690938 42102 691174
rect 41546 690618 41782 690854
rect 41866 690618 42102 690854
rect 41546 654938 41782 655174
rect 41866 654938 42102 655174
rect 41546 654618 41782 654854
rect 41866 654618 42102 654854
rect 41546 618938 41782 619174
rect 41866 618938 42102 619174
rect 41546 618618 41782 618854
rect 41866 618618 42102 618854
rect 41546 582938 41782 583174
rect 41866 582938 42102 583174
rect 41546 582618 41782 582854
rect 41866 582618 42102 582854
rect 41546 546938 41782 547174
rect 41866 546938 42102 547174
rect 41546 546618 41782 546854
rect 41866 546618 42102 546854
rect 41546 510938 41782 511174
rect 41866 510938 42102 511174
rect 41546 510618 41782 510854
rect 41866 510618 42102 510854
rect 41546 474938 41782 475174
rect 41866 474938 42102 475174
rect 41546 474618 41782 474854
rect 41866 474618 42102 474854
rect 41546 438938 41782 439174
rect 41866 438938 42102 439174
rect 41546 438618 41782 438854
rect 41866 438618 42102 438854
rect 41546 402938 41782 403174
rect 41866 402938 42102 403174
rect 41546 402618 41782 402854
rect 41866 402618 42102 402854
rect 41546 366938 41782 367174
rect 41866 366938 42102 367174
rect 41546 366618 41782 366854
rect 41866 366618 42102 366854
rect 41546 330938 41782 331174
rect 41866 330938 42102 331174
rect 41546 330618 41782 330854
rect 41866 330618 42102 330854
rect 41546 294938 41782 295174
rect 41866 294938 42102 295174
rect 41546 294618 41782 294854
rect 41866 294618 42102 294854
rect 41546 258938 41782 259174
rect 41866 258938 42102 259174
rect 41546 258618 41782 258854
rect 41866 258618 42102 258854
rect 41546 222938 41782 223174
rect 41866 222938 42102 223174
rect 41546 222618 41782 222854
rect 41866 222618 42102 222854
rect 41546 186938 41782 187174
rect 41866 186938 42102 187174
rect 41546 186618 41782 186854
rect 41866 186618 42102 186854
rect 41546 150938 41782 151174
rect 41866 150938 42102 151174
rect 41546 150618 41782 150854
rect 41866 150618 42102 150854
rect 41546 114938 41782 115174
rect 41866 114938 42102 115174
rect 41546 114618 41782 114854
rect 41866 114618 42102 114854
rect 41546 78938 41782 79174
rect 41866 78938 42102 79174
rect 41546 78618 41782 78854
rect 41866 78618 42102 78854
rect 41546 42938 41782 43174
rect 41866 42938 42102 43174
rect 41546 42618 41782 42854
rect 41866 42618 42102 42854
rect 41546 6938 41782 7174
rect 41866 6938 42102 7174
rect 41546 6618 41782 6854
rect 41866 6618 42102 6854
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 694658 45502 694894
rect 45586 694658 45822 694894
rect 45266 694338 45502 694574
rect 45586 694338 45822 694574
rect 45266 658658 45502 658894
rect 45586 658658 45822 658894
rect 45266 658338 45502 658574
rect 45586 658338 45822 658574
rect 45266 622658 45502 622894
rect 45586 622658 45822 622894
rect 45266 622338 45502 622574
rect 45586 622338 45822 622574
rect 45266 586658 45502 586894
rect 45586 586658 45822 586894
rect 45266 586338 45502 586574
rect 45586 586338 45822 586574
rect 45266 550658 45502 550894
rect 45586 550658 45822 550894
rect 45266 550338 45502 550574
rect 45586 550338 45822 550574
rect 45266 514658 45502 514894
rect 45586 514658 45822 514894
rect 45266 514338 45502 514574
rect 45586 514338 45822 514574
rect 45266 478658 45502 478894
rect 45586 478658 45822 478894
rect 45266 478338 45502 478574
rect 45586 478338 45822 478574
rect 45266 442658 45502 442894
rect 45586 442658 45822 442894
rect 45266 442338 45502 442574
rect 45586 442338 45822 442574
rect 45266 406658 45502 406894
rect 45586 406658 45822 406894
rect 45266 406338 45502 406574
rect 45586 406338 45822 406574
rect 45266 370658 45502 370894
rect 45586 370658 45822 370894
rect 45266 370338 45502 370574
rect 45586 370338 45822 370574
rect 45266 334658 45502 334894
rect 45586 334658 45822 334894
rect 45266 334338 45502 334574
rect 45586 334338 45822 334574
rect 45266 298658 45502 298894
rect 45586 298658 45822 298894
rect 45266 298338 45502 298574
rect 45586 298338 45822 298574
rect 45266 262658 45502 262894
rect 45586 262658 45822 262894
rect 45266 262338 45502 262574
rect 45586 262338 45822 262574
rect 45266 226658 45502 226894
rect 45586 226658 45822 226894
rect 45266 226338 45502 226574
rect 45586 226338 45822 226574
rect 45266 190658 45502 190894
rect 45586 190658 45822 190894
rect 45266 190338 45502 190574
rect 45586 190338 45822 190574
rect 45266 154658 45502 154894
rect 45586 154658 45822 154894
rect 45266 154338 45502 154574
rect 45586 154338 45822 154574
rect 45266 118658 45502 118894
rect 45586 118658 45822 118894
rect 45266 118338 45502 118574
rect 45586 118338 45822 118574
rect 45266 82658 45502 82894
rect 45586 82658 45822 82894
rect 45266 82338 45502 82574
rect 45586 82338 45822 82574
rect 45266 46658 45502 46894
rect 45586 46658 45822 46894
rect 45266 46338 45502 46574
rect 45586 46338 45822 46574
rect 45266 10658 45502 10894
rect 45586 10658 45822 10894
rect 45266 10338 45502 10574
rect 45586 10338 45822 10574
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 48986 698378 49222 698614
rect 49306 698378 49542 698614
rect 48986 698058 49222 698294
rect 49306 698058 49542 698294
rect 48986 662378 49222 662614
rect 49306 662378 49542 662614
rect 48986 662058 49222 662294
rect 49306 662058 49542 662294
rect 48986 626378 49222 626614
rect 49306 626378 49542 626614
rect 48986 626058 49222 626294
rect 49306 626058 49542 626294
rect 48986 590378 49222 590614
rect 49306 590378 49542 590614
rect 48986 590058 49222 590294
rect 49306 590058 49542 590294
rect 48986 554378 49222 554614
rect 49306 554378 49542 554614
rect 48986 554058 49222 554294
rect 49306 554058 49542 554294
rect 48986 518378 49222 518614
rect 49306 518378 49542 518614
rect 48986 518058 49222 518294
rect 49306 518058 49542 518294
rect 48986 482378 49222 482614
rect 49306 482378 49542 482614
rect 48986 482058 49222 482294
rect 49306 482058 49542 482294
rect 48986 446378 49222 446614
rect 49306 446378 49542 446614
rect 48986 446058 49222 446294
rect 49306 446058 49542 446294
rect 48986 410378 49222 410614
rect 49306 410378 49542 410614
rect 48986 410058 49222 410294
rect 49306 410058 49542 410294
rect 48986 374378 49222 374614
rect 49306 374378 49542 374614
rect 48986 374058 49222 374294
rect 49306 374058 49542 374294
rect 48986 338378 49222 338614
rect 49306 338378 49542 338614
rect 48986 338058 49222 338294
rect 49306 338058 49542 338294
rect 48986 302378 49222 302614
rect 49306 302378 49542 302614
rect 48986 302058 49222 302294
rect 49306 302058 49542 302294
rect 48986 266378 49222 266614
rect 49306 266378 49542 266614
rect 48986 266058 49222 266294
rect 49306 266058 49542 266294
rect 48986 230378 49222 230614
rect 49306 230378 49542 230614
rect 48986 230058 49222 230294
rect 49306 230058 49542 230294
rect 48986 194378 49222 194614
rect 49306 194378 49542 194614
rect 48986 194058 49222 194294
rect 49306 194058 49542 194294
rect 48986 158378 49222 158614
rect 49306 158378 49542 158614
rect 48986 158058 49222 158294
rect 49306 158058 49542 158294
rect 48986 122378 49222 122614
rect 49306 122378 49542 122614
rect 48986 122058 49222 122294
rect 49306 122058 49542 122294
rect 48986 86378 49222 86614
rect 49306 86378 49542 86614
rect 48986 86058 49222 86294
rect 49306 86058 49542 86294
rect 48986 50378 49222 50614
rect 49306 50378 49542 50614
rect 48986 50058 49222 50294
rect 49306 50058 49542 50294
rect 48986 14378 49222 14614
rect 49306 14378 49542 14614
rect 48986 14058 49222 14294
rect 49306 14058 49542 14294
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 55826 669218 56062 669454
rect 56146 669218 56382 669454
rect 55826 668898 56062 669134
rect 56146 668898 56382 669134
rect 55826 633218 56062 633454
rect 56146 633218 56382 633454
rect 55826 632898 56062 633134
rect 56146 632898 56382 633134
rect 55826 597218 56062 597454
rect 56146 597218 56382 597454
rect 55826 596898 56062 597134
rect 56146 596898 56382 597134
rect 55826 561218 56062 561454
rect 56146 561218 56382 561454
rect 55826 560898 56062 561134
rect 56146 560898 56382 561134
rect 55826 525218 56062 525454
rect 56146 525218 56382 525454
rect 55826 524898 56062 525134
rect 56146 524898 56382 525134
rect 55826 489218 56062 489454
rect 56146 489218 56382 489454
rect 55826 488898 56062 489134
rect 56146 488898 56382 489134
rect 59546 672938 59782 673174
rect 59866 672938 60102 673174
rect 59546 672618 59782 672854
rect 59866 672618 60102 672854
rect 59546 636938 59782 637174
rect 59866 636938 60102 637174
rect 59546 636618 59782 636854
rect 59866 636618 60102 636854
rect 59546 600938 59782 601174
rect 59866 600938 60102 601174
rect 59546 600618 59782 600854
rect 59866 600618 60102 600854
rect 59546 564938 59782 565174
rect 59866 564938 60102 565174
rect 59546 564618 59782 564854
rect 59866 564618 60102 564854
rect 59546 528938 59782 529174
rect 59866 528938 60102 529174
rect 59546 528618 59782 528854
rect 59866 528618 60102 528854
rect 59546 492938 59782 493174
rect 59866 492938 60102 493174
rect 59546 492618 59782 492854
rect 59866 492618 60102 492854
rect 63266 676658 63502 676894
rect 63586 676658 63822 676894
rect 63266 676338 63502 676574
rect 63586 676338 63822 676574
rect 63266 640658 63502 640894
rect 63586 640658 63822 640894
rect 63266 640338 63502 640574
rect 63586 640338 63822 640574
rect 63266 604658 63502 604894
rect 63586 604658 63822 604894
rect 63266 604338 63502 604574
rect 63586 604338 63822 604574
rect 63266 568658 63502 568894
rect 63586 568658 63822 568894
rect 63266 568338 63502 568574
rect 63586 568338 63822 568574
rect 63266 532658 63502 532894
rect 63586 532658 63822 532894
rect 63266 532338 63502 532574
rect 63586 532338 63822 532574
rect 63266 496658 63502 496894
rect 63586 496658 63822 496894
rect 63266 496338 63502 496574
rect 63586 496338 63822 496574
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 66986 680378 67222 680614
rect 67306 680378 67542 680614
rect 66986 680058 67222 680294
rect 67306 680058 67542 680294
rect 66986 644378 67222 644614
rect 67306 644378 67542 644614
rect 66986 644058 67222 644294
rect 67306 644058 67542 644294
rect 66986 608378 67222 608614
rect 67306 608378 67542 608614
rect 66986 608058 67222 608294
rect 67306 608058 67542 608294
rect 66986 572378 67222 572614
rect 67306 572378 67542 572614
rect 66986 572058 67222 572294
rect 67306 572058 67542 572294
rect 66986 536378 67222 536614
rect 67306 536378 67542 536614
rect 66986 536058 67222 536294
rect 67306 536058 67542 536294
rect 66986 500378 67222 500614
rect 67306 500378 67542 500614
rect 66986 500058 67222 500294
rect 67306 500058 67542 500294
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 73826 687218 74062 687454
rect 74146 687218 74382 687454
rect 73826 686898 74062 687134
rect 74146 686898 74382 687134
rect 73826 651218 74062 651454
rect 74146 651218 74382 651454
rect 73826 650898 74062 651134
rect 74146 650898 74382 651134
rect 73826 615218 74062 615454
rect 74146 615218 74382 615454
rect 73826 614898 74062 615134
rect 74146 614898 74382 615134
rect 73826 579218 74062 579454
rect 74146 579218 74382 579454
rect 73826 578898 74062 579134
rect 74146 578898 74382 579134
rect 73826 543218 74062 543454
rect 74146 543218 74382 543454
rect 73826 542898 74062 543134
rect 74146 542898 74382 543134
rect 73826 507218 74062 507454
rect 74146 507218 74382 507454
rect 73826 506898 74062 507134
rect 74146 506898 74382 507134
rect 77546 690938 77782 691174
rect 77866 690938 78102 691174
rect 77546 690618 77782 690854
rect 77866 690618 78102 690854
rect 77546 654938 77782 655174
rect 77866 654938 78102 655174
rect 77546 654618 77782 654854
rect 77866 654618 78102 654854
rect 77546 618938 77782 619174
rect 77866 618938 78102 619174
rect 77546 618618 77782 618854
rect 77866 618618 78102 618854
rect 77546 582938 77782 583174
rect 77866 582938 78102 583174
rect 77546 582618 77782 582854
rect 77866 582618 78102 582854
rect 77546 546938 77782 547174
rect 77866 546938 78102 547174
rect 77546 546618 77782 546854
rect 77866 546618 78102 546854
rect 77546 510938 77782 511174
rect 77866 510938 78102 511174
rect 77546 510618 77782 510854
rect 77866 510618 78102 510854
rect 81266 694658 81502 694894
rect 81586 694658 81822 694894
rect 81266 694338 81502 694574
rect 81586 694338 81822 694574
rect 81266 658658 81502 658894
rect 81586 658658 81822 658894
rect 81266 658338 81502 658574
rect 81586 658338 81822 658574
rect 81266 622658 81502 622894
rect 81586 622658 81822 622894
rect 81266 622338 81502 622574
rect 81586 622338 81822 622574
rect 81266 586658 81502 586894
rect 81586 586658 81822 586894
rect 81266 586338 81502 586574
rect 81586 586338 81822 586574
rect 81266 550658 81502 550894
rect 81586 550658 81822 550894
rect 81266 550338 81502 550574
rect 81586 550338 81822 550574
rect 81266 514658 81502 514894
rect 81586 514658 81822 514894
rect 81266 514338 81502 514574
rect 81586 514338 81822 514574
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 84986 698378 85222 698614
rect 85306 698378 85542 698614
rect 84986 698058 85222 698294
rect 85306 698058 85542 698294
rect 84986 662378 85222 662614
rect 85306 662378 85542 662614
rect 84986 662058 85222 662294
rect 85306 662058 85542 662294
rect 84986 626378 85222 626614
rect 85306 626378 85542 626614
rect 84986 626058 85222 626294
rect 85306 626058 85542 626294
rect 84986 590378 85222 590614
rect 85306 590378 85542 590614
rect 84986 590058 85222 590294
rect 85306 590058 85542 590294
rect 84986 554378 85222 554614
rect 85306 554378 85542 554614
rect 84986 554058 85222 554294
rect 85306 554058 85542 554294
rect 84986 518378 85222 518614
rect 85306 518378 85542 518614
rect 84986 518058 85222 518294
rect 85306 518058 85542 518294
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 91826 669218 92062 669454
rect 92146 669218 92382 669454
rect 91826 668898 92062 669134
rect 92146 668898 92382 669134
rect 91826 633218 92062 633454
rect 92146 633218 92382 633454
rect 91826 632898 92062 633134
rect 92146 632898 92382 633134
rect 91826 597218 92062 597454
rect 92146 597218 92382 597454
rect 91826 596898 92062 597134
rect 92146 596898 92382 597134
rect 91826 561218 92062 561454
rect 92146 561218 92382 561454
rect 91826 560898 92062 561134
rect 92146 560898 92382 561134
rect 91826 525218 92062 525454
rect 92146 525218 92382 525454
rect 91826 524898 92062 525134
rect 92146 524898 92382 525134
rect 91826 489218 92062 489454
rect 92146 489218 92382 489454
rect 91826 488898 92062 489134
rect 92146 488898 92382 489134
rect 95546 672938 95782 673174
rect 95866 672938 96102 673174
rect 95546 672618 95782 672854
rect 95866 672618 96102 672854
rect 95546 636938 95782 637174
rect 95866 636938 96102 637174
rect 95546 636618 95782 636854
rect 95866 636618 96102 636854
rect 95546 600938 95782 601174
rect 95866 600938 96102 601174
rect 95546 600618 95782 600854
rect 95866 600618 96102 600854
rect 95546 564938 95782 565174
rect 95866 564938 96102 565174
rect 95546 564618 95782 564854
rect 95866 564618 96102 564854
rect 95546 528938 95782 529174
rect 95866 528938 96102 529174
rect 95546 528618 95782 528854
rect 95866 528618 96102 528854
rect 95546 492938 95782 493174
rect 95866 492938 96102 493174
rect 95546 492618 95782 492854
rect 95866 492618 96102 492854
rect 99266 676658 99502 676894
rect 99586 676658 99822 676894
rect 99266 676338 99502 676574
rect 99586 676338 99822 676574
rect 99266 640658 99502 640894
rect 99586 640658 99822 640894
rect 99266 640338 99502 640574
rect 99586 640338 99822 640574
rect 99266 604658 99502 604894
rect 99586 604658 99822 604894
rect 99266 604338 99502 604574
rect 99586 604338 99822 604574
rect 99266 568658 99502 568894
rect 99586 568658 99822 568894
rect 99266 568338 99502 568574
rect 99586 568338 99822 568574
rect 99266 532658 99502 532894
rect 99586 532658 99822 532894
rect 99266 532338 99502 532574
rect 99586 532338 99822 532574
rect 99266 496658 99502 496894
rect 99586 496658 99822 496894
rect 99266 496338 99502 496574
rect 99586 496338 99822 496574
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 102986 680378 103222 680614
rect 103306 680378 103542 680614
rect 102986 680058 103222 680294
rect 103306 680058 103542 680294
rect 102986 644378 103222 644614
rect 103306 644378 103542 644614
rect 102986 644058 103222 644294
rect 103306 644058 103542 644294
rect 102986 608378 103222 608614
rect 103306 608378 103542 608614
rect 102986 608058 103222 608294
rect 103306 608058 103542 608294
rect 102986 572378 103222 572614
rect 103306 572378 103542 572614
rect 102986 572058 103222 572294
rect 103306 572058 103542 572294
rect 102986 536378 103222 536614
rect 103306 536378 103542 536614
rect 102986 536058 103222 536294
rect 103306 536058 103542 536294
rect 102986 500378 103222 500614
rect 103306 500378 103542 500614
rect 102986 500058 103222 500294
rect 103306 500058 103542 500294
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 109826 687218 110062 687454
rect 110146 687218 110382 687454
rect 109826 686898 110062 687134
rect 110146 686898 110382 687134
rect 109826 651218 110062 651454
rect 110146 651218 110382 651454
rect 109826 650898 110062 651134
rect 110146 650898 110382 651134
rect 109826 615218 110062 615454
rect 110146 615218 110382 615454
rect 109826 614898 110062 615134
rect 110146 614898 110382 615134
rect 109826 579218 110062 579454
rect 110146 579218 110382 579454
rect 109826 578898 110062 579134
rect 110146 578898 110382 579134
rect 109826 543218 110062 543454
rect 110146 543218 110382 543454
rect 109826 542898 110062 543134
rect 110146 542898 110382 543134
rect 109826 507218 110062 507454
rect 110146 507218 110382 507454
rect 109826 506898 110062 507134
rect 110146 506898 110382 507134
rect 113546 690938 113782 691174
rect 113866 690938 114102 691174
rect 113546 690618 113782 690854
rect 113866 690618 114102 690854
rect 113546 654938 113782 655174
rect 113866 654938 114102 655174
rect 113546 654618 113782 654854
rect 113866 654618 114102 654854
rect 113546 618938 113782 619174
rect 113866 618938 114102 619174
rect 113546 618618 113782 618854
rect 113866 618618 114102 618854
rect 113546 582938 113782 583174
rect 113866 582938 114102 583174
rect 113546 582618 113782 582854
rect 113866 582618 114102 582854
rect 113546 546938 113782 547174
rect 113866 546938 114102 547174
rect 113546 546618 113782 546854
rect 113866 546618 114102 546854
rect 113546 510938 113782 511174
rect 113866 510938 114102 511174
rect 113546 510618 113782 510854
rect 113866 510618 114102 510854
rect 117266 694658 117502 694894
rect 117586 694658 117822 694894
rect 117266 694338 117502 694574
rect 117586 694338 117822 694574
rect 117266 658658 117502 658894
rect 117586 658658 117822 658894
rect 117266 658338 117502 658574
rect 117586 658338 117822 658574
rect 117266 622658 117502 622894
rect 117586 622658 117822 622894
rect 117266 622338 117502 622574
rect 117586 622338 117822 622574
rect 117266 586658 117502 586894
rect 117586 586658 117822 586894
rect 117266 586338 117502 586574
rect 117586 586338 117822 586574
rect 117266 550658 117502 550894
rect 117586 550658 117822 550894
rect 117266 550338 117502 550574
rect 117586 550338 117822 550574
rect 117266 514658 117502 514894
rect 117586 514658 117822 514894
rect 117266 514338 117502 514574
rect 117586 514338 117822 514574
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 120986 698378 121222 698614
rect 121306 698378 121542 698614
rect 120986 698058 121222 698294
rect 121306 698058 121542 698294
rect 120986 662378 121222 662614
rect 121306 662378 121542 662614
rect 120986 662058 121222 662294
rect 121306 662058 121542 662294
rect 120986 626378 121222 626614
rect 121306 626378 121542 626614
rect 120986 626058 121222 626294
rect 121306 626058 121542 626294
rect 120986 590378 121222 590614
rect 121306 590378 121542 590614
rect 120986 590058 121222 590294
rect 121306 590058 121542 590294
rect 120986 554378 121222 554614
rect 121306 554378 121542 554614
rect 120986 554058 121222 554294
rect 121306 554058 121542 554294
rect 120986 518378 121222 518614
rect 121306 518378 121542 518614
rect 120986 518058 121222 518294
rect 121306 518058 121542 518294
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 127826 669218 128062 669454
rect 128146 669218 128382 669454
rect 127826 668898 128062 669134
rect 128146 668898 128382 669134
rect 127826 633218 128062 633454
rect 128146 633218 128382 633454
rect 127826 632898 128062 633134
rect 128146 632898 128382 633134
rect 127826 597218 128062 597454
rect 128146 597218 128382 597454
rect 127826 596898 128062 597134
rect 128146 596898 128382 597134
rect 127826 561218 128062 561454
rect 128146 561218 128382 561454
rect 127826 560898 128062 561134
rect 128146 560898 128382 561134
rect 127826 525218 128062 525454
rect 128146 525218 128382 525454
rect 127826 524898 128062 525134
rect 128146 524898 128382 525134
rect 127826 489218 128062 489454
rect 128146 489218 128382 489454
rect 127826 488898 128062 489134
rect 128146 488898 128382 489134
rect 131546 672938 131782 673174
rect 131866 672938 132102 673174
rect 131546 672618 131782 672854
rect 131866 672618 132102 672854
rect 131546 636938 131782 637174
rect 131866 636938 132102 637174
rect 131546 636618 131782 636854
rect 131866 636618 132102 636854
rect 131546 600938 131782 601174
rect 131866 600938 132102 601174
rect 131546 600618 131782 600854
rect 131866 600618 132102 600854
rect 131546 564938 131782 565174
rect 131866 564938 132102 565174
rect 131546 564618 131782 564854
rect 131866 564618 132102 564854
rect 131546 528938 131782 529174
rect 131866 528938 132102 529174
rect 131546 528618 131782 528854
rect 131866 528618 132102 528854
rect 131546 492938 131782 493174
rect 131866 492938 132102 493174
rect 131546 492618 131782 492854
rect 131866 492618 132102 492854
rect 135266 676658 135502 676894
rect 135586 676658 135822 676894
rect 135266 676338 135502 676574
rect 135586 676338 135822 676574
rect 135266 640658 135502 640894
rect 135586 640658 135822 640894
rect 135266 640338 135502 640574
rect 135586 640338 135822 640574
rect 135266 604658 135502 604894
rect 135586 604658 135822 604894
rect 135266 604338 135502 604574
rect 135586 604338 135822 604574
rect 135266 568658 135502 568894
rect 135586 568658 135822 568894
rect 135266 568338 135502 568574
rect 135586 568338 135822 568574
rect 135266 532658 135502 532894
rect 135586 532658 135822 532894
rect 135266 532338 135502 532574
rect 135586 532338 135822 532574
rect 135266 496658 135502 496894
rect 135586 496658 135822 496894
rect 135266 496338 135502 496574
rect 135586 496338 135822 496574
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 138986 680378 139222 680614
rect 139306 680378 139542 680614
rect 138986 680058 139222 680294
rect 139306 680058 139542 680294
rect 138986 644378 139222 644614
rect 139306 644378 139542 644614
rect 138986 644058 139222 644294
rect 139306 644058 139542 644294
rect 138986 608378 139222 608614
rect 139306 608378 139542 608614
rect 138986 608058 139222 608294
rect 139306 608058 139542 608294
rect 138986 572378 139222 572614
rect 139306 572378 139542 572614
rect 138986 572058 139222 572294
rect 139306 572058 139542 572294
rect 138986 536378 139222 536614
rect 139306 536378 139542 536614
rect 138986 536058 139222 536294
rect 139306 536058 139542 536294
rect 138986 500378 139222 500614
rect 139306 500378 139542 500614
rect 138986 500058 139222 500294
rect 139306 500058 139542 500294
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 145826 687218 146062 687454
rect 146146 687218 146382 687454
rect 145826 686898 146062 687134
rect 146146 686898 146382 687134
rect 145826 651218 146062 651454
rect 146146 651218 146382 651454
rect 145826 650898 146062 651134
rect 146146 650898 146382 651134
rect 145826 615218 146062 615454
rect 146146 615218 146382 615454
rect 145826 614898 146062 615134
rect 146146 614898 146382 615134
rect 145826 579218 146062 579454
rect 146146 579218 146382 579454
rect 145826 578898 146062 579134
rect 146146 578898 146382 579134
rect 145826 543218 146062 543454
rect 146146 543218 146382 543454
rect 145826 542898 146062 543134
rect 146146 542898 146382 543134
rect 145826 507218 146062 507454
rect 146146 507218 146382 507454
rect 145826 506898 146062 507134
rect 146146 506898 146382 507134
rect 149546 690938 149782 691174
rect 149866 690938 150102 691174
rect 149546 690618 149782 690854
rect 149866 690618 150102 690854
rect 149546 654938 149782 655174
rect 149866 654938 150102 655174
rect 149546 654618 149782 654854
rect 149866 654618 150102 654854
rect 149546 618938 149782 619174
rect 149866 618938 150102 619174
rect 149546 618618 149782 618854
rect 149866 618618 150102 618854
rect 149546 582938 149782 583174
rect 149866 582938 150102 583174
rect 149546 582618 149782 582854
rect 149866 582618 150102 582854
rect 149546 546938 149782 547174
rect 149866 546938 150102 547174
rect 149546 546618 149782 546854
rect 149866 546618 150102 546854
rect 149546 510938 149782 511174
rect 149866 510938 150102 511174
rect 149546 510618 149782 510854
rect 149866 510618 150102 510854
rect 153266 694658 153502 694894
rect 153586 694658 153822 694894
rect 153266 694338 153502 694574
rect 153586 694338 153822 694574
rect 153266 658658 153502 658894
rect 153586 658658 153822 658894
rect 153266 658338 153502 658574
rect 153586 658338 153822 658574
rect 153266 622658 153502 622894
rect 153586 622658 153822 622894
rect 153266 622338 153502 622574
rect 153586 622338 153822 622574
rect 153266 586658 153502 586894
rect 153586 586658 153822 586894
rect 153266 586338 153502 586574
rect 153586 586338 153822 586574
rect 153266 550658 153502 550894
rect 153586 550658 153822 550894
rect 153266 550338 153502 550574
rect 153586 550338 153822 550574
rect 153266 514658 153502 514894
rect 153586 514658 153822 514894
rect 153266 514338 153502 514574
rect 153586 514338 153822 514574
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 156986 698378 157222 698614
rect 157306 698378 157542 698614
rect 156986 698058 157222 698294
rect 157306 698058 157542 698294
rect 156986 662378 157222 662614
rect 157306 662378 157542 662614
rect 156986 662058 157222 662294
rect 157306 662058 157542 662294
rect 156986 626378 157222 626614
rect 157306 626378 157542 626614
rect 156986 626058 157222 626294
rect 157306 626058 157542 626294
rect 156986 590378 157222 590614
rect 157306 590378 157542 590614
rect 156986 590058 157222 590294
rect 157306 590058 157542 590294
rect 156986 554378 157222 554614
rect 157306 554378 157542 554614
rect 156986 554058 157222 554294
rect 157306 554058 157542 554294
rect 156986 518378 157222 518614
rect 157306 518378 157542 518614
rect 156986 518058 157222 518294
rect 157306 518058 157542 518294
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 163826 669218 164062 669454
rect 164146 669218 164382 669454
rect 163826 668898 164062 669134
rect 164146 668898 164382 669134
rect 163826 633218 164062 633454
rect 164146 633218 164382 633454
rect 163826 632898 164062 633134
rect 164146 632898 164382 633134
rect 163826 597218 164062 597454
rect 164146 597218 164382 597454
rect 163826 596898 164062 597134
rect 164146 596898 164382 597134
rect 163826 561218 164062 561454
rect 164146 561218 164382 561454
rect 163826 560898 164062 561134
rect 164146 560898 164382 561134
rect 163826 525218 164062 525454
rect 164146 525218 164382 525454
rect 163826 524898 164062 525134
rect 164146 524898 164382 525134
rect 163826 489218 164062 489454
rect 164146 489218 164382 489454
rect 163826 488898 164062 489134
rect 164146 488898 164382 489134
rect 167546 672938 167782 673174
rect 167866 672938 168102 673174
rect 167546 672618 167782 672854
rect 167866 672618 168102 672854
rect 167546 636938 167782 637174
rect 167866 636938 168102 637174
rect 167546 636618 167782 636854
rect 167866 636618 168102 636854
rect 167546 600938 167782 601174
rect 167866 600938 168102 601174
rect 167546 600618 167782 600854
rect 167866 600618 168102 600854
rect 167546 564938 167782 565174
rect 167866 564938 168102 565174
rect 167546 564618 167782 564854
rect 167866 564618 168102 564854
rect 167546 528938 167782 529174
rect 167866 528938 168102 529174
rect 167546 528618 167782 528854
rect 167866 528618 168102 528854
rect 167546 492938 167782 493174
rect 167866 492938 168102 493174
rect 167546 492618 167782 492854
rect 167866 492618 168102 492854
rect 171266 676658 171502 676894
rect 171586 676658 171822 676894
rect 171266 676338 171502 676574
rect 171586 676338 171822 676574
rect 171266 640658 171502 640894
rect 171586 640658 171822 640894
rect 171266 640338 171502 640574
rect 171586 640338 171822 640574
rect 171266 604658 171502 604894
rect 171586 604658 171822 604894
rect 171266 604338 171502 604574
rect 171586 604338 171822 604574
rect 171266 568658 171502 568894
rect 171586 568658 171822 568894
rect 171266 568338 171502 568574
rect 171586 568338 171822 568574
rect 171266 532658 171502 532894
rect 171586 532658 171822 532894
rect 171266 532338 171502 532574
rect 171586 532338 171822 532574
rect 171266 496658 171502 496894
rect 171586 496658 171822 496894
rect 171266 496338 171502 496574
rect 171586 496338 171822 496574
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 174986 680378 175222 680614
rect 175306 680378 175542 680614
rect 174986 680058 175222 680294
rect 175306 680058 175542 680294
rect 174986 644378 175222 644614
rect 175306 644378 175542 644614
rect 174986 644058 175222 644294
rect 175306 644058 175542 644294
rect 174986 608378 175222 608614
rect 175306 608378 175542 608614
rect 174986 608058 175222 608294
rect 175306 608058 175542 608294
rect 174986 572378 175222 572614
rect 175306 572378 175542 572614
rect 174986 572058 175222 572294
rect 175306 572058 175542 572294
rect 174986 536378 175222 536614
rect 175306 536378 175542 536614
rect 174986 536058 175222 536294
rect 175306 536058 175542 536294
rect 174986 500378 175222 500614
rect 175306 500378 175542 500614
rect 174986 500058 175222 500294
rect 175306 500058 175542 500294
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 181826 687218 182062 687454
rect 182146 687218 182382 687454
rect 181826 686898 182062 687134
rect 182146 686898 182382 687134
rect 181826 651218 182062 651454
rect 182146 651218 182382 651454
rect 181826 650898 182062 651134
rect 182146 650898 182382 651134
rect 181826 615218 182062 615454
rect 182146 615218 182382 615454
rect 181826 614898 182062 615134
rect 182146 614898 182382 615134
rect 181826 579218 182062 579454
rect 182146 579218 182382 579454
rect 181826 578898 182062 579134
rect 182146 578898 182382 579134
rect 181826 543218 182062 543454
rect 182146 543218 182382 543454
rect 181826 542898 182062 543134
rect 182146 542898 182382 543134
rect 181826 507218 182062 507454
rect 182146 507218 182382 507454
rect 181826 506898 182062 507134
rect 182146 506898 182382 507134
rect 185546 690938 185782 691174
rect 185866 690938 186102 691174
rect 185546 690618 185782 690854
rect 185866 690618 186102 690854
rect 185546 654938 185782 655174
rect 185866 654938 186102 655174
rect 185546 654618 185782 654854
rect 185866 654618 186102 654854
rect 185546 618938 185782 619174
rect 185866 618938 186102 619174
rect 185546 618618 185782 618854
rect 185866 618618 186102 618854
rect 185546 582938 185782 583174
rect 185866 582938 186102 583174
rect 185546 582618 185782 582854
rect 185866 582618 186102 582854
rect 185546 546938 185782 547174
rect 185866 546938 186102 547174
rect 185546 546618 185782 546854
rect 185866 546618 186102 546854
rect 185546 510938 185782 511174
rect 185866 510938 186102 511174
rect 185546 510618 185782 510854
rect 185866 510618 186102 510854
rect 189266 694658 189502 694894
rect 189586 694658 189822 694894
rect 189266 694338 189502 694574
rect 189586 694338 189822 694574
rect 189266 658658 189502 658894
rect 189586 658658 189822 658894
rect 189266 658338 189502 658574
rect 189586 658338 189822 658574
rect 189266 622658 189502 622894
rect 189586 622658 189822 622894
rect 189266 622338 189502 622574
rect 189586 622338 189822 622574
rect 189266 586658 189502 586894
rect 189586 586658 189822 586894
rect 189266 586338 189502 586574
rect 189586 586338 189822 586574
rect 189266 550658 189502 550894
rect 189586 550658 189822 550894
rect 189266 550338 189502 550574
rect 189586 550338 189822 550574
rect 189266 514658 189502 514894
rect 189586 514658 189822 514894
rect 189266 514338 189502 514574
rect 189586 514338 189822 514574
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 192986 698378 193222 698614
rect 193306 698378 193542 698614
rect 192986 698058 193222 698294
rect 193306 698058 193542 698294
rect 192986 662378 193222 662614
rect 193306 662378 193542 662614
rect 192986 662058 193222 662294
rect 193306 662058 193542 662294
rect 192986 626378 193222 626614
rect 193306 626378 193542 626614
rect 192986 626058 193222 626294
rect 193306 626058 193542 626294
rect 192986 590378 193222 590614
rect 193306 590378 193542 590614
rect 192986 590058 193222 590294
rect 193306 590058 193542 590294
rect 192986 554378 193222 554614
rect 193306 554378 193542 554614
rect 192986 554058 193222 554294
rect 193306 554058 193542 554294
rect 192986 518378 193222 518614
rect 193306 518378 193542 518614
rect 192986 518058 193222 518294
rect 193306 518058 193542 518294
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 199826 669218 200062 669454
rect 200146 669218 200382 669454
rect 199826 668898 200062 669134
rect 200146 668898 200382 669134
rect 199826 633218 200062 633454
rect 200146 633218 200382 633454
rect 199826 632898 200062 633134
rect 200146 632898 200382 633134
rect 199826 597218 200062 597454
rect 200146 597218 200382 597454
rect 199826 596898 200062 597134
rect 200146 596898 200382 597134
rect 199826 561218 200062 561454
rect 200146 561218 200382 561454
rect 199826 560898 200062 561134
rect 200146 560898 200382 561134
rect 199826 525218 200062 525454
rect 200146 525218 200382 525454
rect 199826 524898 200062 525134
rect 200146 524898 200382 525134
rect 199826 489218 200062 489454
rect 200146 489218 200382 489454
rect 199826 488898 200062 489134
rect 200146 488898 200382 489134
rect 61008 471218 61244 471454
rect 61008 470898 61244 471134
rect 195376 471218 195612 471454
rect 195376 470898 195612 471134
rect 55826 453218 56062 453454
rect 56146 453218 56382 453454
rect 55826 452898 56062 453134
rect 56146 452898 56382 453134
rect 60328 453218 60564 453454
rect 60328 452898 60564 453134
rect 196056 453218 196292 453454
rect 196056 452898 196292 453134
rect 199826 453218 200062 453454
rect 200146 453218 200382 453454
rect 199826 452898 200062 453134
rect 200146 452898 200382 453134
rect 61008 435218 61244 435454
rect 61008 434898 61244 435134
rect 195376 435218 195612 435454
rect 195376 434898 195612 435134
rect 55826 417218 56062 417454
rect 56146 417218 56382 417454
rect 55826 416898 56062 417134
rect 56146 416898 56382 417134
rect 60328 417218 60564 417454
rect 60328 416898 60564 417134
rect 196056 417218 196292 417454
rect 196056 416898 196292 417134
rect 199826 417218 200062 417454
rect 200146 417218 200382 417454
rect 199826 416898 200062 417134
rect 200146 416898 200382 417134
rect 55826 381218 56062 381454
rect 56146 381218 56382 381454
rect 55826 380898 56062 381134
rect 56146 380898 56382 381134
rect 55826 345218 56062 345454
rect 56146 345218 56382 345454
rect 55826 344898 56062 345134
rect 56146 344898 56382 345134
rect 55826 309218 56062 309454
rect 56146 309218 56382 309454
rect 55826 308898 56062 309134
rect 56146 308898 56382 309134
rect 55826 273218 56062 273454
rect 56146 273218 56382 273454
rect 55826 272898 56062 273134
rect 56146 272898 56382 273134
rect 55826 237218 56062 237454
rect 56146 237218 56382 237454
rect 55826 236898 56062 237134
rect 56146 236898 56382 237134
rect 59546 384938 59782 385174
rect 59866 384938 60102 385174
rect 59546 384618 59782 384854
rect 59866 384618 60102 384854
rect 59546 348938 59782 349174
rect 59866 348938 60102 349174
rect 59546 348618 59782 348854
rect 59866 348618 60102 348854
rect 59546 312938 59782 313174
rect 59866 312938 60102 313174
rect 59546 312618 59782 312854
rect 59866 312618 60102 312854
rect 59546 276938 59782 277174
rect 59866 276938 60102 277174
rect 59546 276618 59782 276854
rect 59866 276618 60102 276854
rect 59546 240938 59782 241174
rect 59866 240938 60102 241174
rect 59546 240618 59782 240854
rect 59866 240618 60102 240854
rect 63266 388658 63502 388894
rect 63586 388658 63822 388894
rect 63266 388338 63502 388574
rect 63586 388338 63822 388574
rect 63266 352658 63502 352894
rect 63586 352658 63822 352894
rect 63266 352338 63502 352574
rect 63586 352338 63822 352574
rect 63266 316658 63502 316894
rect 63586 316658 63822 316894
rect 63266 316338 63502 316574
rect 63586 316338 63822 316574
rect 63266 280658 63502 280894
rect 63586 280658 63822 280894
rect 63266 280338 63502 280574
rect 63586 280338 63822 280574
rect 63266 244658 63502 244894
rect 63586 244658 63822 244894
rect 63266 244338 63502 244574
rect 63586 244338 63822 244574
rect 66986 392378 67222 392614
rect 67306 392378 67542 392614
rect 66986 392058 67222 392294
rect 67306 392058 67542 392294
rect 66986 356378 67222 356614
rect 67306 356378 67542 356614
rect 66986 356058 67222 356294
rect 67306 356058 67542 356294
rect 66986 320378 67222 320614
rect 67306 320378 67542 320614
rect 66986 320058 67222 320294
rect 67306 320058 67542 320294
rect 66986 284378 67222 284614
rect 67306 284378 67542 284614
rect 66986 284058 67222 284294
rect 67306 284058 67542 284294
rect 66986 248378 67222 248614
rect 67306 248378 67542 248614
rect 66986 248058 67222 248294
rect 67306 248058 67542 248294
rect 73826 363218 74062 363454
rect 74146 363218 74382 363454
rect 73826 362898 74062 363134
rect 74146 362898 74382 363134
rect 73826 327218 74062 327454
rect 74146 327218 74382 327454
rect 73826 326898 74062 327134
rect 74146 326898 74382 327134
rect 73826 291218 74062 291454
rect 74146 291218 74382 291454
rect 73826 290898 74062 291134
rect 74146 290898 74382 291134
rect 73826 255218 74062 255454
rect 74146 255218 74382 255454
rect 73826 254898 74062 255134
rect 74146 254898 74382 255134
rect 77546 366938 77782 367174
rect 77866 366938 78102 367174
rect 77546 366618 77782 366854
rect 77866 366618 78102 366854
rect 77546 330938 77782 331174
rect 77866 330938 78102 331174
rect 77546 330618 77782 330854
rect 77866 330618 78102 330854
rect 77546 294938 77782 295174
rect 77866 294938 78102 295174
rect 77546 294618 77782 294854
rect 77866 294618 78102 294854
rect 77546 258938 77782 259174
rect 77866 258938 78102 259174
rect 77546 258618 77782 258854
rect 77866 258618 78102 258854
rect 81266 370658 81502 370894
rect 81586 370658 81822 370894
rect 81266 370338 81502 370574
rect 81586 370338 81822 370574
rect 81266 334658 81502 334894
rect 81586 334658 81822 334894
rect 81266 334338 81502 334574
rect 81586 334338 81822 334574
rect 81266 298658 81502 298894
rect 81586 298658 81822 298894
rect 81266 298338 81502 298574
rect 81586 298338 81822 298574
rect 81266 262658 81502 262894
rect 81586 262658 81822 262894
rect 81266 262338 81502 262574
rect 81586 262338 81822 262574
rect 84986 374378 85222 374614
rect 85306 374378 85542 374614
rect 84986 374058 85222 374294
rect 85306 374058 85542 374294
rect 84986 338378 85222 338614
rect 85306 338378 85542 338614
rect 84986 338058 85222 338294
rect 85306 338058 85542 338294
rect 84986 302378 85222 302614
rect 85306 302378 85542 302614
rect 84986 302058 85222 302294
rect 85306 302058 85542 302294
rect 84986 266378 85222 266614
rect 85306 266378 85542 266614
rect 84986 266058 85222 266294
rect 85306 266058 85542 266294
rect 84986 230378 85222 230614
rect 85306 230378 85542 230614
rect 84986 230058 85222 230294
rect 85306 230058 85542 230294
rect 91826 381218 92062 381454
rect 92146 381218 92382 381454
rect 91826 380898 92062 381134
rect 92146 380898 92382 381134
rect 91826 345218 92062 345454
rect 92146 345218 92382 345454
rect 91826 344898 92062 345134
rect 92146 344898 92382 345134
rect 91826 309218 92062 309454
rect 92146 309218 92382 309454
rect 91826 308898 92062 309134
rect 92146 308898 92382 309134
rect 91826 273218 92062 273454
rect 92146 273218 92382 273454
rect 91826 272898 92062 273134
rect 92146 272898 92382 273134
rect 91826 237218 92062 237454
rect 92146 237218 92382 237454
rect 91826 236898 92062 237134
rect 92146 236898 92382 237134
rect 95546 384938 95782 385174
rect 95866 384938 96102 385174
rect 95546 384618 95782 384854
rect 95866 384618 96102 384854
rect 95546 348938 95782 349174
rect 95866 348938 96102 349174
rect 95546 348618 95782 348854
rect 95866 348618 96102 348854
rect 95546 312938 95782 313174
rect 95866 312938 96102 313174
rect 95546 312618 95782 312854
rect 95866 312618 96102 312854
rect 95546 276938 95782 277174
rect 95866 276938 96102 277174
rect 95546 276618 95782 276854
rect 95866 276618 96102 276854
rect 95546 240938 95782 241174
rect 95866 240938 96102 241174
rect 95546 240618 95782 240854
rect 95866 240618 96102 240854
rect 99266 388658 99502 388894
rect 99586 388658 99822 388894
rect 99266 388338 99502 388574
rect 99586 388338 99822 388574
rect 99266 352658 99502 352894
rect 99586 352658 99822 352894
rect 99266 352338 99502 352574
rect 99586 352338 99822 352574
rect 99266 316658 99502 316894
rect 99586 316658 99822 316894
rect 99266 316338 99502 316574
rect 99586 316338 99822 316574
rect 99266 280658 99502 280894
rect 99586 280658 99822 280894
rect 99266 280338 99502 280574
rect 99586 280338 99822 280574
rect 99266 244658 99502 244894
rect 99586 244658 99822 244894
rect 99266 244338 99502 244574
rect 99586 244338 99822 244574
rect 102986 392378 103222 392614
rect 103306 392378 103542 392614
rect 102986 392058 103222 392294
rect 103306 392058 103542 392294
rect 102986 356378 103222 356614
rect 103306 356378 103542 356614
rect 102986 356058 103222 356294
rect 103306 356058 103542 356294
rect 102986 320378 103222 320614
rect 103306 320378 103542 320614
rect 102986 320058 103222 320294
rect 103306 320058 103542 320294
rect 102986 284378 103222 284614
rect 103306 284378 103542 284614
rect 102986 284058 103222 284294
rect 103306 284058 103542 284294
rect 102986 248378 103222 248614
rect 103306 248378 103542 248614
rect 102986 248058 103222 248294
rect 103306 248058 103542 248294
rect 109826 363218 110062 363454
rect 110146 363218 110382 363454
rect 109826 362898 110062 363134
rect 110146 362898 110382 363134
rect 109826 327218 110062 327454
rect 110146 327218 110382 327454
rect 109826 326898 110062 327134
rect 110146 326898 110382 327134
rect 109826 291218 110062 291454
rect 110146 291218 110382 291454
rect 109826 290898 110062 291134
rect 110146 290898 110382 291134
rect 109826 255218 110062 255454
rect 110146 255218 110382 255454
rect 109826 254898 110062 255134
rect 110146 254898 110382 255134
rect 113546 366938 113782 367174
rect 113866 366938 114102 367174
rect 113546 366618 113782 366854
rect 113866 366618 114102 366854
rect 113546 330938 113782 331174
rect 113866 330938 114102 331174
rect 113546 330618 113782 330854
rect 113866 330618 114102 330854
rect 113546 294938 113782 295174
rect 113866 294938 114102 295174
rect 113546 294618 113782 294854
rect 113866 294618 114102 294854
rect 113546 258938 113782 259174
rect 113866 258938 114102 259174
rect 113546 258618 113782 258854
rect 113866 258618 114102 258854
rect 117266 370658 117502 370894
rect 117586 370658 117822 370894
rect 117266 370338 117502 370574
rect 117586 370338 117822 370574
rect 117266 334658 117502 334894
rect 117586 334658 117822 334894
rect 117266 334338 117502 334574
rect 117586 334338 117822 334574
rect 117266 298658 117502 298894
rect 117586 298658 117822 298894
rect 117266 298338 117502 298574
rect 117586 298338 117822 298574
rect 117266 262658 117502 262894
rect 117586 262658 117822 262894
rect 117266 262338 117502 262574
rect 117586 262338 117822 262574
rect 120986 374378 121222 374614
rect 121306 374378 121542 374614
rect 120986 374058 121222 374294
rect 121306 374058 121542 374294
rect 120986 338378 121222 338614
rect 121306 338378 121542 338614
rect 120986 338058 121222 338294
rect 121306 338058 121542 338294
rect 120986 302378 121222 302614
rect 121306 302378 121542 302614
rect 120986 302058 121222 302294
rect 121306 302058 121542 302294
rect 120986 266378 121222 266614
rect 121306 266378 121542 266614
rect 120986 266058 121222 266294
rect 121306 266058 121542 266294
rect 120986 230378 121222 230614
rect 121306 230378 121542 230614
rect 120986 230058 121222 230294
rect 121306 230058 121542 230294
rect 127826 381218 128062 381454
rect 128146 381218 128382 381454
rect 127826 380898 128062 381134
rect 128146 380898 128382 381134
rect 127826 345218 128062 345454
rect 128146 345218 128382 345454
rect 127826 344898 128062 345134
rect 128146 344898 128382 345134
rect 127826 309218 128062 309454
rect 128146 309218 128382 309454
rect 127826 308898 128062 309134
rect 128146 308898 128382 309134
rect 127826 273218 128062 273454
rect 128146 273218 128382 273454
rect 127826 272898 128062 273134
rect 128146 272898 128382 273134
rect 127826 237218 128062 237454
rect 128146 237218 128382 237454
rect 127826 236898 128062 237134
rect 128146 236898 128382 237134
rect 131546 384938 131782 385174
rect 131866 384938 132102 385174
rect 131546 384618 131782 384854
rect 131866 384618 132102 384854
rect 131546 348938 131782 349174
rect 131866 348938 132102 349174
rect 131546 348618 131782 348854
rect 131866 348618 132102 348854
rect 131546 312938 131782 313174
rect 131866 312938 132102 313174
rect 131546 312618 131782 312854
rect 131866 312618 132102 312854
rect 131546 276938 131782 277174
rect 131866 276938 132102 277174
rect 131546 276618 131782 276854
rect 131866 276618 132102 276854
rect 131546 240938 131782 241174
rect 131866 240938 132102 241174
rect 131546 240618 131782 240854
rect 131866 240618 132102 240854
rect 135266 388658 135502 388894
rect 135586 388658 135822 388894
rect 135266 388338 135502 388574
rect 135586 388338 135822 388574
rect 135266 352658 135502 352894
rect 135586 352658 135822 352894
rect 135266 352338 135502 352574
rect 135586 352338 135822 352574
rect 135266 316658 135502 316894
rect 135586 316658 135822 316894
rect 135266 316338 135502 316574
rect 135586 316338 135822 316574
rect 135266 280658 135502 280894
rect 135586 280658 135822 280894
rect 135266 280338 135502 280574
rect 135586 280338 135822 280574
rect 135266 244658 135502 244894
rect 135586 244658 135822 244894
rect 135266 244338 135502 244574
rect 135586 244338 135822 244574
rect 138986 392378 139222 392614
rect 139306 392378 139542 392614
rect 138986 392058 139222 392294
rect 139306 392058 139542 392294
rect 138986 356378 139222 356614
rect 139306 356378 139542 356614
rect 138986 356058 139222 356294
rect 139306 356058 139542 356294
rect 138986 320378 139222 320614
rect 139306 320378 139542 320614
rect 138986 320058 139222 320294
rect 139306 320058 139542 320294
rect 138986 284378 139222 284614
rect 139306 284378 139542 284614
rect 138986 284058 139222 284294
rect 139306 284058 139542 284294
rect 138986 248378 139222 248614
rect 139306 248378 139542 248614
rect 138986 248058 139222 248294
rect 139306 248058 139542 248294
rect 145826 363218 146062 363454
rect 146146 363218 146382 363454
rect 145826 362898 146062 363134
rect 146146 362898 146382 363134
rect 145826 327218 146062 327454
rect 146146 327218 146382 327454
rect 145826 326898 146062 327134
rect 146146 326898 146382 327134
rect 145826 291218 146062 291454
rect 146146 291218 146382 291454
rect 145826 290898 146062 291134
rect 146146 290898 146382 291134
rect 145826 255218 146062 255454
rect 146146 255218 146382 255454
rect 145826 254898 146062 255134
rect 146146 254898 146382 255134
rect 149546 366938 149782 367174
rect 149866 366938 150102 367174
rect 149546 366618 149782 366854
rect 149866 366618 150102 366854
rect 149546 330938 149782 331174
rect 149866 330938 150102 331174
rect 149546 330618 149782 330854
rect 149866 330618 150102 330854
rect 149546 294938 149782 295174
rect 149866 294938 150102 295174
rect 149546 294618 149782 294854
rect 149866 294618 150102 294854
rect 149546 258938 149782 259174
rect 149866 258938 150102 259174
rect 149546 258618 149782 258854
rect 149866 258618 150102 258854
rect 153266 370658 153502 370894
rect 153586 370658 153822 370894
rect 153266 370338 153502 370574
rect 153586 370338 153822 370574
rect 153266 334658 153502 334894
rect 153586 334658 153822 334894
rect 153266 334338 153502 334574
rect 153586 334338 153822 334574
rect 153266 298658 153502 298894
rect 153586 298658 153822 298894
rect 153266 298338 153502 298574
rect 153586 298338 153822 298574
rect 153266 262658 153502 262894
rect 153586 262658 153822 262894
rect 153266 262338 153502 262574
rect 153586 262338 153822 262574
rect 156986 374378 157222 374614
rect 157306 374378 157542 374614
rect 156986 374058 157222 374294
rect 157306 374058 157542 374294
rect 156986 338378 157222 338614
rect 157306 338378 157542 338614
rect 156986 338058 157222 338294
rect 157306 338058 157542 338294
rect 156986 302378 157222 302614
rect 157306 302378 157542 302614
rect 156986 302058 157222 302294
rect 157306 302058 157542 302294
rect 156986 266378 157222 266614
rect 157306 266378 157542 266614
rect 156986 266058 157222 266294
rect 157306 266058 157542 266294
rect 156986 230378 157222 230614
rect 157306 230378 157542 230614
rect 156986 230058 157222 230294
rect 157306 230058 157542 230294
rect 163826 381218 164062 381454
rect 164146 381218 164382 381454
rect 163826 380898 164062 381134
rect 164146 380898 164382 381134
rect 163826 345218 164062 345454
rect 164146 345218 164382 345454
rect 163826 344898 164062 345134
rect 164146 344898 164382 345134
rect 163826 309218 164062 309454
rect 164146 309218 164382 309454
rect 163826 308898 164062 309134
rect 164146 308898 164382 309134
rect 163826 273218 164062 273454
rect 164146 273218 164382 273454
rect 163826 272898 164062 273134
rect 164146 272898 164382 273134
rect 163826 237218 164062 237454
rect 164146 237218 164382 237454
rect 163826 236898 164062 237134
rect 164146 236898 164382 237134
rect 167546 384938 167782 385174
rect 167866 384938 168102 385174
rect 167546 384618 167782 384854
rect 167866 384618 168102 384854
rect 167546 348938 167782 349174
rect 167866 348938 168102 349174
rect 167546 348618 167782 348854
rect 167866 348618 168102 348854
rect 167546 312938 167782 313174
rect 167866 312938 168102 313174
rect 167546 312618 167782 312854
rect 167866 312618 168102 312854
rect 167546 276938 167782 277174
rect 167866 276938 168102 277174
rect 167546 276618 167782 276854
rect 167866 276618 168102 276854
rect 167546 240938 167782 241174
rect 167866 240938 168102 241174
rect 167546 240618 167782 240854
rect 167866 240618 168102 240854
rect 171266 388658 171502 388894
rect 171586 388658 171822 388894
rect 171266 388338 171502 388574
rect 171586 388338 171822 388574
rect 171266 352658 171502 352894
rect 171586 352658 171822 352894
rect 171266 352338 171502 352574
rect 171586 352338 171822 352574
rect 171266 316658 171502 316894
rect 171586 316658 171822 316894
rect 171266 316338 171502 316574
rect 171586 316338 171822 316574
rect 171266 280658 171502 280894
rect 171586 280658 171822 280894
rect 171266 280338 171502 280574
rect 171586 280338 171822 280574
rect 171266 244658 171502 244894
rect 171586 244658 171822 244894
rect 171266 244338 171502 244574
rect 171586 244338 171822 244574
rect 174986 392378 175222 392614
rect 175306 392378 175542 392614
rect 174986 392058 175222 392294
rect 175306 392058 175542 392294
rect 174986 356378 175222 356614
rect 175306 356378 175542 356614
rect 174986 356058 175222 356294
rect 175306 356058 175542 356294
rect 174986 320378 175222 320614
rect 175306 320378 175542 320614
rect 174986 320058 175222 320294
rect 175306 320058 175542 320294
rect 174986 284378 175222 284614
rect 175306 284378 175542 284614
rect 174986 284058 175222 284294
rect 175306 284058 175542 284294
rect 174986 248378 175222 248614
rect 175306 248378 175542 248614
rect 174986 248058 175222 248294
rect 175306 248058 175542 248294
rect 181826 363218 182062 363454
rect 182146 363218 182382 363454
rect 181826 362898 182062 363134
rect 182146 362898 182382 363134
rect 181826 327218 182062 327454
rect 182146 327218 182382 327454
rect 181826 326898 182062 327134
rect 182146 326898 182382 327134
rect 181826 291218 182062 291454
rect 182146 291218 182382 291454
rect 181826 290898 182062 291134
rect 182146 290898 182382 291134
rect 181826 255218 182062 255454
rect 182146 255218 182382 255454
rect 181826 254898 182062 255134
rect 182146 254898 182382 255134
rect 185546 366938 185782 367174
rect 185866 366938 186102 367174
rect 185546 366618 185782 366854
rect 185866 366618 186102 366854
rect 185546 330938 185782 331174
rect 185866 330938 186102 331174
rect 185546 330618 185782 330854
rect 185866 330618 186102 330854
rect 185546 294938 185782 295174
rect 185866 294938 186102 295174
rect 185546 294618 185782 294854
rect 185866 294618 186102 294854
rect 185546 258938 185782 259174
rect 185866 258938 186102 259174
rect 185546 258618 185782 258854
rect 185866 258618 186102 258854
rect 189266 370658 189502 370894
rect 189586 370658 189822 370894
rect 189266 370338 189502 370574
rect 189586 370338 189822 370574
rect 189266 334658 189502 334894
rect 189586 334658 189822 334894
rect 189266 334338 189502 334574
rect 189586 334338 189822 334574
rect 189266 298658 189502 298894
rect 189586 298658 189822 298894
rect 189266 298338 189502 298574
rect 189586 298338 189822 298574
rect 189266 262658 189502 262894
rect 189586 262658 189822 262894
rect 189266 262338 189502 262574
rect 189586 262338 189822 262574
rect 192986 374378 193222 374614
rect 193306 374378 193542 374614
rect 192986 374058 193222 374294
rect 193306 374058 193542 374294
rect 192986 338378 193222 338614
rect 193306 338378 193542 338614
rect 192986 338058 193222 338294
rect 193306 338058 193542 338294
rect 192986 302378 193222 302614
rect 193306 302378 193542 302614
rect 192986 302058 193222 302294
rect 193306 302058 193542 302294
rect 192986 266378 193222 266614
rect 193306 266378 193542 266614
rect 192986 266058 193222 266294
rect 193306 266058 193542 266294
rect 192986 230378 193222 230614
rect 193306 230378 193542 230614
rect 192986 230058 193222 230294
rect 193306 230058 193542 230294
rect 199826 381218 200062 381454
rect 200146 381218 200382 381454
rect 199826 380898 200062 381134
rect 200146 380898 200382 381134
rect 199826 345218 200062 345454
rect 200146 345218 200382 345454
rect 199826 344898 200062 345134
rect 200146 344898 200382 345134
rect 199826 309218 200062 309454
rect 200146 309218 200382 309454
rect 199826 308898 200062 309134
rect 200146 308898 200382 309134
rect 199826 273218 200062 273454
rect 200146 273218 200382 273454
rect 199826 272898 200062 273134
rect 200146 272898 200382 273134
rect 199826 237218 200062 237454
rect 200146 237218 200382 237454
rect 199826 236898 200062 237134
rect 200146 236898 200382 237134
rect 203546 672938 203782 673174
rect 203866 672938 204102 673174
rect 203546 672618 203782 672854
rect 203866 672618 204102 672854
rect 203546 636938 203782 637174
rect 203866 636938 204102 637174
rect 203546 636618 203782 636854
rect 203866 636618 204102 636854
rect 203546 600938 203782 601174
rect 203866 600938 204102 601174
rect 203546 600618 203782 600854
rect 203866 600618 204102 600854
rect 203546 564938 203782 565174
rect 203866 564938 204102 565174
rect 203546 564618 203782 564854
rect 203866 564618 204102 564854
rect 203546 528938 203782 529174
rect 203866 528938 204102 529174
rect 203546 528618 203782 528854
rect 203866 528618 204102 528854
rect 203546 492938 203782 493174
rect 203866 492938 204102 493174
rect 203546 492618 203782 492854
rect 203866 492618 204102 492854
rect 203546 456938 203782 457174
rect 203866 456938 204102 457174
rect 203546 456618 203782 456854
rect 203866 456618 204102 456854
rect 203546 420938 203782 421174
rect 203866 420938 204102 421174
rect 203546 420618 203782 420854
rect 203866 420618 204102 420854
rect 203546 384938 203782 385174
rect 203866 384938 204102 385174
rect 203546 384618 203782 384854
rect 203866 384618 204102 384854
rect 203546 348938 203782 349174
rect 203866 348938 204102 349174
rect 203546 348618 203782 348854
rect 203866 348618 204102 348854
rect 203546 312938 203782 313174
rect 203866 312938 204102 313174
rect 203546 312618 203782 312854
rect 203866 312618 204102 312854
rect 203546 276938 203782 277174
rect 203866 276938 204102 277174
rect 203546 276618 203782 276854
rect 203866 276618 204102 276854
rect 203546 240938 203782 241174
rect 203866 240938 204102 241174
rect 203546 240618 203782 240854
rect 203866 240618 204102 240854
rect 207266 676658 207502 676894
rect 207586 676658 207822 676894
rect 207266 676338 207502 676574
rect 207586 676338 207822 676574
rect 207266 640658 207502 640894
rect 207586 640658 207822 640894
rect 207266 640338 207502 640574
rect 207586 640338 207822 640574
rect 207266 604658 207502 604894
rect 207586 604658 207822 604894
rect 207266 604338 207502 604574
rect 207586 604338 207822 604574
rect 207266 568658 207502 568894
rect 207586 568658 207822 568894
rect 207266 568338 207502 568574
rect 207586 568338 207822 568574
rect 207266 532658 207502 532894
rect 207586 532658 207822 532894
rect 207266 532338 207502 532574
rect 207586 532338 207822 532574
rect 207266 496658 207502 496894
rect 207586 496658 207822 496894
rect 207266 496338 207502 496574
rect 207586 496338 207822 496574
rect 207266 460658 207502 460894
rect 207586 460658 207822 460894
rect 207266 460338 207502 460574
rect 207586 460338 207822 460574
rect 207266 424658 207502 424894
rect 207586 424658 207822 424894
rect 207266 424338 207502 424574
rect 207586 424338 207822 424574
rect 207266 388658 207502 388894
rect 207586 388658 207822 388894
rect 207266 388338 207502 388574
rect 207586 388338 207822 388574
rect 207266 352658 207502 352894
rect 207586 352658 207822 352894
rect 207266 352338 207502 352574
rect 207586 352338 207822 352574
rect 207266 316658 207502 316894
rect 207586 316658 207822 316894
rect 207266 316338 207502 316574
rect 207586 316338 207822 316574
rect 207266 280658 207502 280894
rect 207586 280658 207822 280894
rect 207266 280338 207502 280574
rect 207586 280338 207822 280574
rect 207266 244658 207502 244894
rect 207586 244658 207822 244894
rect 207266 244338 207502 244574
rect 207586 244338 207822 244574
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 210986 680378 211222 680614
rect 211306 680378 211542 680614
rect 210986 680058 211222 680294
rect 211306 680058 211542 680294
rect 210986 644378 211222 644614
rect 211306 644378 211542 644614
rect 210986 644058 211222 644294
rect 211306 644058 211542 644294
rect 210986 608378 211222 608614
rect 211306 608378 211542 608614
rect 210986 608058 211222 608294
rect 211306 608058 211542 608294
rect 210986 572378 211222 572614
rect 211306 572378 211542 572614
rect 210986 572058 211222 572294
rect 211306 572058 211542 572294
rect 210986 536378 211222 536614
rect 211306 536378 211542 536614
rect 210986 536058 211222 536294
rect 211306 536058 211542 536294
rect 210986 500378 211222 500614
rect 211306 500378 211542 500614
rect 210986 500058 211222 500294
rect 211306 500058 211542 500294
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 217826 687218 218062 687454
rect 218146 687218 218382 687454
rect 217826 686898 218062 687134
rect 218146 686898 218382 687134
rect 217826 651218 218062 651454
rect 218146 651218 218382 651454
rect 217826 650898 218062 651134
rect 218146 650898 218382 651134
rect 217826 615218 218062 615454
rect 218146 615218 218382 615454
rect 217826 614898 218062 615134
rect 218146 614898 218382 615134
rect 217826 579218 218062 579454
rect 218146 579218 218382 579454
rect 217826 578898 218062 579134
rect 218146 578898 218382 579134
rect 217826 543218 218062 543454
rect 218146 543218 218382 543454
rect 217826 542898 218062 543134
rect 218146 542898 218382 543134
rect 217826 507218 218062 507454
rect 218146 507218 218382 507454
rect 217826 506898 218062 507134
rect 218146 506898 218382 507134
rect 221546 690938 221782 691174
rect 221866 690938 222102 691174
rect 221546 690618 221782 690854
rect 221866 690618 222102 690854
rect 221546 654938 221782 655174
rect 221866 654938 222102 655174
rect 221546 654618 221782 654854
rect 221866 654618 222102 654854
rect 221546 618938 221782 619174
rect 221866 618938 222102 619174
rect 221546 618618 221782 618854
rect 221866 618618 222102 618854
rect 221546 582938 221782 583174
rect 221866 582938 222102 583174
rect 221546 582618 221782 582854
rect 221866 582618 222102 582854
rect 221546 546938 221782 547174
rect 221866 546938 222102 547174
rect 221546 546618 221782 546854
rect 221866 546618 222102 546854
rect 221546 510938 221782 511174
rect 221866 510938 222102 511174
rect 221546 510618 221782 510854
rect 221866 510618 222102 510854
rect 210986 464378 211222 464614
rect 211306 464378 211542 464614
rect 210986 464058 211222 464294
rect 211306 464058 211542 464294
rect 210986 428378 211222 428614
rect 211306 428378 211542 428614
rect 210986 428058 211222 428294
rect 211306 428058 211542 428294
rect 210986 392378 211222 392614
rect 211306 392378 211542 392614
rect 210986 392058 211222 392294
rect 211306 392058 211542 392294
rect 210986 356378 211222 356614
rect 211306 356378 211542 356614
rect 210986 356058 211222 356294
rect 211306 356058 211542 356294
rect 210986 320378 211222 320614
rect 211306 320378 211542 320614
rect 210986 320058 211222 320294
rect 211306 320058 211542 320294
rect 210986 284378 211222 284614
rect 211306 284378 211542 284614
rect 210986 284058 211222 284294
rect 211306 284058 211542 284294
rect 210986 248378 211222 248614
rect 211306 248378 211542 248614
rect 210986 248058 211222 248294
rect 211306 248058 211542 248294
rect 217826 363218 218062 363454
rect 218146 363218 218382 363454
rect 217826 362898 218062 363134
rect 218146 362898 218382 363134
rect 217826 327218 218062 327454
rect 218146 327218 218382 327454
rect 217826 326898 218062 327134
rect 218146 326898 218382 327134
rect 217826 291218 218062 291454
rect 218146 291218 218382 291454
rect 217826 290898 218062 291134
rect 218146 290898 218382 291134
rect 217826 255218 218062 255454
rect 218146 255218 218382 255454
rect 217826 254898 218062 255134
rect 218146 254898 218382 255134
rect 225266 694658 225502 694894
rect 225586 694658 225822 694894
rect 225266 694338 225502 694574
rect 225586 694338 225822 694574
rect 225266 658658 225502 658894
rect 225586 658658 225822 658894
rect 225266 658338 225502 658574
rect 225586 658338 225822 658574
rect 225266 622658 225502 622894
rect 225586 622658 225822 622894
rect 225266 622338 225502 622574
rect 225586 622338 225822 622574
rect 225266 586658 225502 586894
rect 225586 586658 225822 586894
rect 225266 586338 225502 586574
rect 225586 586338 225822 586574
rect 225266 550658 225502 550894
rect 225586 550658 225822 550894
rect 225266 550338 225502 550574
rect 225586 550338 225822 550574
rect 225266 514658 225502 514894
rect 225586 514658 225822 514894
rect 225266 514338 225502 514574
rect 225586 514338 225822 514574
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 228986 698378 229222 698614
rect 229306 698378 229542 698614
rect 228986 698058 229222 698294
rect 229306 698058 229542 698294
rect 228986 662378 229222 662614
rect 229306 662378 229542 662614
rect 228986 662058 229222 662294
rect 229306 662058 229542 662294
rect 228986 626378 229222 626614
rect 229306 626378 229542 626614
rect 228986 626058 229222 626294
rect 229306 626058 229542 626294
rect 228986 590378 229222 590614
rect 229306 590378 229542 590614
rect 228986 590058 229222 590294
rect 229306 590058 229542 590294
rect 228986 554378 229222 554614
rect 229306 554378 229542 554614
rect 228986 554058 229222 554294
rect 229306 554058 229542 554294
rect 228986 518378 229222 518614
rect 229306 518378 229542 518614
rect 228986 518058 229222 518294
rect 229306 518058 229542 518294
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 235826 669218 236062 669454
rect 236146 669218 236382 669454
rect 235826 668898 236062 669134
rect 236146 668898 236382 669134
rect 235826 633218 236062 633454
rect 236146 633218 236382 633454
rect 235826 632898 236062 633134
rect 236146 632898 236382 633134
rect 235826 597218 236062 597454
rect 236146 597218 236382 597454
rect 235826 596898 236062 597134
rect 236146 596898 236382 597134
rect 235826 561218 236062 561454
rect 236146 561218 236382 561454
rect 235826 560898 236062 561134
rect 236146 560898 236382 561134
rect 235826 525218 236062 525454
rect 236146 525218 236382 525454
rect 235826 524898 236062 525134
rect 236146 524898 236382 525134
rect 235826 489218 236062 489454
rect 236146 489218 236382 489454
rect 235826 488898 236062 489134
rect 236146 488898 236382 489134
rect 239546 672938 239782 673174
rect 239866 672938 240102 673174
rect 239546 672618 239782 672854
rect 239866 672618 240102 672854
rect 239546 636938 239782 637174
rect 239866 636938 240102 637174
rect 239546 636618 239782 636854
rect 239866 636618 240102 636854
rect 239546 600938 239782 601174
rect 239866 600938 240102 601174
rect 239546 600618 239782 600854
rect 239866 600618 240102 600854
rect 239546 564938 239782 565174
rect 239866 564938 240102 565174
rect 239546 564618 239782 564854
rect 239866 564618 240102 564854
rect 239546 528938 239782 529174
rect 239866 528938 240102 529174
rect 239546 528618 239782 528854
rect 239866 528618 240102 528854
rect 239546 492938 239782 493174
rect 239866 492938 240102 493174
rect 239546 492618 239782 492854
rect 239866 492618 240102 492854
rect 243266 676658 243502 676894
rect 243586 676658 243822 676894
rect 243266 676338 243502 676574
rect 243586 676338 243822 676574
rect 243266 640658 243502 640894
rect 243586 640658 243822 640894
rect 243266 640338 243502 640574
rect 243586 640338 243822 640574
rect 243266 604658 243502 604894
rect 243586 604658 243822 604894
rect 243266 604338 243502 604574
rect 243586 604338 243822 604574
rect 243266 568658 243502 568894
rect 243586 568658 243822 568894
rect 243266 568338 243502 568574
rect 243586 568338 243822 568574
rect 243266 532658 243502 532894
rect 243586 532658 243822 532894
rect 243266 532338 243502 532574
rect 243586 532338 243822 532574
rect 243266 496658 243502 496894
rect 243586 496658 243822 496894
rect 243266 496338 243502 496574
rect 243586 496338 243822 496574
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 246986 680378 247222 680614
rect 247306 680378 247542 680614
rect 246986 680058 247222 680294
rect 247306 680058 247542 680294
rect 246986 644378 247222 644614
rect 247306 644378 247542 644614
rect 246986 644058 247222 644294
rect 247306 644058 247542 644294
rect 246986 608378 247222 608614
rect 247306 608378 247542 608614
rect 246986 608058 247222 608294
rect 247306 608058 247542 608294
rect 246986 572378 247222 572614
rect 247306 572378 247542 572614
rect 246986 572058 247222 572294
rect 247306 572058 247542 572294
rect 246986 536378 247222 536614
rect 247306 536378 247542 536614
rect 246986 536058 247222 536294
rect 247306 536058 247542 536294
rect 246986 500378 247222 500614
rect 247306 500378 247542 500614
rect 246986 500058 247222 500294
rect 247306 500058 247542 500294
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 253826 687218 254062 687454
rect 254146 687218 254382 687454
rect 253826 686898 254062 687134
rect 254146 686898 254382 687134
rect 253826 651218 254062 651454
rect 254146 651218 254382 651454
rect 253826 650898 254062 651134
rect 254146 650898 254382 651134
rect 253826 615218 254062 615454
rect 254146 615218 254382 615454
rect 253826 614898 254062 615134
rect 254146 614898 254382 615134
rect 253826 579218 254062 579454
rect 254146 579218 254382 579454
rect 253826 578898 254062 579134
rect 254146 578898 254382 579134
rect 253826 543218 254062 543454
rect 254146 543218 254382 543454
rect 253826 542898 254062 543134
rect 254146 542898 254382 543134
rect 253826 507218 254062 507454
rect 254146 507218 254382 507454
rect 253826 506898 254062 507134
rect 254146 506898 254382 507134
rect 257546 690938 257782 691174
rect 257866 690938 258102 691174
rect 257546 690618 257782 690854
rect 257866 690618 258102 690854
rect 257546 654938 257782 655174
rect 257866 654938 258102 655174
rect 257546 654618 257782 654854
rect 257866 654618 258102 654854
rect 257546 618938 257782 619174
rect 257866 618938 258102 619174
rect 257546 618618 257782 618854
rect 257866 618618 258102 618854
rect 257546 582938 257782 583174
rect 257866 582938 258102 583174
rect 257546 582618 257782 582854
rect 257866 582618 258102 582854
rect 257546 546938 257782 547174
rect 257866 546938 258102 547174
rect 257546 546618 257782 546854
rect 257866 546618 258102 546854
rect 257546 510938 257782 511174
rect 257866 510938 258102 511174
rect 257546 510618 257782 510854
rect 257866 510618 258102 510854
rect 261266 694658 261502 694894
rect 261586 694658 261822 694894
rect 261266 694338 261502 694574
rect 261586 694338 261822 694574
rect 261266 658658 261502 658894
rect 261586 658658 261822 658894
rect 261266 658338 261502 658574
rect 261586 658338 261822 658574
rect 261266 622658 261502 622894
rect 261586 622658 261822 622894
rect 261266 622338 261502 622574
rect 261586 622338 261822 622574
rect 261266 586658 261502 586894
rect 261586 586658 261822 586894
rect 261266 586338 261502 586574
rect 261586 586338 261822 586574
rect 261266 550658 261502 550894
rect 261586 550658 261822 550894
rect 261266 550338 261502 550574
rect 261586 550338 261822 550574
rect 261266 514658 261502 514894
rect 261586 514658 261822 514894
rect 261266 514338 261502 514574
rect 261586 514338 261822 514574
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 264986 698378 265222 698614
rect 265306 698378 265542 698614
rect 264986 698058 265222 698294
rect 265306 698058 265542 698294
rect 264986 662378 265222 662614
rect 265306 662378 265542 662614
rect 264986 662058 265222 662294
rect 265306 662058 265542 662294
rect 264986 626378 265222 626614
rect 265306 626378 265542 626614
rect 264986 626058 265222 626294
rect 265306 626058 265542 626294
rect 264986 590378 265222 590614
rect 265306 590378 265542 590614
rect 264986 590058 265222 590294
rect 265306 590058 265542 590294
rect 264986 554378 265222 554614
rect 265306 554378 265542 554614
rect 264986 554058 265222 554294
rect 265306 554058 265542 554294
rect 264986 518378 265222 518614
rect 265306 518378 265542 518614
rect 264986 518058 265222 518294
rect 265306 518058 265542 518294
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 271826 669218 272062 669454
rect 272146 669218 272382 669454
rect 271826 668898 272062 669134
rect 272146 668898 272382 669134
rect 271826 633218 272062 633454
rect 272146 633218 272382 633454
rect 271826 632898 272062 633134
rect 272146 632898 272382 633134
rect 271826 597218 272062 597454
rect 272146 597218 272382 597454
rect 271826 596898 272062 597134
rect 272146 596898 272382 597134
rect 271826 561218 272062 561454
rect 272146 561218 272382 561454
rect 271826 560898 272062 561134
rect 272146 560898 272382 561134
rect 271826 525218 272062 525454
rect 272146 525218 272382 525454
rect 271826 524898 272062 525134
rect 272146 524898 272382 525134
rect 271826 489218 272062 489454
rect 272146 489218 272382 489454
rect 271826 488898 272062 489134
rect 272146 488898 272382 489134
rect 275546 672938 275782 673174
rect 275866 672938 276102 673174
rect 275546 672618 275782 672854
rect 275866 672618 276102 672854
rect 275546 636938 275782 637174
rect 275866 636938 276102 637174
rect 275546 636618 275782 636854
rect 275866 636618 276102 636854
rect 275546 600938 275782 601174
rect 275866 600938 276102 601174
rect 275546 600618 275782 600854
rect 275866 600618 276102 600854
rect 275546 564938 275782 565174
rect 275866 564938 276102 565174
rect 275546 564618 275782 564854
rect 275866 564618 276102 564854
rect 275546 528938 275782 529174
rect 275866 528938 276102 529174
rect 275546 528618 275782 528854
rect 275866 528618 276102 528854
rect 275546 492938 275782 493174
rect 275866 492938 276102 493174
rect 275546 492618 275782 492854
rect 275866 492618 276102 492854
rect 279266 676658 279502 676894
rect 279586 676658 279822 676894
rect 279266 676338 279502 676574
rect 279586 676338 279822 676574
rect 279266 640658 279502 640894
rect 279586 640658 279822 640894
rect 279266 640338 279502 640574
rect 279586 640338 279822 640574
rect 279266 604658 279502 604894
rect 279586 604658 279822 604894
rect 279266 604338 279502 604574
rect 279586 604338 279822 604574
rect 279266 568658 279502 568894
rect 279586 568658 279822 568894
rect 279266 568338 279502 568574
rect 279586 568338 279822 568574
rect 279266 532658 279502 532894
rect 279586 532658 279822 532894
rect 279266 532338 279502 532574
rect 279586 532338 279822 532574
rect 279266 496658 279502 496894
rect 279586 496658 279822 496894
rect 279266 496338 279502 496574
rect 279586 496338 279822 496574
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 282986 680378 283222 680614
rect 283306 680378 283542 680614
rect 282986 680058 283222 680294
rect 283306 680058 283542 680294
rect 282986 644378 283222 644614
rect 283306 644378 283542 644614
rect 282986 644058 283222 644294
rect 283306 644058 283542 644294
rect 282986 608378 283222 608614
rect 283306 608378 283542 608614
rect 282986 608058 283222 608294
rect 283306 608058 283542 608294
rect 282986 572378 283222 572614
rect 283306 572378 283542 572614
rect 282986 572058 283222 572294
rect 283306 572058 283542 572294
rect 282986 536378 283222 536614
rect 283306 536378 283542 536614
rect 282986 536058 283222 536294
rect 283306 536058 283542 536294
rect 282986 500378 283222 500614
rect 283306 500378 283542 500614
rect 282986 500058 283222 500294
rect 283306 500058 283542 500294
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 289826 687218 290062 687454
rect 290146 687218 290382 687454
rect 289826 686898 290062 687134
rect 290146 686898 290382 687134
rect 289826 651218 290062 651454
rect 290146 651218 290382 651454
rect 289826 650898 290062 651134
rect 290146 650898 290382 651134
rect 289826 615218 290062 615454
rect 290146 615218 290382 615454
rect 289826 614898 290062 615134
rect 290146 614898 290382 615134
rect 289826 579218 290062 579454
rect 290146 579218 290382 579454
rect 289826 578898 290062 579134
rect 290146 578898 290382 579134
rect 289826 543218 290062 543454
rect 290146 543218 290382 543454
rect 289826 542898 290062 543134
rect 290146 542898 290382 543134
rect 289826 507218 290062 507454
rect 290146 507218 290382 507454
rect 289826 506898 290062 507134
rect 290146 506898 290382 507134
rect 293546 690938 293782 691174
rect 293866 690938 294102 691174
rect 293546 690618 293782 690854
rect 293866 690618 294102 690854
rect 293546 654938 293782 655174
rect 293866 654938 294102 655174
rect 293546 654618 293782 654854
rect 293866 654618 294102 654854
rect 293546 618938 293782 619174
rect 293866 618938 294102 619174
rect 293546 618618 293782 618854
rect 293866 618618 294102 618854
rect 293546 582938 293782 583174
rect 293866 582938 294102 583174
rect 293546 582618 293782 582854
rect 293866 582618 294102 582854
rect 293546 546938 293782 547174
rect 293866 546938 294102 547174
rect 293546 546618 293782 546854
rect 293866 546618 294102 546854
rect 293546 510938 293782 511174
rect 293866 510938 294102 511174
rect 293546 510618 293782 510854
rect 293866 510618 294102 510854
rect 297266 694658 297502 694894
rect 297586 694658 297822 694894
rect 297266 694338 297502 694574
rect 297586 694338 297822 694574
rect 297266 658658 297502 658894
rect 297586 658658 297822 658894
rect 297266 658338 297502 658574
rect 297586 658338 297822 658574
rect 297266 622658 297502 622894
rect 297586 622658 297822 622894
rect 297266 622338 297502 622574
rect 297586 622338 297822 622574
rect 297266 586658 297502 586894
rect 297586 586658 297822 586894
rect 297266 586338 297502 586574
rect 297586 586338 297822 586574
rect 297266 550658 297502 550894
rect 297586 550658 297822 550894
rect 297266 550338 297502 550574
rect 297586 550338 297822 550574
rect 297266 514658 297502 514894
rect 297586 514658 297822 514894
rect 297266 514338 297502 514574
rect 297586 514338 297822 514574
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 300986 698378 301222 698614
rect 301306 698378 301542 698614
rect 300986 698058 301222 698294
rect 301306 698058 301542 698294
rect 300986 662378 301222 662614
rect 301306 662378 301542 662614
rect 300986 662058 301222 662294
rect 301306 662058 301542 662294
rect 300986 626378 301222 626614
rect 301306 626378 301542 626614
rect 300986 626058 301222 626294
rect 301306 626058 301542 626294
rect 300986 590378 301222 590614
rect 301306 590378 301542 590614
rect 300986 590058 301222 590294
rect 301306 590058 301542 590294
rect 300986 554378 301222 554614
rect 301306 554378 301542 554614
rect 300986 554058 301222 554294
rect 301306 554058 301542 554294
rect 300986 518378 301222 518614
rect 301306 518378 301542 518614
rect 300986 518058 301222 518294
rect 301306 518058 301542 518294
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 307826 669218 308062 669454
rect 308146 669218 308382 669454
rect 307826 668898 308062 669134
rect 308146 668898 308382 669134
rect 307826 633218 308062 633454
rect 308146 633218 308382 633454
rect 307826 632898 308062 633134
rect 308146 632898 308382 633134
rect 307826 597218 308062 597454
rect 308146 597218 308382 597454
rect 307826 596898 308062 597134
rect 308146 596898 308382 597134
rect 307826 561218 308062 561454
rect 308146 561218 308382 561454
rect 307826 560898 308062 561134
rect 308146 560898 308382 561134
rect 307826 525218 308062 525454
rect 308146 525218 308382 525454
rect 307826 524898 308062 525134
rect 308146 524898 308382 525134
rect 307826 489218 308062 489454
rect 308146 489218 308382 489454
rect 307826 488898 308062 489134
rect 308146 488898 308382 489134
rect 311546 672938 311782 673174
rect 311866 672938 312102 673174
rect 311546 672618 311782 672854
rect 311866 672618 312102 672854
rect 311546 636938 311782 637174
rect 311866 636938 312102 637174
rect 311546 636618 311782 636854
rect 311866 636618 312102 636854
rect 311546 600938 311782 601174
rect 311866 600938 312102 601174
rect 311546 600618 311782 600854
rect 311866 600618 312102 600854
rect 311546 564938 311782 565174
rect 311866 564938 312102 565174
rect 311546 564618 311782 564854
rect 311866 564618 312102 564854
rect 311546 528938 311782 529174
rect 311866 528938 312102 529174
rect 311546 528618 311782 528854
rect 311866 528618 312102 528854
rect 311546 492938 311782 493174
rect 311866 492938 312102 493174
rect 311546 492618 311782 492854
rect 311866 492618 312102 492854
rect 315266 676658 315502 676894
rect 315586 676658 315822 676894
rect 315266 676338 315502 676574
rect 315586 676338 315822 676574
rect 315266 640658 315502 640894
rect 315586 640658 315822 640894
rect 315266 640338 315502 640574
rect 315586 640338 315822 640574
rect 315266 604658 315502 604894
rect 315586 604658 315822 604894
rect 315266 604338 315502 604574
rect 315586 604338 315822 604574
rect 315266 568658 315502 568894
rect 315586 568658 315822 568894
rect 315266 568338 315502 568574
rect 315586 568338 315822 568574
rect 315266 532658 315502 532894
rect 315586 532658 315822 532894
rect 315266 532338 315502 532574
rect 315586 532338 315822 532574
rect 315266 496658 315502 496894
rect 315586 496658 315822 496894
rect 315266 496338 315502 496574
rect 315586 496338 315822 496574
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 318986 680378 319222 680614
rect 319306 680378 319542 680614
rect 318986 680058 319222 680294
rect 319306 680058 319542 680294
rect 318986 644378 319222 644614
rect 319306 644378 319542 644614
rect 318986 644058 319222 644294
rect 319306 644058 319542 644294
rect 318986 608378 319222 608614
rect 319306 608378 319542 608614
rect 318986 608058 319222 608294
rect 319306 608058 319542 608294
rect 318986 572378 319222 572614
rect 319306 572378 319542 572614
rect 318986 572058 319222 572294
rect 319306 572058 319542 572294
rect 318986 536378 319222 536614
rect 319306 536378 319542 536614
rect 318986 536058 319222 536294
rect 319306 536058 319542 536294
rect 318986 500378 319222 500614
rect 319306 500378 319542 500614
rect 318986 500058 319222 500294
rect 319306 500058 319542 500294
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 325826 687218 326062 687454
rect 326146 687218 326382 687454
rect 325826 686898 326062 687134
rect 326146 686898 326382 687134
rect 325826 651218 326062 651454
rect 326146 651218 326382 651454
rect 325826 650898 326062 651134
rect 326146 650898 326382 651134
rect 325826 615218 326062 615454
rect 326146 615218 326382 615454
rect 325826 614898 326062 615134
rect 326146 614898 326382 615134
rect 325826 579218 326062 579454
rect 326146 579218 326382 579454
rect 325826 578898 326062 579134
rect 326146 578898 326382 579134
rect 325826 543218 326062 543454
rect 326146 543218 326382 543454
rect 325826 542898 326062 543134
rect 326146 542898 326382 543134
rect 325826 507218 326062 507454
rect 326146 507218 326382 507454
rect 325826 506898 326062 507134
rect 326146 506898 326382 507134
rect 329546 690938 329782 691174
rect 329866 690938 330102 691174
rect 329546 690618 329782 690854
rect 329866 690618 330102 690854
rect 329546 654938 329782 655174
rect 329866 654938 330102 655174
rect 329546 654618 329782 654854
rect 329866 654618 330102 654854
rect 329546 618938 329782 619174
rect 329866 618938 330102 619174
rect 329546 618618 329782 618854
rect 329866 618618 330102 618854
rect 329546 582938 329782 583174
rect 329866 582938 330102 583174
rect 329546 582618 329782 582854
rect 329866 582618 330102 582854
rect 329546 546938 329782 547174
rect 329866 546938 330102 547174
rect 329546 546618 329782 546854
rect 329866 546618 330102 546854
rect 329546 510938 329782 511174
rect 329866 510938 330102 511174
rect 329546 510618 329782 510854
rect 329866 510618 330102 510854
rect 333266 694658 333502 694894
rect 333586 694658 333822 694894
rect 333266 694338 333502 694574
rect 333586 694338 333822 694574
rect 333266 658658 333502 658894
rect 333586 658658 333822 658894
rect 333266 658338 333502 658574
rect 333586 658338 333822 658574
rect 333266 622658 333502 622894
rect 333586 622658 333822 622894
rect 333266 622338 333502 622574
rect 333586 622338 333822 622574
rect 333266 586658 333502 586894
rect 333586 586658 333822 586894
rect 333266 586338 333502 586574
rect 333586 586338 333822 586574
rect 333266 550658 333502 550894
rect 333586 550658 333822 550894
rect 333266 550338 333502 550574
rect 333586 550338 333822 550574
rect 333266 514658 333502 514894
rect 333586 514658 333822 514894
rect 333266 514338 333502 514574
rect 333586 514338 333822 514574
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 336986 698378 337222 698614
rect 337306 698378 337542 698614
rect 336986 698058 337222 698294
rect 337306 698058 337542 698294
rect 336986 662378 337222 662614
rect 337306 662378 337542 662614
rect 336986 662058 337222 662294
rect 337306 662058 337542 662294
rect 336986 626378 337222 626614
rect 337306 626378 337542 626614
rect 336986 626058 337222 626294
rect 337306 626058 337542 626294
rect 336986 590378 337222 590614
rect 337306 590378 337542 590614
rect 336986 590058 337222 590294
rect 337306 590058 337542 590294
rect 336986 554378 337222 554614
rect 337306 554378 337542 554614
rect 336986 554058 337222 554294
rect 337306 554058 337542 554294
rect 336986 518378 337222 518614
rect 337306 518378 337542 518614
rect 336986 518058 337222 518294
rect 337306 518058 337542 518294
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 343826 669218 344062 669454
rect 344146 669218 344382 669454
rect 343826 668898 344062 669134
rect 344146 668898 344382 669134
rect 343826 633218 344062 633454
rect 344146 633218 344382 633454
rect 343826 632898 344062 633134
rect 344146 632898 344382 633134
rect 343826 597218 344062 597454
rect 344146 597218 344382 597454
rect 343826 596898 344062 597134
rect 344146 596898 344382 597134
rect 343826 561218 344062 561454
rect 344146 561218 344382 561454
rect 343826 560898 344062 561134
rect 344146 560898 344382 561134
rect 343826 525218 344062 525454
rect 344146 525218 344382 525454
rect 343826 524898 344062 525134
rect 344146 524898 344382 525134
rect 343826 489218 344062 489454
rect 344146 489218 344382 489454
rect 343826 488898 344062 489134
rect 344146 488898 344382 489134
rect 347546 672938 347782 673174
rect 347866 672938 348102 673174
rect 347546 672618 347782 672854
rect 347866 672618 348102 672854
rect 347546 636938 347782 637174
rect 347866 636938 348102 637174
rect 347546 636618 347782 636854
rect 347866 636618 348102 636854
rect 347546 600938 347782 601174
rect 347866 600938 348102 601174
rect 347546 600618 347782 600854
rect 347866 600618 348102 600854
rect 347546 564938 347782 565174
rect 347866 564938 348102 565174
rect 347546 564618 347782 564854
rect 347866 564618 348102 564854
rect 347546 528938 347782 529174
rect 347866 528938 348102 529174
rect 347546 528618 347782 528854
rect 347866 528618 348102 528854
rect 347546 492938 347782 493174
rect 347866 492938 348102 493174
rect 347546 492618 347782 492854
rect 347866 492618 348102 492854
rect 351266 676658 351502 676894
rect 351586 676658 351822 676894
rect 351266 676338 351502 676574
rect 351586 676338 351822 676574
rect 351266 640658 351502 640894
rect 351586 640658 351822 640894
rect 351266 640338 351502 640574
rect 351586 640338 351822 640574
rect 351266 604658 351502 604894
rect 351586 604658 351822 604894
rect 351266 604338 351502 604574
rect 351586 604338 351822 604574
rect 351266 568658 351502 568894
rect 351586 568658 351822 568894
rect 351266 568338 351502 568574
rect 351586 568338 351822 568574
rect 351266 532658 351502 532894
rect 351586 532658 351822 532894
rect 351266 532338 351502 532574
rect 351586 532338 351822 532574
rect 351266 496658 351502 496894
rect 351586 496658 351822 496894
rect 351266 496338 351502 496574
rect 351586 496338 351822 496574
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 354986 680378 355222 680614
rect 355306 680378 355542 680614
rect 354986 680058 355222 680294
rect 355306 680058 355542 680294
rect 354986 644378 355222 644614
rect 355306 644378 355542 644614
rect 354986 644058 355222 644294
rect 355306 644058 355542 644294
rect 354986 608378 355222 608614
rect 355306 608378 355542 608614
rect 354986 608058 355222 608294
rect 355306 608058 355542 608294
rect 354986 572378 355222 572614
rect 355306 572378 355542 572614
rect 354986 572058 355222 572294
rect 355306 572058 355542 572294
rect 354986 536378 355222 536614
rect 355306 536378 355542 536614
rect 354986 536058 355222 536294
rect 355306 536058 355542 536294
rect 354986 500378 355222 500614
rect 355306 500378 355542 500614
rect 354986 500058 355222 500294
rect 355306 500058 355542 500294
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 361826 687218 362062 687454
rect 362146 687218 362382 687454
rect 361826 686898 362062 687134
rect 362146 686898 362382 687134
rect 361826 651218 362062 651454
rect 362146 651218 362382 651454
rect 361826 650898 362062 651134
rect 362146 650898 362382 651134
rect 361826 615218 362062 615454
rect 362146 615218 362382 615454
rect 361826 614898 362062 615134
rect 362146 614898 362382 615134
rect 361826 579218 362062 579454
rect 362146 579218 362382 579454
rect 361826 578898 362062 579134
rect 362146 578898 362382 579134
rect 361826 543218 362062 543454
rect 362146 543218 362382 543454
rect 361826 542898 362062 543134
rect 362146 542898 362382 543134
rect 361826 507218 362062 507454
rect 362146 507218 362382 507454
rect 361826 506898 362062 507134
rect 362146 506898 362382 507134
rect 221008 471218 221244 471454
rect 221008 470898 221244 471134
rect 355376 471218 355612 471454
rect 355376 470898 355612 471134
rect 361826 471218 362062 471454
rect 362146 471218 362382 471454
rect 361826 470898 362062 471134
rect 362146 470898 362382 471134
rect 220328 453218 220564 453454
rect 220328 452898 220564 453134
rect 356056 453218 356292 453454
rect 356056 452898 356292 453134
rect 221008 435218 221244 435454
rect 221008 434898 221244 435134
rect 355376 435218 355612 435454
rect 355376 434898 355612 435134
rect 361826 435218 362062 435454
rect 362146 435218 362382 435454
rect 361826 434898 362062 435134
rect 362146 434898 362382 435134
rect 220328 417218 220564 417454
rect 220328 416898 220564 417134
rect 356056 417218 356292 417454
rect 356056 416898 356292 417134
rect 221546 366938 221782 367174
rect 221866 366938 222102 367174
rect 221546 366618 221782 366854
rect 221866 366618 222102 366854
rect 221546 330938 221782 331174
rect 221866 330938 222102 331174
rect 221546 330618 221782 330854
rect 221866 330618 222102 330854
rect 221546 294938 221782 295174
rect 221866 294938 222102 295174
rect 221546 294618 221782 294854
rect 221866 294618 222102 294854
rect 221546 258938 221782 259174
rect 221866 258938 222102 259174
rect 221546 258618 221782 258854
rect 221866 258618 222102 258854
rect 64250 219218 64486 219454
rect 64250 218898 64486 219134
rect 94970 219218 95206 219454
rect 94970 218898 95206 219134
rect 125690 219218 125926 219454
rect 125690 218898 125926 219134
rect 156410 219218 156646 219454
rect 156410 218898 156646 219134
rect 187130 219218 187366 219454
rect 187130 218898 187366 219134
rect 217850 219218 218086 219454
rect 217850 218898 218086 219134
rect 55826 201218 56062 201454
rect 56146 201218 56382 201454
rect 55826 200898 56062 201134
rect 56146 200898 56382 201134
rect 79610 201218 79846 201454
rect 79610 200898 79846 201134
rect 110330 201218 110566 201454
rect 110330 200898 110566 201134
rect 141050 201218 141286 201454
rect 141050 200898 141286 201134
rect 171770 201218 172006 201454
rect 171770 200898 172006 201134
rect 202490 201218 202726 201454
rect 202490 200898 202726 201134
rect 64250 183218 64486 183454
rect 64250 182898 64486 183134
rect 94970 183218 95206 183454
rect 94970 182898 95206 183134
rect 125690 183218 125926 183454
rect 125690 182898 125926 183134
rect 156410 183218 156646 183454
rect 156410 182898 156646 183134
rect 187130 183218 187366 183454
rect 187130 182898 187366 183134
rect 217850 183218 218086 183454
rect 217850 182898 218086 183134
rect 55826 165218 56062 165454
rect 56146 165218 56382 165454
rect 55826 164898 56062 165134
rect 56146 164898 56382 165134
rect 79610 165218 79846 165454
rect 79610 164898 79846 165134
rect 110330 165218 110566 165454
rect 110330 164898 110566 165134
rect 141050 165218 141286 165454
rect 141050 164898 141286 165134
rect 171770 165218 172006 165454
rect 171770 164898 172006 165134
rect 202490 165218 202726 165454
rect 202490 164898 202726 165134
rect 64250 147218 64486 147454
rect 64250 146898 64486 147134
rect 94970 147218 95206 147454
rect 94970 146898 95206 147134
rect 125690 147218 125926 147454
rect 125690 146898 125926 147134
rect 156410 147218 156646 147454
rect 156410 146898 156646 147134
rect 187130 147218 187366 147454
rect 187130 146898 187366 147134
rect 217850 147218 218086 147454
rect 217850 146898 218086 147134
rect 55826 129218 56062 129454
rect 56146 129218 56382 129454
rect 55826 128898 56062 129134
rect 56146 128898 56382 129134
rect 79610 129218 79846 129454
rect 79610 128898 79846 129134
rect 110330 129218 110566 129454
rect 110330 128898 110566 129134
rect 141050 129218 141286 129454
rect 141050 128898 141286 129134
rect 171770 129218 172006 129454
rect 171770 128898 172006 129134
rect 202490 129218 202726 129454
rect 202490 128898 202726 129134
rect 64250 111218 64486 111454
rect 64250 110898 64486 111134
rect 94970 111218 95206 111454
rect 94970 110898 95206 111134
rect 125690 111218 125926 111454
rect 125690 110898 125926 111134
rect 156410 111218 156646 111454
rect 156410 110898 156646 111134
rect 187130 111218 187366 111454
rect 187130 110898 187366 111134
rect 217850 111218 218086 111454
rect 217850 110898 218086 111134
rect 55826 93218 56062 93454
rect 56146 93218 56382 93454
rect 55826 92898 56062 93134
rect 56146 92898 56382 93134
rect 79610 93218 79846 93454
rect 79610 92898 79846 93134
rect 110330 93218 110566 93454
rect 110330 92898 110566 93134
rect 141050 93218 141286 93454
rect 141050 92898 141286 93134
rect 171770 93218 172006 93454
rect 171770 92898 172006 93134
rect 202490 93218 202726 93454
rect 202490 92898 202726 93134
rect 64250 75218 64486 75454
rect 64250 74898 64486 75134
rect 94970 75218 95206 75454
rect 94970 74898 95206 75134
rect 125690 75218 125926 75454
rect 125690 74898 125926 75134
rect 156410 75218 156646 75454
rect 156410 74898 156646 75134
rect 187130 75218 187366 75454
rect 187130 74898 187366 75134
rect 217850 75218 218086 75454
rect 217850 74898 218086 75134
rect 225266 370658 225502 370894
rect 225586 370658 225822 370894
rect 225266 370338 225502 370574
rect 225586 370338 225822 370574
rect 225266 334658 225502 334894
rect 225586 334658 225822 334894
rect 225266 334338 225502 334574
rect 225586 334338 225822 334574
rect 225266 298658 225502 298894
rect 225586 298658 225822 298894
rect 225266 298338 225502 298574
rect 225586 298338 225822 298574
rect 225266 262658 225502 262894
rect 225586 262658 225822 262894
rect 225266 262338 225502 262574
rect 225586 262338 225822 262574
rect 55826 57218 56062 57454
rect 56146 57218 56382 57454
rect 55826 56898 56062 57134
rect 56146 56898 56382 57134
rect 55826 21218 56062 21454
rect 56146 21218 56382 21454
rect 55826 20898 56062 21134
rect 56146 20898 56382 21134
rect 55826 -1542 56062 -1306
rect 56146 -1542 56382 -1306
rect 55826 -1862 56062 -1626
rect 56146 -1862 56382 -1626
rect 59546 24938 59782 25174
rect 59866 24938 60102 25174
rect 59546 24618 59782 24854
rect 59866 24618 60102 24854
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 28658 63502 28894
rect 63586 28658 63822 28894
rect 63266 28338 63502 28574
rect 63586 28338 63822 28574
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 66986 32378 67222 32614
rect 67306 32378 67542 32614
rect 66986 32058 67222 32294
rect 67306 32058 67542 32294
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 73826 39218 74062 39454
rect 74146 39218 74382 39454
rect 73826 38898 74062 39134
rect 74146 38898 74382 39134
rect 73826 3218 74062 3454
rect 74146 3218 74382 3454
rect 73826 2898 74062 3134
rect 74146 2898 74382 3134
rect 73826 -582 74062 -346
rect 74146 -582 74382 -346
rect 73826 -902 74062 -666
rect 74146 -902 74382 -666
rect 77546 42938 77782 43174
rect 77866 42938 78102 43174
rect 77546 42618 77782 42854
rect 77866 42618 78102 42854
rect 77546 6938 77782 7174
rect 77866 6938 78102 7174
rect 77546 6618 77782 6854
rect 77866 6618 78102 6854
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 46658 81502 46894
rect 81586 46658 81822 46894
rect 81266 46338 81502 46574
rect 81586 46338 81822 46574
rect 81266 10658 81502 10894
rect 81586 10658 81822 10894
rect 81266 10338 81502 10574
rect 81586 10338 81822 10574
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 84986 50378 85222 50614
rect 85306 50378 85542 50614
rect 84986 50058 85222 50294
rect 85306 50058 85542 50294
rect 84986 14378 85222 14614
rect 85306 14378 85542 14614
rect 84986 14058 85222 14294
rect 85306 14058 85542 14294
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 91826 57218 92062 57454
rect 92146 57218 92382 57454
rect 91826 56898 92062 57134
rect 92146 56898 92382 57134
rect 91826 21218 92062 21454
rect 92146 21218 92382 21454
rect 91826 20898 92062 21134
rect 92146 20898 92382 21134
rect 91826 -1542 92062 -1306
rect 92146 -1542 92382 -1306
rect 91826 -1862 92062 -1626
rect 92146 -1862 92382 -1626
rect 95546 24938 95782 25174
rect 95866 24938 96102 25174
rect 95546 24618 95782 24854
rect 95866 24618 96102 24854
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 28658 99502 28894
rect 99586 28658 99822 28894
rect 99266 28338 99502 28574
rect 99586 28338 99822 28574
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 102986 32378 103222 32614
rect 103306 32378 103542 32614
rect 102986 32058 103222 32294
rect 103306 32058 103542 32294
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 109826 39218 110062 39454
rect 110146 39218 110382 39454
rect 109826 38898 110062 39134
rect 110146 38898 110382 39134
rect 109826 3218 110062 3454
rect 110146 3218 110382 3454
rect 109826 2898 110062 3134
rect 110146 2898 110382 3134
rect 109826 -582 110062 -346
rect 110146 -582 110382 -346
rect 109826 -902 110062 -666
rect 110146 -902 110382 -666
rect 113546 42938 113782 43174
rect 113866 42938 114102 43174
rect 113546 42618 113782 42854
rect 113866 42618 114102 42854
rect 113546 6938 113782 7174
rect 113866 6938 114102 7174
rect 113546 6618 113782 6854
rect 113866 6618 114102 6854
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 46658 117502 46894
rect 117586 46658 117822 46894
rect 117266 46338 117502 46574
rect 117586 46338 117822 46574
rect 117266 10658 117502 10894
rect 117586 10658 117822 10894
rect 117266 10338 117502 10574
rect 117586 10338 117822 10574
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 120986 50378 121222 50614
rect 121306 50378 121542 50614
rect 120986 50058 121222 50294
rect 121306 50058 121542 50294
rect 120986 14378 121222 14614
rect 121306 14378 121542 14614
rect 120986 14058 121222 14294
rect 121306 14058 121542 14294
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 127826 57218 128062 57454
rect 128146 57218 128382 57454
rect 127826 56898 128062 57134
rect 128146 56898 128382 57134
rect 127826 21218 128062 21454
rect 128146 21218 128382 21454
rect 127826 20898 128062 21134
rect 128146 20898 128382 21134
rect 127826 -1542 128062 -1306
rect 128146 -1542 128382 -1306
rect 127826 -1862 128062 -1626
rect 128146 -1862 128382 -1626
rect 131546 24938 131782 25174
rect 131866 24938 132102 25174
rect 131546 24618 131782 24854
rect 131866 24618 132102 24854
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 28658 135502 28894
rect 135586 28658 135822 28894
rect 135266 28338 135502 28574
rect 135586 28338 135822 28574
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 138986 32378 139222 32614
rect 139306 32378 139542 32614
rect 138986 32058 139222 32294
rect 139306 32058 139542 32294
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 145826 39218 146062 39454
rect 146146 39218 146382 39454
rect 145826 38898 146062 39134
rect 146146 38898 146382 39134
rect 145826 3218 146062 3454
rect 146146 3218 146382 3454
rect 145826 2898 146062 3134
rect 146146 2898 146382 3134
rect 145826 -582 146062 -346
rect 146146 -582 146382 -346
rect 145826 -902 146062 -666
rect 146146 -902 146382 -666
rect 149546 42938 149782 43174
rect 149866 42938 150102 43174
rect 149546 42618 149782 42854
rect 149866 42618 150102 42854
rect 149546 6938 149782 7174
rect 149866 6938 150102 7174
rect 149546 6618 149782 6854
rect 149866 6618 150102 6854
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 46658 153502 46894
rect 153586 46658 153822 46894
rect 153266 46338 153502 46574
rect 153586 46338 153822 46574
rect 153266 10658 153502 10894
rect 153586 10658 153822 10894
rect 153266 10338 153502 10574
rect 153586 10338 153822 10574
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 156986 50378 157222 50614
rect 157306 50378 157542 50614
rect 156986 50058 157222 50294
rect 157306 50058 157542 50294
rect 156986 14378 157222 14614
rect 157306 14378 157542 14614
rect 156986 14058 157222 14294
rect 157306 14058 157542 14294
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 163826 57218 164062 57454
rect 164146 57218 164382 57454
rect 163826 56898 164062 57134
rect 164146 56898 164382 57134
rect 163826 21218 164062 21454
rect 164146 21218 164382 21454
rect 163826 20898 164062 21134
rect 164146 20898 164382 21134
rect 163826 -1542 164062 -1306
rect 164146 -1542 164382 -1306
rect 163826 -1862 164062 -1626
rect 164146 -1862 164382 -1626
rect 167546 24938 167782 25174
rect 167866 24938 168102 25174
rect 167546 24618 167782 24854
rect 167866 24618 168102 24854
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 28658 171502 28894
rect 171586 28658 171822 28894
rect 171266 28338 171502 28574
rect 171586 28338 171822 28574
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 174986 32378 175222 32614
rect 175306 32378 175542 32614
rect 174986 32058 175222 32294
rect 175306 32058 175542 32294
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 181826 39218 182062 39454
rect 182146 39218 182382 39454
rect 181826 38898 182062 39134
rect 182146 38898 182382 39134
rect 181826 3218 182062 3454
rect 182146 3218 182382 3454
rect 181826 2898 182062 3134
rect 182146 2898 182382 3134
rect 181826 -582 182062 -346
rect 182146 -582 182382 -346
rect 181826 -902 182062 -666
rect 182146 -902 182382 -666
rect 185546 42938 185782 43174
rect 185866 42938 186102 43174
rect 185546 42618 185782 42854
rect 185866 42618 186102 42854
rect 185546 6938 185782 7174
rect 185866 6938 186102 7174
rect 185546 6618 185782 6854
rect 185866 6618 186102 6854
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 46658 189502 46894
rect 189586 46658 189822 46894
rect 189266 46338 189502 46574
rect 189586 46338 189822 46574
rect 189266 10658 189502 10894
rect 189586 10658 189822 10894
rect 189266 10338 189502 10574
rect 189586 10338 189822 10574
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 192986 50378 193222 50614
rect 193306 50378 193542 50614
rect 192986 50058 193222 50294
rect 193306 50058 193542 50294
rect 192986 14378 193222 14614
rect 193306 14378 193542 14614
rect 192986 14058 193222 14294
rect 193306 14058 193542 14294
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 199826 57218 200062 57454
rect 200146 57218 200382 57454
rect 199826 56898 200062 57134
rect 200146 56898 200382 57134
rect 199826 21218 200062 21454
rect 200146 21218 200382 21454
rect 199826 20898 200062 21134
rect 200146 20898 200382 21134
rect 199826 -1542 200062 -1306
rect 200146 -1542 200382 -1306
rect 199826 -1862 200062 -1626
rect 200146 -1862 200382 -1626
rect 203546 24938 203782 25174
rect 203866 24938 204102 25174
rect 203546 24618 203782 24854
rect 203866 24618 204102 24854
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 28658 207502 28894
rect 207586 28658 207822 28894
rect 207266 28338 207502 28574
rect 207586 28338 207822 28574
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 210986 32378 211222 32614
rect 211306 32378 211542 32614
rect 210986 32058 211222 32294
rect 211306 32058 211542 32294
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 217826 39218 218062 39454
rect 218146 39218 218382 39454
rect 217826 38898 218062 39134
rect 218146 38898 218382 39134
rect 217826 3218 218062 3454
rect 218146 3218 218382 3454
rect 217826 2898 218062 3134
rect 218146 2898 218382 3134
rect 217826 -582 218062 -346
rect 218146 -582 218382 -346
rect 217826 -902 218062 -666
rect 218146 -902 218382 -666
rect 228986 374378 229222 374614
rect 229306 374378 229542 374614
rect 228986 374058 229222 374294
rect 229306 374058 229542 374294
rect 228986 338378 229222 338614
rect 229306 338378 229542 338614
rect 228986 338058 229222 338294
rect 229306 338058 229542 338294
rect 228986 302378 229222 302614
rect 229306 302378 229542 302614
rect 228986 302058 229222 302294
rect 229306 302058 229542 302294
rect 228986 266378 229222 266614
rect 229306 266378 229542 266614
rect 228986 266058 229222 266294
rect 229306 266058 229542 266294
rect 228986 230378 229222 230614
rect 229306 230378 229542 230614
rect 228986 230058 229222 230294
rect 229306 230058 229542 230294
rect 228986 194378 229222 194614
rect 229306 194378 229542 194614
rect 228986 194058 229222 194294
rect 229306 194058 229542 194294
rect 228986 158378 229222 158614
rect 229306 158378 229542 158614
rect 228986 158058 229222 158294
rect 229306 158058 229542 158294
rect 228986 122378 229222 122614
rect 229306 122378 229542 122614
rect 228986 122058 229222 122294
rect 229306 122058 229542 122294
rect 228986 86378 229222 86614
rect 229306 86378 229542 86614
rect 228986 86058 229222 86294
rect 229306 86058 229542 86294
rect 221546 42938 221782 43174
rect 221866 42938 222102 43174
rect 221546 42618 221782 42854
rect 221866 42618 222102 42854
rect 221546 6938 221782 7174
rect 221866 6938 222102 7174
rect 221546 6618 221782 6854
rect 221866 6618 222102 6854
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 46658 225502 46894
rect 225586 46658 225822 46894
rect 225266 46338 225502 46574
rect 225586 46338 225822 46574
rect 225266 10658 225502 10894
rect 225586 10658 225822 10894
rect 225266 10338 225502 10574
rect 225586 10338 225822 10574
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 228986 50378 229222 50614
rect 229306 50378 229542 50614
rect 228986 50058 229222 50294
rect 229306 50058 229542 50294
rect 228986 14378 229222 14614
rect 229306 14378 229542 14614
rect 228986 14058 229222 14294
rect 229306 14058 229542 14294
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 235826 381218 236062 381454
rect 236146 381218 236382 381454
rect 235826 380898 236062 381134
rect 236146 380898 236382 381134
rect 235826 345218 236062 345454
rect 236146 345218 236382 345454
rect 235826 344898 236062 345134
rect 236146 344898 236382 345134
rect 235826 309218 236062 309454
rect 236146 309218 236382 309454
rect 235826 308898 236062 309134
rect 236146 308898 236382 309134
rect 235826 273218 236062 273454
rect 236146 273218 236382 273454
rect 235826 272898 236062 273134
rect 236146 272898 236382 273134
rect 235826 237218 236062 237454
rect 236146 237218 236382 237454
rect 235826 236898 236062 237134
rect 236146 236898 236382 237134
rect 235826 201218 236062 201454
rect 236146 201218 236382 201454
rect 235826 200898 236062 201134
rect 236146 200898 236382 201134
rect 235826 165218 236062 165454
rect 236146 165218 236382 165454
rect 235826 164898 236062 165134
rect 236146 164898 236382 165134
rect 235826 129218 236062 129454
rect 236146 129218 236382 129454
rect 235826 128898 236062 129134
rect 236146 128898 236382 129134
rect 235826 93218 236062 93454
rect 236146 93218 236382 93454
rect 235826 92898 236062 93134
rect 236146 92898 236382 93134
rect 235826 57218 236062 57454
rect 236146 57218 236382 57454
rect 235826 56898 236062 57134
rect 236146 56898 236382 57134
rect 235826 21218 236062 21454
rect 236146 21218 236382 21454
rect 235826 20898 236062 21134
rect 236146 20898 236382 21134
rect 235826 -1542 236062 -1306
rect 236146 -1542 236382 -1306
rect 235826 -1862 236062 -1626
rect 236146 -1862 236382 -1626
rect 239546 384938 239782 385174
rect 239866 384938 240102 385174
rect 239546 384618 239782 384854
rect 239866 384618 240102 384854
rect 239546 348938 239782 349174
rect 239866 348938 240102 349174
rect 239546 348618 239782 348854
rect 239866 348618 240102 348854
rect 239546 312938 239782 313174
rect 239866 312938 240102 313174
rect 239546 312618 239782 312854
rect 239866 312618 240102 312854
rect 239546 276938 239782 277174
rect 239866 276938 240102 277174
rect 239546 276618 239782 276854
rect 239866 276618 240102 276854
rect 239546 240938 239782 241174
rect 239866 240938 240102 241174
rect 239546 240618 239782 240854
rect 239866 240618 240102 240854
rect 239546 204938 239782 205174
rect 239866 204938 240102 205174
rect 239546 204618 239782 204854
rect 239866 204618 240102 204854
rect 239546 168938 239782 169174
rect 239866 168938 240102 169174
rect 239546 168618 239782 168854
rect 239866 168618 240102 168854
rect 239546 132938 239782 133174
rect 239866 132938 240102 133174
rect 239546 132618 239782 132854
rect 239866 132618 240102 132854
rect 239546 96938 239782 97174
rect 239866 96938 240102 97174
rect 239546 96618 239782 96854
rect 239866 96618 240102 96854
rect 239546 60938 239782 61174
rect 239866 60938 240102 61174
rect 239546 60618 239782 60854
rect 239866 60618 240102 60854
rect 239546 24938 239782 25174
rect 239866 24938 240102 25174
rect 239546 24618 239782 24854
rect 239866 24618 240102 24854
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 388658 243502 388894
rect 243586 388658 243822 388894
rect 243266 388338 243502 388574
rect 243586 388338 243822 388574
rect 243266 352658 243502 352894
rect 243586 352658 243822 352894
rect 243266 352338 243502 352574
rect 243586 352338 243822 352574
rect 243266 316658 243502 316894
rect 243586 316658 243822 316894
rect 243266 316338 243502 316574
rect 243586 316338 243822 316574
rect 243266 280658 243502 280894
rect 243586 280658 243822 280894
rect 243266 280338 243502 280574
rect 243586 280338 243822 280574
rect 243266 244658 243502 244894
rect 243586 244658 243822 244894
rect 243266 244338 243502 244574
rect 243586 244338 243822 244574
rect 243266 208658 243502 208894
rect 243586 208658 243822 208894
rect 243266 208338 243502 208574
rect 243586 208338 243822 208574
rect 243266 172658 243502 172894
rect 243586 172658 243822 172894
rect 243266 172338 243502 172574
rect 243586 172338 243822 172574
rect 243266 136658 243502 136894
rect 243586 136658 243822 136894
rect 243266 136338 243502 136574
rect 243586 136338 243822 136574
rect 243266 100658 243502 100894
rect 243586 100658 243822 100894
rect 243266 100338 243502 100574
rect 243586 100338 243822 100574
rect 243266 64658 243502 64894
rect 243586 64658 243822 64894
rect 243266 64338 243502 64574
rect 243586 64338 243822 64574
rect 243266 28658 243502 28894
rect 243586 28658 243822 28894
rect 243266 28338 243502 28574
rect 243586 28338 243822 28574
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 246986 392378 247222 392614
rect 247306 392378 247542 392614
rect 246986 392058 247222 392294
rect 247306 392058 247542 392294
rect 246986 356378 247222 356614
rect 247306 356378 247542 356614
rect 246986 356058 247222 356294
rect 247306 356058 247542 356294
rect 246986 320378 247222 320614
rect 247306 320378 247542 320614
rect 246986 320058 247222 320294
rect 247306 320058 247542 320294
rect 246986 284378 247222 284614
rect 247306 284378 247542 284614
rect 246986 284058 247222 284294
rect 247306 284058 247542 284294
rect 246986 248378 247222 248614
rect 247306 248378 247542 248614
rect 246986 248058 247222 248294
rect 247306 248058 247542 248294
rect 246986 212378 247222 212614
rect 247306 212378 247542 212614
rect 246986 212058 247222 212294
rect 247306 212058 247542 212294
rect 246986 176378 247222 176614
rect 247306 176378 247542 176614
rect 246986 176058 247222 176294
rect 247306 176058 247542 176294
rect 246986 140378 247222 140614
rect 247306 140378 247542 140614
rect 246986 140058 247222 140294
rect 247306 140058 247542 140294
rect 246986 104378 247222 104614
rect 247306 104378 247542 104614
rect 246986 104058 247222 104294
rect 247306 104058 247542 104294
rect 246986 68378 247222 68614
rect 247306 68378 247542 68614
rect 246986 68058 247222 68294
rect 247306 68058 247542 68294
rect 246986 32378 247222 32614
rect 247306 32378 247542 32614
rect 246986 32058 247222 32294
rect 247306 32058 247542 32294
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 253826 363218 254062 363454
rect 254146 363218 254382 363454
rect 253826 362898 254062 363134
rect 254146 362898 254382 363134
rect 253826 327218 254062 327454
rect 254146 327218 254382 327454
rect 253826 326898 254062 327134
rect 254146 326898 254382 327134
rect 253826 291218 254062 291454
rect 254146 291218 254382 291454
rect 253826 290898 254062 291134
rect 254146 290898 254382 291134
rect 253826 255218 254062 255454
rect 254146 255218 254382 255454
rect 253826 254898 254062 255134
rect 254146 254898 254382 255134
rect 253826 219218 254062 219454
rect 254146 219218 254382 219454
rect 253826 218898 254062 219134
rect 254146 218898 254382 219134
rect 253826 183218 254062 183454
rect 254146 183218 254382 183454
rect 253826 182898 254062 183134
rect 254146 182898 254382 183134
rect 253826 147218 254062 147454
rect 254146 147218 254382 147454
rect 253826 146898 254062 147134
rect 254146 146898 254382 147134
rect 253826 111218 254062 111454
rect 254146 111218 254382 111454
rect 253826 110898 254062 111134
rect 254146 110898 254382 111134
rect 253826 75218 254062 75454
rect 254146 75218 254382 75454
rect 253826 74898 254062 75134
rect 254146 74898 254382 75134
rect 253826 39218 254062 39454
rect 254146 39218 254382 39454
rect 253826 38898 254062 39134
rect 254146 38898 254382 39134
rect 253826 3218 254062 3454
rect 254146 3218 254382 3454
rect 253826 2898 254062 3134
rect 254146 2898 254382 3134
rect 253826 -582 254062 -346
rect 254146 -582 254382 -346
rect 253826 -902 254062 -666
rect 254146 -902 254382 -666
rect 257546 366938 257782 367174
rect 257866 366938 258102 367174
rect 257546 366618 257782 366854
rect 257866 366618 258102 366854
rect 257546 330938 257782 331174
rect 257866 330938 258102 331174
rect 257546 330618 257782 330854
rect 257866 330618 258102 330854
rect 257546 294938 257782 295174
rect 257866 294938 258102 295174
rect 257546 294618 257782 294854
rect 257866 294618 258102 294854
rect 257546 258938 257782 259174
rect 257866 258938 258102 259174
rect 257546 258618 257782 258854
rect 257866 258618 258102 258854
rect 257546 222938 257782 223174
rect 257866 222938 258102 223174
rect 257546 222618 257782 222854
rect 257866 222618 258102 222854
rect 257546 186938 257782 187174
rect 257866 186938 258102 187174
rect 257546 186618 257782 186854
rect 257866 186618 258102 186854
rect 257546 150938 257782 151174
rect 257866 150938 258102 151174
rect 257546 150618 257782 150854
rect 257866 150618 258102 150854
rect 257546 114938 257782 115174
rect 257866 114938 258102 115174
rect 257546 114618 257782 114854
rect 257866 114618 258102 114854
rect 257546 78938 257782 79174
rect 257866 78938 258102 79174
rect 257546 78618 257782 78854
rect 257866 78618 258102 78854
rect 257546 42938 257782 43174
rect 257866 42938 258102 43174
rect 257546 42618 257782 42854
rect 257866 42618 258102 42854
rect 257546 6938 257782 7174
rect 257866 6938 258102 7174
rect 257546 6618 257782 6854
rect 257866 6618 258102 6854
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 370658 261502 370894
rect 261586 370658 261822 370894
rect 261266 370338 261502 370574
rect 261586 370338 261822 370574
rect 261266 334658 261502 334894
rect 261586 334658 261822 334894
rect 261266 334338 261502 334574
rect 261586 334338 261822 334574
rect 261266 298658 261502 298894
rect 261586 298658 261822 298894
rect 261266 298338 261502 298574
rect 261586 298338 261822 298574
rect 261266 262658 261502 262894
rect 261586 262658 261822 262894
rect 261266 262338 261502 262574
rect 261586 262338 261822 262574
rect 261266 226658 261502 226894
rect 261586 226658 261822 226894
rect 261266 226338 261502 226574
rect 261586 226338 261822 226574
rect 261266 190658 261502 190894
rect 261586 190658 261822 190894
rect 261266 190338 261502 190574
rect 261586 190338 261822 190574
rect 261266 154658 261502 154894
rect 261586 154658 261822 154894
rect 261266 154338 261502 154574
rect 261586 154338 261822 154574
rect 261266 118658 261502 118894
rect 261586 118658 261822 118894
rect 261266 118338 261502 118574
rect 261586 118338 261822 118574
rect 261266 82658 261502 82894
rect 261586 82658 261822 82894
rect 261266 82338 261502 82574
rect 261586 82338 261822 82574
rect 261266 46658 261502 46894
rect 261586 46658 261822 46894
rect 261266 46338 261502 46574
rect 261586 46338 261822 46574
rect 261266 10658 261502 10894
rect 261586 10658 261822 10894
rect 261266 10338 261502 10574
rect 261586 10338 261822 10574
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 264986 374378 265222 374614
rect 265306 374378 265542 374614
rect 264986 374058 265222 374294
rect 265306 374058 265542 374294
rect 264986 338378 265222 338614
rect 265306 338378 265542 338614
rect 264986 338058 265222 338294
rect 265306 338058 265542 338294
rect 264986 302378 265222 302614
rect 265306 302378 265542 302614
rect 264986 302058 265222 302294
rect 265306 302058 265542 302294
rect 264986 266378 265222 266614
rect 265306 266378 265542 266614
rect 264986 266058 265222 266294
rect 265306 266058 265542 266294
rect 264986 230378 265222 230614
rect 265306 230378 265542 230614
rect 264986 230058 265222 230294
rect 265306 230058 265542 230294
rect 264986 194378 265222 194614
rect 265306 194378 265542 194614
rect 264986 194058 265222 194294
rect 265306 194058 265542 194294
rect 264986 158378 265222 158614
rect 265306 158378 265542 158614
rect 264986 158058 265222 158294
rect 265306 158058 265542 158294
rect 264986 122378 265222 122614
rect 265306 122378 265542 122614
rect 264986 122058 265222 122294
rect 265306 122058 265542 122294
rect 264986 86378 265222 86614
rect 265306 86378 265542 86614
rect 264986 86058 265222 86294
rect 265306 86058 265542 86294
rect 264986 50378 265222 50614
rect 265306 50378 265542 50614
rect 264986 50058 265222 50294
rect 265306 50058 265542 50294
rect 264986 14378 265222 14614
rect 265306 14378 265542 14614
rect 264986 14058 265222 14294
rect 265306 14058 265542 14294
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 271826 381218 272062 381454
rect 272146 381218 272382 381454
rect 271826 380898 272062 381134
rect 272146 380898 272382 381134
rect 271826 345218 272062 345454
rect 272146 345218 272382 345454
rect 271826 344898 272062 345134
rect 272146 344898 272382 345134
rect 271826 309218 272062 309454
rect 272146 309218 272382 309454
rect 271826 308898 272062 309134
rect 272146 308898 272382 309134
rect 271826 273218 272062 273454
rect 272146 273218 272382 273454
rect 271826 272898 272062 273134
rect 272146 272898 272382 273134
rect 271826 237218 272062 237454
rect 272146 237218 272382 237454
rect 271826 236898 272062 237134
rect 272146 236898 272382 237134
rect 271826 201218 272062 201454
rect 272146 201218 272382 201454
rect 271826 200898 272062 201134
rect 272146 200898 272382 201134
rect 271826 165218 272062 165454
rect 272146 165218 272382 165454
rect 271826 164898 272062 165134
rect 272146 164898 272382 165134
rect 271826 129218 272062 129454
rect 272146 129218 272382 129454
rect 271826 128898 272062 129134
rect 272146 128898 272382 129134
rect 271826 93218 272062 93454
rect 272146 93218 272382 93454
rect 271826 92898 272062 93134
rect 272146 92898 272382 93134
rect 271826 57218 272062 57454
rect 272146 57218 272382 57454
rect 271826 56898 272062 57134
rect 272146 56898 272382 57134
rect 271826 21218 272062 21454
rect 272146 21218 272382 21454
rect 271826 20898 272062 21134
rect 272146 20898 272382 21134
rect 271826 -1542 272062 -1306
rect 272146 -1542 272382 -1306
rect 271826 -1862 272062 -1626
rect 272146 -1862 272382 -1626
rect 275546 384938 275782 385174
rect 275866 384938 276102 385174
rect 275546 384618 275782 384854
rect 275866 384618 276102 384854
rect 275546 348938 275782 349174
rect 275866 348938 276102 349174
rect 275546 348618 275782 348854
rect 275866 348618 276102 348854
rect 275546 312938 275782 313174
rect 275866 312938 276102 313174
rect 275546 312618 275782 312854
rect 275866 312618 276102 312854
rect 275546 276938 275782 277174
rect 275866 276938 276102 277174
rect 275546 276618 275782 276854
rect 275866 276618 276102 276854
rect 275546 240938 275782 241174
rect 275866 240938 276102 241174
rect 275546 240618 275782 240854
rect 275866 240618 276102 240854
rect 275546 204938 275782 205174
rect 275866 204938 276102 205174
rect 275546 204618 275782 204854
rect 275866 204618 276102 204854
rect 275546 168938 275782 169174
rect 275866 168938 276102 169174
rect 275546 168618 275782 168854
rect 275866 168618 276102 168854
rect 275546 132938 275782 133174
rect 275866 132938 276102 133174
rect 275546 132618 275782 132854
rect 275866 132618 276102 132854
rect 275546 96938 275782 97174
rect 275866 96938 276102 97174
rect 275546 96618 275782 96854
rect 275866 96618 276102 96854
rect 275546 60938 275782 61174
rect 275866 60938 276102 61174
rect 275546 60618 275782 60854
rect 275866 60618 276102 60854
rect 275546 24938 275782 25174
rect 275866 24938 276102 25174
rect 275546 24618 275782 24854
rect 275866 24618 276102 24854
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 388658 279502 388894
rect 279586 388658 279822 388894
rect 279266 388338 279502 388574
rect 279586 388338 279822 388574
rect 279266 352658 279502 352894
rect 279586 352658 279822 352894
rect 279266 352338 279502 352574
rect 279586 352338 279822 352574
rect 279266 316658 279502 316894
rect 279586 316658 279822 316894
rect 279266 316338 279502 316574
rect 279586 316338 279822 316574
rect 279266 280658 279502 280894
rect 279586 280658 279822 280894
rect 279266 280338 279502 280574
rect 279586 280338 279822 280574
rect 279266 244658 279502 244894
rect 279586 244658 279822 244894
rect 279266 244338 279502 244574
rect 279586 244338 279822 244574
rect 279266 208658 279502 208894
rect 279586 208658 279822 208894
rect 279266 208338 279502 208574
rect 279586 208338 279822 208574
rect 279266 172658 279502 172894
rect 279586 172658 279822 172894
rect 279266 172338 279502 172574
rect 279586 172338 279822 172574
rect 279266 136658 279502 136894
rect 279586 136658 279822 136894
rect 279266 136338 279502 136574
rect 279586 136338 279822 136574
rect 279266 100658 279502 100894
rect 279586 100658 279822 100894
rect 279266 100338 279502 100574
rect 279586 100338 279822 100574
rect 279266 64658 279502 64894
rect 279586 64658 279822 64894
rect 279266 64338 279502 64574
rect 279586 64338 279822 64574
rect 279266 28658 279502 28894
rect 279586 28658 279822 28894
rect 279266 28338 279502 28574
rect 279586 28338 279822 28574
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 282986 392378 283222 392614
rect 283306 392378 283542 392614
rect 282986 392058 283222 392294
rect 283306 392058 283542 392294
rect 282986 356378 283222 356614
rect 283306 356378 283542 356614
rect 282986 356058 283222 356294
rect 283306 356058 283542 356294
rect 282986 320378 283222 320614
rect 283306 320378 283542 320614
rect 282986 320058 283222 320294
rect 283306 320058 283542 320294
rect 282986 284378 283222 284614
rect 283306 284378 283542 284614
rect 282986 284058 283222 284294
rect 283306 284058 283542 284294
rect 282986 248378 283222 248614
rect 283306 248378 283542 248614
rect 282986 248058 283222 248294
rect 283306 248058 283542 248294
rect 282986 212378 283222 212614
rect 283306 212378 283542 212614
rect 282986 212058 283222 212294
rect 283306 212058 283542 212294
rect 282986 176378 283222 176614
rect 283306 176378 283542 176614
rect 282986 176058 283222 176294
rect 283306 176058 283542 176294
rect 282986 140378 283222 140614
rect 283306 140378 283542 140614
rect 282986 140058 283222 140294
rect 283306 140058 283542 140294
rect 282986 104378 283222 104614
rect 283306 104378 283542 104614
rect 282986 104058 283222 104294
rect 283306 104058 283542 104294
rect 282986 68378 283222 68614
rect 283306 68378 283542 68614
rect 282986 68058 283222 68294
rect 283306 68058 283542 68294
rect 282986 32378 283222 32614
rect 283306 32378 283542 32614
rect 282986 32058 283222 32294
rect 283306 32058 283542 32294
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 289826 363218 290062 363454
rect 290146 363218 290382 363454
rect 289826 362898 290062 363134
rect 290146 362898 290382 363134
rect 289826 327218 290062 327454
rect 290146 327218 290382 327454
rect 289826 326898 290062 327134
rect 290146 326898 290382 327134
rect 289826 291218 290062 291454
rect 290146 291218 290382 291454
rect 289826 290898 290062 291134
rect 290146 290898 290382 291134
rect 289826 255218 290062 255454
rect 290146 255218 290382 255454
rect 289826 254898 290062 255134
rect 290146 254898 290382 255134
rect 289826 219218 290062 219454
rect 290146 219218 290382 219454
rect 289826 218898 290062 219134
rect 290146 218898 290382 219134
rect 289826 183218 290062 183454
rect 290146 183218 290382 183454
rect 289826 182898 290062 183134
rect 290146 182898 290382 183134
rect 289826 147218 290062 147454
rect 290146 147218 290382 147454
rect 289826 146898 290062 147134
rect 290146 146898 290382 147134
rect 289826 111218 290062 111454
rect 290146 111218 290382 111454
rect 289826 110898 290062 111134
rect 290146 110898 290382 111134
rect 289826 75218 290062 75454
rect 290146 75218 290382 75454
rect 289826 74898 290062 75134
rect 290146 74898 290382 75134
rect 289826 39218 290062 39454
rect 290146 39218 290382 39454
rect 289826 38898 290062 39134
rect 290146 38898 290382 39134
rect 289826 3218 290062 3454
rect 290146 3218 290382 3454
rect 289826 2898 290062 3134
rect 290146 2898 290382 3134
rect 289826 -582 290062 -346
rect 290146 -582 290382 -346
rect 289826 -902 290062 -666
rect 290146 -902 290382 -666
rect 293546 366938 293782 367174
rect 293866 366938 294102 367174
rect 293546 366618 293782 366854
rect 293866 366618 294102 366854
rect 293546 330938 293782 331174
rect 293866 330938 294102 331174
rect 293546 330618 293782 330854
rect 293866 330618 294102 330854
rect 293546 294938 293782 295174
rect 293866 294938 294102 295174
rect 293546 294618 293782 294854
rect 293866 294618 294102 294854
rect 293546 258938 293782 259174
rect 293866 258938 294102 259174
rect 293546 258618 293782 258854
rect 293866 258618 294102 258854
rect 293546 222938 293782 223174
rect 293866 222938 294102 223174
rect 293546 222618 293782 222854
rect 293866 222618 294102 222854
rect 293546 186938 293782 187174
rect 293866 186938 294102 187174
rect 293546 186618 293782 186854
rect 293866 186618 294102 186854
rect 293546 150938 293782 151174
rect 293866 150938 294102 151174
rect 293546 150618 293782 150854
rect 293866 150618 294102 150854
rect 293546 114938 293782 115174
rect 293866 114938 294102 115174
rect 293546 114618 293782 114854
rect 293866 114618 294102 114854
rect 293546 78938 293782 79174
rect 293866 78938 294102 79174
rect 293546 78618 293782 78854
rect 293866 78618 294102 78854
rect 293546 42938 293782 43174
rect 293866 42938 294102 43174
rect 293546 42618 293782 42854
rect 293866 42618 294102 42854
rect 293546 6938 293782 7174
rect 293866 6938 294102 7174
rect 293546 6618 293782 6854
rect 293866 6618 294102 6854
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 370658 297502 370894
rect 297586 370658 297822 370894
rect 297266 370338 297502 370574
rect 297586 370338 297822 370574
rect 297266 334658 297502 334894
rect 297586 334658 297822 334894
rect 297266 334338 297502 334574
rect 297586 334338 297822 334574
rect 297266 298658 297502 298894
rect 297586 298658 297822 298894
rect 297266 298338 297502 298574
rect 297586 298338 297822 298574
rect 297266 262658 297502 262894
rect 297586 262658 297822 262894
rect 297266 262338 297502 262574
rect 297586 262338 297822 262574
rect 297266 226658 297502 226894
rect 297586 226658 297822 226894
rect 297266 226338 297502 226574
rect 297586 226338 297822 226574
rect 297266 190658 297502 190894
rect 297586 190658 297822 190894
rect 297266 190338 297502 190574
rect 297586 190338 297822 190574
rect 297266 154658 297502 154894
rect 297586 154658 297822 154894
rect 297266 154338 297502 154574
rect 297586 154338 297822 154574
rect 297266 118658 297502 118894
rect 297586 118658 297822 118894
rect 297266 118338 297502 118574
rect 297586 118338 297822 118574
rect 297266 82658 297502 82894
rect 297586 82658 297822 82894
rect 297266 82338 297502 82574
rect 297586 82338 297822 82574
rect 297266 46658 297502 46894
rect 297586 46658 297822 46894
rect 297266 46338 297502 46574
rect 297586 46338 297822 46574
rect 297266 10658 297502 10894
rect 297586 10658 297822 10894
rect 297266 10338 297502 10574
rect 297586 10338 297822 10574
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 300986 374378 301222 374614
rect 301306 374378 301542 374614
rect 300986 374058 301222 374294
rect 301306 374058 301542 374294
rect 300986 338378 301222 338614
rect 301306 338378 301542 338614
rect 300986 338058 301222 338294
rect 301306 338058 301542 338294
rect 300986 302378 301222 302614
rect 301306 302378 301542 302614
rect 300986 302058 301222 302294
rect 301306 302058 301542 302294
rect 300986 266378 301222 266614
rect 301306 266378 301542 266614
rect 300986 266058 301222 266294
rect 301306 266058 301542 266294
rect 300986 230378 301222 230614
rect 301306 230378 301542 230614
rect 300986 230058 301222 230294
rect 301306 230058 301542 230294
rect 300986 194378 301222 194614
rect 301306 194378 301542 194614
rect 300986 194058 301222 194294
rect 301306 194058 301542 194294
rect 300986 158378 301222 158614
rect 301306 158378 301542 158614
rect 300986 158058 301222 158294
rect 301306 158058 301542 158294
rect 300986 122378 301222 122614
rect 301306 122378 301542 122614
rect 300986 122058 301222 122294
rect 301306 122058 301542 122294
rect 300986 86378 301222 86614
rect 301306 86378 301542 86614
rect 300986 86058 301222 86294
rect 301306 86058 301542 86294
rect 300986 50378 301222 50614
rect 301306 50378 301542 50614
rect 300986 50058 301222 50294
rect 301306 50058 301542 50294
rect 300986 14378 301222 14614
rect 301306 14378 301542 14614
rect 300986 14058 301222 14294
rect 301306 14058 301542 14294
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 307826 381218 308062 381454
rect 308146 381218 308382 381454
rect 307826 380898 308062 381134
rect 308146 380898 308382 381134
rect 307826 345218 308062 345454
rect 308146 345218 308382 345454
rect 307826 344898 308062 345134
rect 308146 344898 308382 345134
rect 307826 309218 308062 309454
rect 308146 309218 308382 309454
rect 307826 308898 308062 309134
rect 308146 308898 308382 309134
rect 307826 273218 308062 273454
rect 308146 273218 308382 273454
rect 307826 272898 308062 273134
rect 308146 272898 308382 273134
rect 307826 237218 308062 237454
rect 308146 237218 308382 237454
rect 307826 236898 308062 237134
rect 308146 236898 308382 237134
rect 307826 201218 308062 201454
rect 308146 201218 308382 201454
rect 307826 200898 308062 201134
rect 308146 200898 308382 201134
rect 307826 165218 308062 165454
rect 308146 165218 308382 165454
rect 307826 164898 308062 165134
rect 308146 164898 308382 165134
rect 307826 129218 308062 129454
rect 308146 129218 308382 129454
rect 307826 128898 308062 129134
rect 308146 128898 308382 129134
rect 307826 93218 308062 93454
rect 308146 93218 308382 93454
rect 307826 92898 308062 93134
rect 308146 92898 308382 93134
rect 307826 57218 308062 57454
rect 308146 57218 308382 57454
rect 307826 56898 308062 57134
rect 308146 56898 308382 57134
rect 307826 21218 308062 21454
rect 308146 21218 308382 21454
rect 307826 20898 308062 21134
rect 308146 20898 308382 21134
rect 307826 -1542 308062 -1306
rect 308146 -1542 308382 -1306
rect 307826 -1862 308062 -1626
rect 308146 -1862 308382 -1626
rect 311546 384938 311782 385174
rect 311866 384938 312102 385174
rect 311546 384618 311782 384854
rect 311866 384618 312102 384854
rect 311546 348938 311782 349174
rect 311866 348938 312102 349174
rect 311546 348618 311782 348854
rect 311866 348618 312102 348854
rect 311546 312938 311782 313174
rect 311866 312938 312102 313174
rect 311546 312618 311782 312854
rect 311866 312618 312102 312854
rect 311546 276938 311782 277174
rect 311866 276938 312102 277174
rect 311546 276618 311782 276854
rect 311866 276618 312102 276854
rect 311546 240938 311782 241174
rect 311866 240938 312102 241174
rect 311546 240618 311782 240854
rect 311866 240618 312102 240854
rect 311546 204938 311782 205174
rect 311866 204938 312102 205174
rect 311546 204618 311782 204854
rect 311866 204618 312102 204854
rect 311546 168938 311782 169174
rect 311866 168938 312102 169174
rect 311546 168618 311782 168854
rect 311866 168618 312102 168854
rect 311546 132938 311782 133174
rect 311866 132938 312102 133174
rect 311546 132618 311782 132854
rect 311866 132618 312102 132854
rect 311546 96938 311782 97174
rect 311866 96938 312102 97174
rect 311546 96618 311782 96854
rect 311866 96618 312102 96854
rect 311546 60938 311782 61174
rect 311866 60938 312102 61174
rect 311546 60618 311782 60854
rect 311866 60618 312102 60854
rect 311546 24938 311782 25174
rect 311866 24938 312102 25174
rect 311546 24618 311782 24854
rect 311866 24618 312102 24854
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 388658 315502 388894
rect 315586 388658 315822 388894
rect 315266 388338 315502 388574
rect 315586 388338 315822 388574
rect 315266 352658 315502 352894
rect 315586 352658 315822 352894
rect 315266 352338 315502 352574
rect 315586 352338 315822 352574
rect 315266 316658 315502 316894
rect 315586 316658 315822 316894
rect 315266 316338 315502 316574
rect 315586 316338 315822 316574
rect 315266 280658 315502 280894
rect 315586 280658 315822 280894
rect 315266 280338 315502 280574
rect 315586 280338 315822 280574
rect 315266 244658 315502 244894
rect 315586 244658 315822 244894
rect 315266 244338 315502 244574
rect 315586 244338 315822 244574
rect 315266 208658 315502 208894
rect 315586 208658 315822 208894
rect 315266 208338 315502 208574
rect 315586 208338 315822 208574
rect 315266 172658 315502 172894
rect 315586 172658 315822 172894
rect 315266 172338 315502 172574
rect 315586 172338 315822 172574
rect 315266 136658 315502 136894
rect 315586 136658 315822 136894
rect 315266 136338 315502 136574
rect 315586 136338 315822 136574
rect 315266 100658 315502 100894
rect 315586 100658 315822 100894
rect 315266 100338 315502 100574
rect 315586 100338 315822 100574
rect 315266 64658 315502 64894
rect 315586 64658 315822 64894
rect 315266 64338 315502 64574
rect 315586 64338 315822 64574
rect 315266 28658 315502 28894
rect 315586 28658 315822 28894
rect 315266 28338 315502 28574
rect 315586 28338 315822 28574
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 318986 392378 319222 392614
rect 319306 392378 319542 392614
rect 318986 392058 319222 392294
rect 319306 392058 319542 392294
rect 318986 356378 319222 356614
rect 319306 356378 319542 356614
rect 318986 356058 319222 356294
rect 319306 356058 319542 356294
rect 318986 320378 319222 320614
rect 319306 320378 319542 320614
rect 318986 320058 319222 320294
rect 319306 320058 319542 320294
rect 318986 284378 319222 284614
rect 319306 284378 319542 284614
rect 318986 284058 319222 284294
rect 319306 284058 319542 284294
rect 318986 248378 319222 248614
rect 319306 248378 319542 248614
rect 318986 248058 319222 248294
rect 319306 248058 319542 248294
rect 318986 212378 319222 212614
rect 319306 212378 319542 212614
rect 318986 212058 319222 212294
rect 319306 212058 319542 212294
rect 318986 176378 319222 176614
rect 319306 176378 319542 176614
rect 318986 176058 319222 176294
rect 319306 176058 319542 176294
rect 318986 140378 319222 140614
rect 319306 140378 319542 140614
rect 318986 140058 319222 140294
rect 319306 140058 319542 140294
rect 318986 104378 319222 104614
rect 319306 104378 319542 104614
rect 318986 104058 319222 104294
rect 319306 104058 319542 104294
rect 318986 68378 319222 68614
rect 319306 68378 319542 68614
rect 318986 68058 319222 68294
rect 319306 68058 319542 68294
rect 318986 32378 319222 32614
rect 319306 32378 319542 32614
rect 318986 32058 319222 32294
rect 319306 32058 319542 32294
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 325826 363218 326062 363454
rect 326146 363218 326382 363454
rect 325826 362898 326062 363134
rect 326146 362898 326382 363134
rect 325826 327218 326062 327454
rect 326146 327218 326382 327454
rect 325826 326898 326062 327134
rect 326146 326898 326382 327134
rect 325826 291218 326062 291454
rect 326146 291218 326382 291454
rect 325826 290898 326062 291134
rect 326146 290898 326382 291134
rect 325826 255218 326062 255454
rect 326146 255218 326382 255454
rect 325826 254898 326062 255134
rect 326146 254898 326382 255134
rect 325826 219218 326062 219454
rect 326146 219218 326382 219454
rect 325826 218898 326062 219134
rect 326146 218898 326382 219134
rect 325826 183218 326062 183454
rect 326146 183218 326382 183454
rect 325826 182898 326062 183134
rect 326146 182898 326382 183134
rect 325826 147218 326062 147454
rect 326146 147218 326382 147454
rect 325826 146898 326062 147134
rect 326146 146898 326382 147134
rect 325826 111218 326062 111454
rect 326146 111218 326382 111454
rect 325826 110898 326062 111134
rect 326146 110898 326382 111134
rect 325826 75218 326062 75454
rect 326146 75218 326382 75454
rect 325826 74898 326062 75134
rect 326146 74898 326382 75134
rect 325826 39218 326062 39454
rect 326146 39218 326382 39454
rect 325826 38898 326062 39134
rect 326146 38898 326382 39134
rect 325826 3218 326062 3454
rect 326146 3218 326382 3454
rect 325826 2898 326062 3134
rect 326146 2898 326382 3134
rect 325826 -582 326062 -346
rect 326146 -582 326382 -346
rect 325826 -902 326062 -666
rect 326146 -902 326382 -666
rect 329546 366938 329782 367174
rect 329866 366938 330102 367174
rect 329546 366618 329782 366854
rect 329866 366618 330102 366854
rect 329546 330938 329782 331174
rect 329866 330938 330102 331174
rect 329546 330618 329782 330854
rect 329866 330618 330102 330854
rect 329546 294938 329782 295174
rect 329866 294938 330102 295174
rect 329546 294618 329782 294854
rect 329866 294618 330102 294854
rect 329546 258938 329782 259174
rect 329866 258938 330102 259174
rect 329546 258618 329782 258854
rect 329866 258618 330102 258854
rect 329546 222938 329782 223174
rect 329866 222938 330102 223174
rect 329546 222618 329782 222854
rect 329866 222618 330102 222854
rect 329546 186938 329782 187174
rect 329866 186938 330102 187174
rect 329546 186618 329782 186854
rect 329866 186618 330102 186854
rect 329546 150938 329782 151174
rect 329866 150938 330102 151174
rect 329546 150618 329782 150854
rect 329866 150618 330102 150854
rect 329546 114938 329782 115174
rect 329866 114938 330102 115174
rect 329546 114618 329782 114854
rect 329866 114618 330102 114854
rect 329546 78938 329782 79174
rect 329866 78938 330102 79174
rect 329546 78618 329782 78854
rect 329866 78618 330102 78854
rect 329546 42938 329782 43174
rect 329866 42938 330102 43174
rect 329546 42618 329782 42854
rect 329866 42618 330102 42854
rect 329546 6938 329782 7174
rect 329866 6938 330102 7174
rect 329546 6618 329782 6854
rect 329866 6618 330102 6854
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 370658 333502 370894
rect 333586 370658 333822 370894
rect 333266 370338 333502 370574
rect 333586 370338 333822 370574
rect 333266 334658 333502 334894
rect 333586 334658 333822 334894
rect 333266 334338 333502 334574
rect 333586 334338 333822 334574
rect 333266 298658 333502 298894
rect 333586 298658 333822 298894
rect 333266 298338 333502 298574
rect 333586 298338 333822 298574
rect 333266 262658 333502 262894
rect 333586 262658 333822 262894
rect 333266 262338 333502 262574
rect 333586 262338 333822 262574
rect 333266 226658 333502 226894
rect 333586 226658 333822 226894
rect 333266 226338 333502 226574
rect 333586 226338 333822 226574
rect 333266 190658 333502 190894
rect 333586 190658 333822 190894
rect 333266 190338 333502 190574
rect 333586 190338 333822 190574
rect 333266 154658 333502 154894
rect 333586 154658 333822 154894
rect 333266 154338 333502 154574
rect 333586 154338 333822 154574
rect 333266 118658 333502 118894
rect 333586 118658 333822 118894
rect 333266 118338 333502 118574
rect 333586 118338 333822 118574
rect 333266 82658 333502 82894
rect 333586 82658 333822 82894
rect 333266 82338 333502 82574
rect 333586 82338 333822 82574
rect 333266 46658 333502 46894
rect 333586 46658 333822 46894
rect 333266 46338 333502 46574
rect 333586 46338 333822 46574
rect 333266 10658 333502 10894
rect 333586 10658 333822 10894
rect 333266 10338 333502 10574
rect 333586 10338 333822 10574
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 361826 399218 362062 399454
rect 362146 399218 362382 399454
rect 361826 398898 362062 399134
rect 362146 398898 362382 399134
rect 336986 374378 337222 374614
rect 337306 374378 337542 374614
rect 336986 374058 337222 374294
rect 337306 374058 337542 374294
rect 336986 338378 337222 338614
rect 337306 338378 337542 338614
rect 336986 338058 337222 338294
rect 337306 338058 337542 338294
rect 336986 302378 337222 302614
rect 337306 302378 337542 302614
rect 336986 302058 337222 302294
rect 337306 302058 337542 302294
rect 336986 266378 337222 266614
rect 337306 266378 337542 266614
rect 336986 266058 337222 266294
rect 337306 266058 337542 266294
rect 336986 230378 337222 230614
rect 337306 230378 337542 230614
rect 336986 230058 337222 230294
rect 337306 230058 337542 230294
rect 336986 194378 337222 194614
rect 337306 194378 337542 194614
rect 336986 194058 337222 194294
rect 337306 194058 337542 194294
rect 336986 158378 337222 158614
rect 337306 158378 337542 158614
rect 336986 158058 337222 158294
rect 337306 158058 337542 158294
rect 336986 122378 337222 122614
rect 337306 122378 337542 122614
rect 336986 122058 337222 122294
rect 337306 122058 337542 122294
rect 336986 86378 337222 86614
rect 337306 86378 337542 86614
rect 336986 86058 337222 86294
rect 337306 86058 337542 86294
rect 336986 50378 337222 50614
rect 337306 50378 337542 50614
rect 336986 50058 337222 50294
rect 337306 50058 337542 50294
rect 336986 14378 337222 14614
rect 337306 14378 337542 14614
rect 336986 14058 337222 14294
rect 337306 14058 337542 14294
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 343826 381218 344062 381454
rect 344146 381218 344382 381454
rect 343826 380898 344062 381134
rect 344146 380898 344382 381134
rect 343826 345218 344062 345454
rect 344146 345218 344382 345454
rect 343826 344898 344062 345134
rect 344146 344898 344382 345134
rect 343826 309218 344062 309454
rect 344146 309218 344382 309454
rect 343826 308898 344062 309134
rect 344146 308898 344382 309134
rect 343826 273218 344062 273454
rect 344146 273218 344382 273454
rect 343826 272898 344062 273134
rect 344146 272898 344382 273134
rect 343826 237218 344062 237454
rect 344146 237218 344382 237454
rect 343826 236898 344062 237134
rect 344146 236898 344382 237134
rect 343826 201218 344062 201454
rect 344146 201218 344382 201454
rect 343826 200898 344062 201134
rect 344146 200898 344382 201134
rect 343826 165218 344062 165454
rect 344146 165218 344382 165454
rect 343826 164898 344062 165134
rect 344146 164898 344382 165134
rect 343826 129218 344062 129454
rect 344146 129218 344382 129454
rect 343826 128898 344062 129134
rect 344146 128898 344382 129134
rect 343826 93218 344062 93454
rect 344146 93218 344382 93454
rect 343826 92898 344062 93134
rect 344146 92898 344382 93134
rect 343826 57218 344062 57454
rect 344146 57218 344382 57454
rect 343826 56898 344062 57134
rect 344146 56898 344382 57134
rect 343826 21218 344062 21454
rect 344146 21218 344382 21454
rect 343826 20898 344062 21134
rect 344146 20898 344382 21134
rect 343826 -1542 344062 -1306
rect 344146 -1542 344382 -1306
rect 343826 -1862 344062 -1626
rect 344146 -1862 344382 -1626
rect 347546 384938 347782 385174
rect 347866 384938 348102 385174
rect 347546 384618 347782 384854
rect 347866 384618 348102 384854
rect 347546 348938 347782 349174
rect 347866 348938 348102 349174
rect 347546 348618 347782 348854
rect 347866 348618 348102 348854
rect 347546 312938 347782 313174
rect 347866 312938 348102 313174
rect 347546 312618 347782 312854
rect 347866 312618 348102 312854
rect 347546 276938 347782 277174
rect 347866 276938 348102 277174
rect 347546 276618 347782 276854
rect 347866 276618 348102 276854
rect 347546 240938 347782 241174
rect 347866 240938 348102 241174
rect 347546 240618 347782 240854
rect 347866 240618 348102 240854
rect 347546 204938 347782 205174
rect 347866 204938 348102 205174
rect 347546 204618 347782 204854
rect 347866 204618 348102 204854
rect 347546 168938 347782 169174
rect 347866 168938 348102 169174
rect 347546 168618 347782 168854
rect 347866 168618 348102 168854
rect 347546 132938 347782 133174
rect 347866 132938 348102 133174
rect 347546 132618 347782 132854
rect 347866 132618 348102 132854
rect 347546 96938 347782 97174
rect 347866 96938 348102 97174
rect 347546 96618 347782 96854
rect 347866 96618 348102 96854
rect 347546 60938 347782 61174
rect 347866 60938 348102 61174
rect 347546 60618 347782 60854
rect 347866 60618 348102 60854
rect 347546 24938 347782 25174
rect 347866 24938 348102 25174
rect 347546 24618 347782 24854
rect 347866 24618 348102 24854
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 388658 351502 388894
rect 351586 388658 351822 388894
rect 351266 388338 351502 388574
rect 351586 388338 351822 388574
rect 351266 352658 351502 352894
rect 351586 352658 351822 352894
rect 351266 352338 351502 352574
rect 351586 352338 351822 352574
rect 351266 316658 351502 316894
rect 351586 316658 351822 316894
rect 351266 316338 351502 316574
rect 351586 316338 351822 316574
rect 351266 280658 351502 280894
rect 351586 280658 351822 280894
rect 351266 280338 351502 280574
rect 351586 280338 351822 280574
rect 351266 244658 351502 244894
rect 351586 244658 351822 244894
rect 351266 244338 351502 244574
rect 351586 244338 351822 244574
rect 351266 208658 351502 208894
rect 351586 208658 351822 208894
rect 351266 208338 351502 208574
rect 351586 208338 351822 208574
rect 351266 172658 351502 172894
rect 351586 172658 351822 172894
rect 351266 172338 351502 172574
rect 351586 172338 351822 172574
rect 351266 136658 351502 136894
rect 351586 136658 351822 136894
rect 351266 136338 351502 136574
rect 351586 136338 351822 136574
rect 351266 100658 351502 100894
rect 351586 100658 351822 100894
rect 351266 100338 351502 100574
rect 351586 100338 351822 100574
rect 351266 64658 351502 64894
rect 351586 64658 351822 64894
rect 351266 64338 351502 64574
rect 351586 64338 351822 64574
rect 351266 28658 351502 28894
rect 351586 28658 351822 28894
rect 351266 28338 351502 28574
rect 351586 28338 351822 28574
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 354986 392378 355222 392614
rect 355306 392378 355542 392614
rect 354986 392058 355222 392294
rect 355306 392058 355542 392294
rect 354986 356378 355222 356614
rect 355306 356378 355542 356614
rect 354986 356058 355222 356294
rect 355306 356058 355542 356294
rect 354986 320378 355222 320614
rect 355306 320378 355542 320614
rect 354986 320058 355222 320294
rect 355306 320058 355542 320294
rect 354986 284378 355222 284614
rect 355306 284378 355542 284614
rect 354986 284058 355222 284294
rect 355306 284058 355542 284294
rect 354986 248378 355222 248614
rect 355306 248378 355542 248614
rect 354986 248058 355222 248294
rect 355306 248058 355542 248294
rect 354986 212378 355222 212614
rect 355306 212378 355542 212614
rect 354986 212058 355222 212294
rect 355306 212058 355542 212294
rect 354986 176378 355222 176614
rect 355306 176378 355542 176614
rect 354986 176058 355222 176294
rect 355306 176058 355542 176294
rect 354986 140378 355222 140614
rect 355306 140378 355542 140614
rect 354986 140058 355222 140294
rect 355306 140058 355542 140294
rect 354986 104378 355222 104614
rect 355306 104378 355542 104614
rect 354986 104058 355222 104294
rect 355306 104058 355542 104294
rect 354986 68378 355222 68614
rect 355306 68378 355542 68614
rect 354986 68058 355222 68294
rect 355306 68058 355542 68294
rect 354986 32378 355222 32614
rect 355306 32378 355542 32614
rect 354986 32058 355222 32294
rect 355306 32058 355542 32294
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 361826 363218 362062 363454
rect 362146 363218 362382 363454
rect 361826 362898 362062 363134
rect 362146 362898 362382 363134
rect 361826 327218 362062 327454
rect 362146 327218 362382 327454
rect 361826 326898 362062 327134
rect 362146 326898 362382 327134
rect 361826 291218 362062 291454
rect 362146 291218 362382 291454
rect 361826 290898 362062 291134
rect 362146 290898 362382 291134
rect 361826 255218 362062 255454
rect 362146 255218 362382 255454
rect 361826 254898 362062 255134
rect 362146 254898 362382 255134
rect 361826 219218 362062 219454
rect 362146 219218 362382 219454
rect 361826 218898 362062 219134
rect 362146 218898 362382 219134
rect 361826 183218 362062 183454
rect 362146 183218 362382 183454
rect 361826 182898 362062 183134
rect 362146 182898 362382 183134
rect 361826 147218 362062 147454
rect 362146 147218 362382 147454
rect 361826 146898 362062 147134
rect 362146 146898 362382 147134
rect 361826 111218 362062 111454
rect 362146 111218 362382 111454
rect 361826 110898 362062 111134
rect 362146 110898 362382 111134
rect 361826 75218 362062 75454
rect 362146 75218 362382 75454
rect 361826 74898 362062 75134
rect 362146 74898 362382 75134
rect 361826 39218 362062 39454
rect 362146 39218 362382 39454
rect 361826 38898 362062 39134
rect 362146 38898 362382 39134
rect 361826 3218 362062 3454
rect 362146 3218 362382 3454
rect 361826 2898 362062 3134
rect 362146 2898 362382 3134
rect 361826 -582 362062 -346
rect 362146 -582 362382 -346
rect 361826 -902 362062 -666
rect 362146 -902 362382 -666
rect 365546 690938 365782 691174
rect 365866 690938 366102 691174
rect 365546 690618 365782 690854
rect 365866 690618 366102 690854
rect 365546 654938 365782 655174
rect 365866 654938 366102 655174
rect 365546 654618 365782 654854
rect 365866 654618 366102 654854
rect 365546 618938 365782 619174
rect 365866 618938 366102 619174
rect 365546 618618 365782 618854
rect 365866 618618 366102 618854
rect 365546 582938 365782 583174
rect 365866 582938 366102 583174
rect 365546 582618 365782 582854
rect 365866 582618 366102 582854
rect 365546 546938 365782 547174
rect 365866 546938 366102 547174
rect 365546 546618 365782 546854
rect 365866 546618 366102 546854
rect 365546 510938 365782 511174
rect 365866 510938 366102 511174
rect 365546 510618 365782 510854
rect 365866 510618 366102 510854
rect 365546 474938 365782 475174
rect 365866 474938 366102 475174
rect 365546 474618 365782 474854
rect 365866 474618 366102 474854
rect 365546 438938 365782 439174
rect 365866 438938 366102 439174
rect 365546 438618 365782 438854
rect 365866 438618 366102 438854
rect 365546 402938 365782 403174
rect 365866 402938 366102 403174
rect 365546 402618 365782 402854
rect 365866 402618 366102 402854
rect 365546 366938 365782 367174
rect 365866 366938 366102 367174
rect 365546 366618 365782 366854
rect 365866 366618 366102 366854
rect 365546 330938 365782 331174
rect 365866 330938 366102 331174
rect 365546 330618 365782 330854
rect 365866 330618 366102 330854
rect 365546 294938 365782 295174
rect 365866 294938 366102 295174
rect 365546 294618 365782 294854
rect 365866 294618 366102 294854
rect 365546 258938 365782 259174
rect 365866 258938 366102 259174
rect 365546 258618 365782 258854
rect 365866 258618 366102 258854
rect 365546 222938 365782 223174
rect 365866 222938 366102 223174
rect 365546 222618 365782 222854
rect 365866 222618 366102 222854
rect 365546 186938 365782 187174
rect 365866 186938 366102 187174
rect 365546 186618 365782 186854
rect 365866 186618 366102 186854
rect 365546 150938 365782 151174
rect 365866 150938 366102 151174
rect 365546 150618 365782 150854
rect 365866 150618 366102 150854
rect 365546 114938 365782 115174
rect 365866 114938 366102 115174
rect 365546 114618 365782 114854
rect 365866 114618 366102 114854
rect 365546 78938 365782 79174
rect 365866 78938 366102 79174
rect 365546 78618 365782 78854
rect 365866 78618 366102 78854
rect 365546 42938 365782 43174
rect 365866 42938 366102 43174
rect 365546 42618 365782 42854
rect 365866 42618 366102 42854
rect 365546 6938 365782 7174
rect 365866 6938 366102 7174
rect 365546 6618 365782 6854
rect 365866 6618 366102 6854
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 694658 369502 694894
rect 369586 694658 369822 694894
rect 369266 694338 369502 694574
rect 369586 694338 369822 694574
rect 369266 658658 369502 658894
rect 369586 658658 369822 658894
rect 369266 658338 369502 658574
rect 369586 658338 369822 658574
rect 369266 622658 369502 622894
rect 369586 622658 369822 622894
rect 369266 622338 369502 622574
rect 369586 622338 369822 622574
rect 369266 586658 369502 586894
rect 369586 586658 369822 586894
rect 369266 586338 369502 586574
rect 369586 586338 369822 586574
rect 369266 550658 369502 550894
rect 369586 550658 369822 550894
rect 369266 550338 369502 550574
rect 369586 550338 369822 550574
rect 369266 514658 369502 514894
rect 369586 514658 369822 514894
rect 369266 514338 369502 514574
rect 369586 514338 369822 514574
rect 369266 478658 369502 478894
rect 369586 478658 369822 478894
rect 369266 478338 369502 478574
rect 369586 478338 369822 478574
rect 369266 442658 369502 442894
rect 369586 442658 369822 442894
rect 369266 442338 369502 442574
rect 369586 442338 369822 442574
rect 369266 406658 369502 406894
rect 369586 406658 369822 406894
rect 369266 406338 369502 406574
rect 369586 406338 369822 406574
rect 369266 370658 369502 370894
rect 369586 370658 369822 370894
rect 369266 370338 369502 370574
rect 369586 370338 369822 370574
rect 369266 334658 369502 334894
rect 369586 334658 369822 334894
rect 369266 334338 369502 334574
rect 369586 334338 369822 334574
rect 369266 298658 369502 298894
rect 369586 298658 369822 298894
rect 369266 298338 369502 298574
rect 369586 298338 369822 298574
rect 369266 262658 369502 262894
rect 369586 262658 369822 262894
rect 369266 262338 369502 262574
rect 369586 262338 369822 262574
rect 369266 226658 369502 226894
rect 369586 226658 369822 226894
rect 369266 226338 369502 226574
rect 369586 226338 369822 226574
rect 369266 190658 369502 190894
rect 369586 190658 369822 190894
rect 369266 190338 369502 190574
rect 369586 190338 369822 190574
rect 369266 154658 369502 154894
rect 369586 154658 369822 154894
rect 369266 154338 369502 154574
rect 369586 154338 369822 154574
rect 369266 118658 369502 118894
rect 369586 118658 369822 118894
rect 369266 118338 369502 118574
rect 369586 118338 369822 118574
rect 369266 82658 369502 82894
rect 369586 82658 369822 82894
rect 369266 82338 369502 82574
rect 369586 82338 369822 82574
rect 369266 46658 369502 46894
rect 369586 46658 369822 46894
rect 369266 46338 369502 46574
rect 369586 46338 369822 46574
rect 369266 10658 369502 10894
rect 369586 10658 369822 10894
rect 369266 10338 369502 10574
rect 369586 10338 369822 10574
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 372986 698378 373222 698614
rect 373306 698378 373542 698614
rect 372986 698058 373222 698294
rect 373306 698058 373542 698294
rect 372986 662378 373222 662614
rect 373306 662378 373542 662614
rect 372986 662058 373222 662294
rect 373306 662058 373542 662294
rect 372986 626378 373222 626614
rect 373306 626378 373542 626614
rect 372986 626058 373222 626294
rect 373306 626058 373542 626294
rect 372986 590378 373222 590614
rect 373306 590378 373542 590614
rect 372986 590058 373222 590294
rect 373306 590058 373542 590294
rect 372986 554378 373222 554614
rect 373306 554378 373542 554614
rect 372986 554058 373222 554294
rect 373306 554058 373542 554294
rect 372986 518378 373222 518614
rect 373306 518378 373542 518614
rect 372986 518058 373222 518294
rect 373306 518058 373542 518294
rect 372986 482378 373222 482614
rect 373306 482378 373542 482614
rect 372986 482058 373222 482294
rect 373306 482058 373542 482294
rect 372986 446378 373222 446614
rect 373306 446378 373542 446614
rect 372986 446058 373222 446294
rect 373306 446058 373542 446294
rect 372986 410378 373222 410614
rect 373306 410378 373542 410614
rect 372986 410058 373222 410294
rect 373306 410058 373542 410294
rect 372986 374378 373222 374614
rect 373306 374378 373542 374614
rect 372986 374058 373222 374294
rect 373306 374058 373542 374294
rect 372986 338378 373222 338614
rect 373306 338378 373542 338614
rect 372986 338058 373222 338294
rect 373306 338058 373542 338294
rect 372986 302378 373222 302614
rect 373306 302378 373542 302614
rect 372986 302058 373222 302294
rect 373306 302058 373542 302294
rect 372986 266378 373222 266614
rect 373306 266378 373542 266614
rect 372986 266058 373222 266294
rect 373306 266058 373542 266294
rect 372986 230378 373222 230614
rect 373306 230378 373542 230614
rect 372986 230058 373222 230294
rect 373306 230058 373542 230294
rect 372986 194378 373222 194614
rect 373306 194378 373542 194614
rect 372986 194058 373222 194294
rect 373306 194058 373542 194294
rect 372986 158378 373222 158614
rect 373306 158378 373542 158614
rect 372986 158058 373222 158294
rect 373306 158058 373542 158294
rect 372986 122378 373222 122614
rect 373306 122378 373542 122614
rect 372986 122058 373222 122294
rect 373306 122058 373542 122294
rect 372986 86378 373222 86614
rect 373306 86378 373542 86614
rect 372986 86058 373222 86294
rect 373306 86058 373542 86294
rect 372986 50378 373222 50614
rect 373306 50378 373542 50614
rect 372986 50058 373222 50294
rect 373306 50058 373542 50294
rect 372986 14378 373222 14614
rect 373306 14378 373542 14614
rect 372986 14058 373222 14294
rect 373306 14058 373542 14294
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 379826 669218 380062 669454
rect 380146 669218 380382 669454
rect 379826 668898 380062 669134
rect 380146 668898 380382 669134
rect 379826 633218 380062 633454
rect 380146 633218 380382 633454
rect 379826 632898 380062 633134
rect 380146 632898 380382 633134
rect 379826 597218 380062 597454
rect 380146 597218 380382 597454
rect 379826 596898 380062 597134
rect 380146 596898 380382 597134
rect 379826 561218 380062 561454
rect 380146 561218 380382 561454
rect 379826 560898 380062 561134
rect 380146 560898 380382 561134
rect 379826 525218 380062 525454
rect 380146 525218 380382 525454
rect 379826 524898 380062 525134
rect 380146 524898 380382 525134
rect 379826 489218 380062 489454
rect 380146 489218 380382 489454
rect 379826 488898 380062 489134
rect 380146 488898 380382 489134
rect 379826 453218 380062 453454
rect 380146 453218 380382 453454
rect 379826 452898 380062 453134
rect 380146 452898 380382 453134
rect 379826 417218 380062 417454
rect 380146 417218 380382 417454
rect 379826 416898 380062 417134
rect 380146 416898 380382 417134
rect 379826 381218 380062 381454
rect 380146 381218 380382 381454
rect 379826 380898 380062 381134
rect 380146 380898 380382 381134
rect 379826 345218 380062 345454
rect 380146 345218 380382 345454
rect 379826 344898 380062 345134
rect 380146 344898 380382 345134
rect 379826 309218 380062 309454
rect 380146 309218 380382 309454
rect 379826 308898 380062 309134
rect 380146 308898 380382 309134
rect 379826 273218 380062 273454
rect 380146 273218 380382 273454
rect 379826 272898 380062 273134
rect 380146 272898 380382 273134
rect 379826 237218 380062 237454
rect 380146 237218 380382 237454
rect 379826 236898 380062 237134
rect 380146 236898 380382 237134
rect 379826 201218 380062 201454
rect 380146 201218 380382 201454
rect 379826 200898 380062 201134
rect 380146 200898 380382 201134
rect 379826 165218 380062 165454
rect 380146 165218 380382 165454
rect 379826 164898 380062 165134
rect 380146 164898 380382 165134
rect 379826 129218 380062 129454
rect 380146 129218 380382 129454
rect 379826 128898 380062 129134
rect 380146 128898 380382 129134
rect 379826 93218 380062 93454
rect 380146 93218 380382 93454
rect 379826 92898 380062 93134
rect 380146 92898 380382 93134
rect 379826 57218 380062 57454
rect 380146 57218 380382 57454
rect 379826 56898 380062 57134
rect 380146 56898 380382 57134
rect 379826 21218 380062 21454
rect 380146 21218 380382 21454
rect 379826 20898 380062 21134
rect 380146 20898 380382 21134
rect 379826 -1542 380062 -1306
rect 380146 -1542 380382 -1306
rect 379826 -1862 380062 -1626
rect 380146 -1862 380382 -1626
rect 383546 672938 383782 673174
rect 383866 672938 384102 673174
rect 383546 672618 383782 672854
rect 383866 672618 384102 672854
rect 383546 636938 383782 637174
rect 383866 636938 384102 637174
rect 383546 636618 383782 636854
rect 383866 636618 384102 636854
rect 383546 600938 383782 601174
rect 383866 600938 384102 601174
rect 383546 600618 383782 600854
rect 383866 600618 384102 600854
rect 383546 564938 383782 565174
rect 383866 564938 384102 565174
rect 383546 564618 383782 564854
rect 383866 564618 384102 564854
rect 383546 528938 383782 529174
rect 383866 528938 384102 529174
rect 383546 528618 383782 528854
rect 383866 528618 384102 528854
rect 383546 492938 383782 493174
rect 383866 492938 384102 493174
rect 383546 492618 383782 492854
rect 383866 492618 384102 492854
rect 383546 456938 383782 457174
rect 383866 456938 384102 457174
rect 383546 456618 383782 456854
rect 383866 456618 384102 456854
rect 383546 420938 383782 421174
rect 383866 420938 384102 421174
rect 383546 420618 383782 420854
rect 383866 420618 384102 420854
rect 383546 384938 383782 385174
rect 383866 384938 384102 385174
rect 383546 384618 383782 384854
rect 383866 384618 384102 384854
rect 383546 348938 383782 349174
rect 383866 348938 384102 349174
rect 383546 348618 383782 348854
rect 383866 348618 384102 348854
rect 383546 312938 383782 313174
rect 383866 312938 384102 313174
rect 383546 312618 383782 312854
rect 383866 312618 384102 312854
rect 383546 276938 383782 277174
rect 383866 276938 384102 277174
rect 383546 276618 383782 276854
rect 383866 276618 384102 276854
rect 383546 240938 383782 241174
rect 383866 240938 384102 241174
rect 383546 240618 383782 240854
rect 383866 240618 384102 240854
rect 383546 204938 383782 205174
rect 383866 204938 384102 205174
rect 383546 204618 383782 204854
rect 383866 204618 384102 204854
rect 383546 168938 383782 169174
rect 383866 168938 384102 169174
rect 383546 168618 383782 168854
rect 383866 168618 384102 168854
rect 383546 132938 383782 133174
rect 383866 132938 384102 133174
rect 383546 132618 383782 132854
rect 383866 132618 384102 132854
rect 383546 96938 383782 97174
rect 383866 96938 384102 97174
rect 383546 96618 383782 96854
rect 383866 96618 384102 96854
rect 383546 60938 383782 61174
rect 383866 60938 384102 61174
rect 383546 60618 383782 60854
rect 383866 60618 384102 60854
rect 383546 24938 383782 25174
rect 383866 24938 384102 25174
rect 383546 24618 383782 24854
rect 383866 24618 384102 24854
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 676658 387502 676894
rect 387586 676658 387822 676894
rect 387266 676338 387502 676574
rect 387586 676338 387822 676574
rect 387266 640658 387502 640894
rect 387586 640658 387822 640894
rect 387266 640338 387502 640574
rect 387586 640338 387822 640574
rect 387266 604658 387502 604894
rect 387586 604658 387822 604894
rect 387266 604338 387502 604574
rect 387586 604338 387822 604574
rect 387266 568658 387502 568894
rect 387586 568658 387822 568894
rect 387266 568338 387502 568574
rect 387586 568338 387822 568574
rect 387266 532658 387502 532894
rect 387586 532658 387822 532894
rect 387266 532338 387502 532574
rect 387586 532338 387822 532574
rect 387266 496658 387502 496894
rect 387586 496658 387822 496894
rect 387266 496338 387502 496574
rect 387586 496338 387822 496574
rect 387266 460658 387502 460894
rect 387586 460658 387822 460894
rect 387266 460338 387502 460574
rect 387586 460338 387822 460574
rect 387266 424658 387502 424894
rect 387586 424658 387822 424894
rect 387266 424338 387502 424574
rect 387586 424338 387822 424574
rect 387266 388658 387502 388894
rect 387586 388658 387822 388894
rect 387266 388338 387502 388574
rect 387586 388338 387822 388574
rect 387266 352658 387502 352894
rect 387586 352658 387822 352894
rect 387266 352338 387502 352574
rect 387586 352338 387822 352574
rect 387266 316658 387502 316894
rect 387586 316658 387822 316894
rect 387266 316338 387502 316574
rect 387586 316338 387822 316574
rect 387266 280658 387502 280894
rect 387586 280658 387822 280894
rect 387266 280338 387502 280574
rect 387586 280338 387822 280574
rect 387266 244658 387502 244894
rect 387586 244658 387822 244894
rect 387266 244338 387502 244574
rect 387586 244338 387822 244574
rect 387266 208658 387502 208894
rect 387586 208658 387822 208894
rect 387266 208338 387502 208574
rect 387586 208338 387822 208574
rect 387266 172658 387502 172894
rect 387586 172658 387822 172894
rect 387266 172338 387502 172574
rect 387586 172338 387822 172574
rect 387266 136658 387502 136894
rect 387586 136658 387822 136894
rect 387266 136338 387502 136574
rect 387586 136338 387822 136574
rect 387266 100658 387502 100894
rect 387586 100658 387822 100894
rect 387266 100338 387502 100574
rect 387586 100338 387822 100574
rect 387266 64658 387502 64894
rect 387586 64658 387822 64894
rect 387266 64338 387502 64574
rect 387586 64338 387822 64574
rect 387266 28658 387502 28894
rect 387586 28658 387822 28894
rect 387266 28338 387502 28574
rect 387586 28338 387822 28574
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 390986 680378 391222 680614
rect 391306 680378 391542 680614
rect 390986 680058 391222 680294
rect 391306 680058 391542 680294
rect 390986 644378 391222 644614
rect 391306 644378 391542 644614
rect 390986 644058 391222 644294
rect 391306 644058 391542 644294
rect 390986 608378 391222 608614
rect 391306 608378 391542 608614
rect 390986 608058 391222 608294
rect 391306 608058 391542 608294
rect 390986 572378 391222 572614
rect 391306 572378 391542 572614
rect 390986 572058 391222 572294
rect 391306 572058 391542 572294
rect 390986 536378 391222 536614
rect 391306 536378 391542 536614
rect 390986 536058 391222 536294
rect 391306 536058 391542 536294
rect 390986 500378 391222 500614
rect 391306 500378 391542 500614
rect 390986 500058 391222 500294
rect 391306 500058 391542 500294
rect 390986 464378 391222 464614
rect 391306 464378 391542 464614
rect 390986 464058 391222 464294
rect 391306 464058 391542 464294
rect 390986 428378 391222 428614
rect 391306 428378 391542 428614
rect 390986 428058 391222 428294
rect 391306 428058 391542 428294
rect 390986 392378 391222 392614
rect 391306 392378 391542 392614
rect 390986 392058 391222 392294
rect 391306 392058 391542 392294
rect 390986 356378 391222 356614
rect 391306 356378 391542 356614
rect 390986 356058 391222 356294
rect 391306 356058 391542 356294
rect 390986 320378 391222 320614
rect 391306 320378 391542 320614
rect 390986 320058 391222 320294
rect 391306 320058 391542 320294
rect 390986 284378 391222 284614
rect 391306 284378 391542 284614
rect 390986 284058 391222 284294
rect 391306 284058 391542 284294
rect 390986 248378 391222 248614
rect 391306 248378 391542 248614
rect 390986 248058 391222 248294
rect 391306 248058 391542 248294
rect 390986 212378 391222 212614
rect 391306 212378 391542 212614
rect 390986 212058 391222 212294
rect 391306 212058 391542 212294
rect 390986 176378 391222 176614
rect 391306 176378 391542 176614
rect 390986 176058 391222 176294
rect 391306 176058 391542 176294
rect 390986 140378 391222 140614
rect 391306 140378 391542 140614
rect 390986 140058 391222 140294
rect 391306 140058 391542 140294
rect 390986 104378 391222 104614
rect 391306 104378 391542 104614
rect 390986 104058 391222 104294
rect 391306 104058 391542 104294
rect 390986 68378 391222 68614
rect 391306 68378 391542 68614
rect 390986 68058 391222 68294
rect 391306 68058 391542 68294
rect 390986 32378 391222 32614
rect 391306 32378 391542 32614
rect 390986 32058 391222 32294
rect 391306 32058 391542 32294
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 397826 687218 398062 687454
rect 398146 687218 398382 687454
rect 397826 686898 398062 687134
rect 398146 686898 398382 687134
rect 397826 651218 398062 651454
rect 398146 651218 398382 651454
rect 397826 650898 398062 651134
rect 398146 650898 398382 651134
rect 397826 615218 398062 615454
rect 398146 615218 398382 615454
rect 397826 614898 398062 615134
rect 398146 614898 398382 615134
rect 397826 579218 398062 579454
rect 398146 579218 398382 579454
rect 397826 578898 398062 579134
rect 398146 578898 398382 579134
rect 397826 543218 398062 543454
rect 398146 543218 398382 543454
rect 397826 542898 398062 543134
rect 398146 542898 398382 543134
rect 397826 507218 398062 507454
rect 398146 507218 398382 507454
rect 397826 506898 398062 507134
rect 398146 506898 398382 507134
rect 397826 471218 398062 471454
rect 398146 471218 398382 471454
rect 397826 470898 398062 471134
rect 398146 470898 398382 471134
rect 397826 435218 398062 435454
rect 398146 435218 398382 435454
rect 397826 434898 398062 435134
rect 398146 434898 398382 435134
rect 397826 399218 398062 399454
rect 398146 399218 398382 399454
rect 397826 398898 398062 399134
rect 398146 398898 398382 399134
rect 397826 363218 398062 363454
rect 398146 363218 398382 363454
rect 397826 362898 398062 363134
rect 398146 362898 398382 363134
rect 397826 327218 398062 327454
rect 398146 327218 398382 327454
rect 397826 326898 398062 327134
rect 398146 326898 398382 327134
rect 397826 291218 398062 291454
rect 398146 291218 398382 291454
rect 397826 290898 398062 291134
rect 398146 290898 398382 291134
rect 397826 255218 398062 255454
rect 398146 255218 398382 255454
rect 397826 254898 398062 255134
rect 398146 254898 398382 255134
rect 397826 219218 398062 219454
rect 398146 219218 398382 219454
rect 397826 218898 398062 219134
rect 398146 218898 398382 219134
rect 397826 183218 398062 183454
rect 398146 183218 398382 183454
rect 397826 182898 398062 183134
rect 398146 182898 398382 183134
rect 397826 147218 398062 147454
rect 398146 147218 398382 147454
rect 397826 146898 398062 147134
rect 398146 146898 398382 147134
rect 397826 111218 398062 111454
rect 398146 111218 398382 111454
rect 397826 110898 398062 111134
rect 398146 110898 398382 111134
rect 397826 75218 398062 75454
rect 398146 75218 398382 75454
rect 397826 74898 398062 75134
rect 398146 74898 398382 75134
rect 397826 39218 398062 39454
rect 398146 39218 398382 39454
rect 397826 38898 398062 39134
rect 398146 38898 398382 39134
rect 397826 3218 398062 3454
rect 398146 3218 398382 3454
rect 397826 2898 398062 3134
rect 398146 2898 398382 3134
rect 397826 -582 398062 -346
rect 398146 -582 398382 -346
rect 397826 -902 398062 -666
rect 398146 -902 398382 -666
rect 401546 690938 401782 691174
rect 401866 690938 402102 691174
rect 401546 690618 401782 690854
rect 401866 690618 402102 690854
rect 401546 654938 401782 655174
rect 401866 654938 402102 655174
rect 401546 654618 401782 654854
rect 401866 654618 402102 654854
rect 401546 618938 401782 619174
rect 401866 618938 402102 619174
rect 401546 618618 401782 618854
rect 401866 618618 402102 618854
rect 401546 582938 401782 583174
rect 401866 582938 402102 583174
rect 401546 582618 401782 582854
rect 401866 582618 402102 582854
rect 401546 546938 401782 547174
rect 401866 546938 402102 547174
rect 401546 546618 401782 546854
rect 401866 546618 402102 546854
rect 401546 510938 401782 511174
rect 401866 510938 402102 511174
rect 401546 510618 401782 510854
rect 401866 510618 402102 510854
rect 401546 474938 401782 475174
rect 401866 474938 402102 475174
rect 401546 474618 401782 474854
rect 401866 474618 402102 474854
rect 401546 438938 401782 439174
rect 401866 438938 402102 439174
rect 401546 438618 401782 438854
rect 401866 438618 402102 438854
rect 401546 402938 401782 403174
rect 401866 402938 402102 403174
rect 401546 402618 401782 402854
rect 401866 402618 402102 402854
rect 401546 366938 401782 367174
rect 401866 366938 402102 367174
rect 401546 366618 401782 366854
rect 401866 366618 402102 366854
rect 401546 330938 401782 331174
rect 401866 330938 402102 331174
rect 401546 330618 401782 330854
rect 401866 330618 402102 330854
rect 401546 294938 401782 295174
rect 401866 294938 402102 295174
rect 401546 294618 401782 294854
rect 401866 294618 402102 294854
rect 401546 258938 401782 259174
rect 401866 258938 402102 259174
rect 401546 258618 401782 258854
rect 401866 258618 402102 258854
rect 401546 222938 401782 223174
rect 401866 222938 402102 223174
rect 401546 222618 401782 222854
rect 401866 222618 402102 222854
rect 401546 186938 401782 187174
rect 401866 186938 402102 187174
rect 401546 186618 401782 186854
rect 401866 186618 402102 186854
rect 401546 150938 401782 151174
rect 401866 150938 402102 151174
rect 401546 150618 401782 150854
rect 401866 150618 402102 150854
rect 401546 114938 401782 115174
rect 401866 114938 402102 115174
rect 401546 114618 401782 114854
rect 401866 114618 402102 114854
rect 401546 78938 401782 79174
rect 401866 78938 402102 79174
rect 401546 78618 401782 78854
rect 401866 78618 402102 78854
rect 401546 42938 401782 43174
rect 401866 42938 402102 43174
rect 401546 42618 401782 42854
rect 401866 42618 402102 42854
rect 401546 6938 401782 7174
rect 401866 6938 402102 7174
rect 401546 6618 401782 6854
rect 401866 6618 402102 6854
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 694658 405502 694894
rect 405586 694658 405822 694894
rect 405266 694338 405502 694574
rect 405586 694338 405822 694574
rect 405266 658658 405502 658894
rect 405586 658658 405822 658894
rect 405266 658338 405502 658574
rect 405586 658338 405822 658574
rect 405266 622658 405502 622894
rect 405586 622658 405822 622894
rect 405266 622338 405502 622574
rect 405586 622338 405822 622574
rect 405266 586658 405502 586894
rect 405586 586658 405822 586894
rect 405266 586338 405502 586574
rect 405586 586338 405822 586574
rect 405266 550658 405502 550894
rect 405586 550658 405822 550894
rect 405266 550338 405502 550574
rect 405586 550338 405822 550574
rect 405266 514658 405502 514894
rect 405586 514658 405822 514894
rect 405266 514338 405502 514574
rect 405586 514338 405822 514574
rect 405266 478658 405502 478894
rect 405586 478658 405822 478894
rect 405266 478338 405502 478574
rect 405586 478338 405822 478574
rect 405266 442658 405502 442894
rect 405586 442658 405822 442894
rect 405266 442338 405502 442574
rect 405586 442338 405822 442574
rect 405266 406658 405502 406894
rect 405586 406658 405822 406894
rect 405266 406338 405502 406574
rect 405586 406338 405822 406574
rect 405266 370658 405502 370894
rect 405586 370658 405822 370894
rect 405266 370338 405502 370574
rect 405586 370338 405822 370574
rect 405266 334658 405502 334894
rect 405586 334658 405822 334894
rect 405266 334338 405502 334574
rect 405586 334338 405822 334574
rect 405266 298658 405502 298894
rect 405586 298658 405822 298894
rect 405266 298338 405502 298574
rect 405586 298338 405822 298574
rect 405266 262658 405502 262894
rect 405586 262658 405822 262894
rect 405266 262338 405502 262574
rect 405586 262338 405822 262574
rect 405266 226658 405502 226894
rect 405586 226658 405822 226894
rect 405266 226338 405502 226574
rect 405586 226338 405822 226574
rect 405266 190658 405502 190894
rect 405586 190658 405822 190894
rect 405266 190338 405502 190574
rect 405586 190338 405822 190574
rect 405266 154658 405502 154894
rect 405586 154658 405822 154894
rect 405266 154338 405502 154574
rect 405586 154338 405822 154574
rect 405266 118658 405502 118894
rect 405586 118658 405822 118894
rect 405266 118338 405502 118574
rect 405586 118338 405822 118574
rect 405266 82658 405502 82894
rect 405586 82658 405822 82894
rect 405266 82338 405502 82574
rect 405586 82338 405822 82574
rect 405266 46658 405502 46894
rect 405586 46658 405822 46894
rect 405266 46338 405502 46574
rect 405586 46338 405822 46574
rect 405266 10658 405502 10894
rect 405586 10658 405822 10894
rect 405266 10338 405502 10574
rect 405586 10338 405822 10574
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 408986 698378 409222 698614
rect 409306 698378 409542 698614
rect 408986 698058 409222 698294
rect 409306 698058 409542 698294
rect 408986 662378 409222 662614
rect 409306 662378 409542 662614
rect 408986 662058 409222 662294
rect 409306 662058 409542 662294
rect 408986 626378 409222 626614
rect 409306 626378 409542 626614
rect 408986 626058 409222 626294
rect 409306 626058 409542 626294
rect 408986 590378 409222 590614
rect 409306 590378 409542 590614
rect 408986 590058 409222 590294
rect 409306 590058 409542 590294
rect 408986 554378 409222 554614
rect 409306 554378 409542 554614
rect 408986 554058 409222 554294
rect 409306 554058 409542 554294
rect 408986 518378 409222 518614
rect 409306 518378 409542 518614
rect 408986 518058 409222 518294
rect 409306 518058 409542 518294
rect 408986 482378 409222 482614
rect 409306 482378 409542 482614
rect 408986 482058 409222 482294
rect 409306 482058 409542 482294
rect 408986 446378 409222 446614
rect 409306 446378 409542 446614
rect 408986 446058 409222 446294
rect 409306 446058 409542 446294
rect 408986 410378 409222 410614
rect 409306 410378 409542 410614
rect 408986 410058 409222 410294
rect 409306 410058 409542 410294
rect 408986 374378 409222 374614
rect 409306 374378 409542 374614
rect 408986 374058 409222 374294
rect 409306 374058 409542 374294
rect 408986 338378 409222 338614
rect 409306 338378 409542 338614
rect 408986 338058 409222 338294
rect 409306 338058 409542 338294
rect 408986 302378 409222 302614
rect 409306 302378 409542 302614
rect 408986 302058 409222 302294
rect 409306 302058 409542 302294
rect 408986 266378 409222 266614
rect 409306 266378 409542 266614
rect 408986 266058 409222 266294
rect 409306 266058 409542 266294
rect 408986 230378 409222 230614
rect 409306 230378 409542 230614
rect 408986 230058 409222 230294
rect 409306 230058 409542 230294
rect 408986 194378 409222 194614
rect 409306 194378 409542 194614
rect 408986 194058 409222 194294
rect 409306 194058 409542 194294
rect 408986 158378 409222 158614
rect 409306 158378 409542 158614
rect 408986 158058 409222 158294
rect 409306 158058 409542 158294
rect 408986 122378 409222 122614
rect 409306 122378 409542 122614
rect 408986 122058 409222 122294
rect 409306 122058 409542 122294
rect 408986 86378 409222 86614
rect 409306 86378 409542 86614
rect 408986 86058 409222 86294
rect 409306 86058 409542 86294
rect 408986 50378 409222 50614
rect 409306 50378 409542 50614
rect 408986 50058 409222 50294
rect 409306 50058 409542 50294
rect 408986 14378 409222 14614
rect 409306 14378 409542 14614
rect 408986 14058 409222 14294
rect 409306 14058 409542 14294
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 415826 669218 416062 669454
rect 416146 669218 416382 669454
rect 415826 668898 416062 669134
rect 416146 668898 416382 669134
rect 415826 633218 416062 633454
rect 416146 633218 416382 633454
rect 415826 632898 416062 633134
rect 416146 632898 416382 633134
rect 415826 597218 416062 597454
rect 416146 597218 416382 597454
rect 415826 596898 416062 597134
rect 416146 596898 416382 597134
rect 415826 561218 416062 561454
rect 416146 561218 416382 561454
rect 415826 560898 416062 561134
rect 416146 560898 416382 561134
rect 415826 525218 416062 525454
rect 416146 525218 416382 525454
rect 415826 524898 416062 525134
rect 416146 524898 416382 525134
rect 415826 489218 416062 489454
rect 416146 489218 416382 489454
rect 415826 488898 416062 489134
rect 416146 488898 416382 489134
rect 415826 453218 416062 453454
rect 416146 453218 416382 453454
rect 415826 452898 416062 453134
rect 416146 452898 416382 453134
rect 415826 417218 416062 417454
rect 416146 417218 416382 417454
rect 415826 416898 416062 417134
rect 416146 416898 416382 417134
rect 415826 381218 416062 381454
rect 416146 381218 416382 381454
rect 415826 380898 416062 381134
rect 416146 380898 416382 381134
rect 415826 345218 416062 345454
rect 416146 345218 416382 345454
rect 415826 344898 416062 345134
rect 416146 344898 416382 345134
rect 415826 309218 416062 309454
rect 416146 309218 416382 309454
rect 415826 308898 416062 309134
rect 416146 308898 416382 309134
rect 415826 273218 416062 273454
rect 416146 273218 416382 273454
rect 415826 272898 416062 273134
rect 416146 272898 416382 273134
rect 415826 237218 416062 237454
rect 416146 237218 416382 237454
rect 415826 236898 416062 237134
rect 416146 236898 416382 237134
rect 415826 201218 416062 201454
rect 416146 201218 416382 201454
rect 415826 200898 416062 201134
rect 416146 200898 416382 201134
rect 415826 165218 416062 165454
rect 416146 165218 416382 165454
rect 415826 164898 416062 165134
rect 416146 164898 416382 165134
rect 415826 129218 416062 129454
rect 416146 129218 416382 129454
rect 415826 128898 416062 129134
rect 416146 128898 416382 129134
rect 415826 93218 416062 93454
rect 416146 93218 416382 93454
rect 415826 92898 416062 93134
rect 416146 92898 416382 93134
rect 415826 57218 416062 57454
rect 416146 57218 416382 57454
rect 415826 56898 416062 57134
rect 416146 56898 416382 57134
rect 415826 21218 416062 21454
rect 416146 21218 416382 21454
rect 415826 20898 416062 21134
rect 416146 20898 416382 21134
rect 415826 -1542 416062 -1306
rect 416146 -1542 416382 -1306
rect 415826 -1862 416062 -1626
rect 416146 -1862 416382 -1626
rect 419546 672938 419782 673174
rect 419866 672938 420102 673174
rect 419546 672618 419782 672854
rect 419866 672618 420102 672854
rect 419546 636938 419782 637174
rect 419866 636938 420102 637174
rect 419546 636618 419782 636854
rect 419866 636618 420102 636854
rect 419546 600938 419782 601174
rect 419866 600938 420102 601174
rect 419546 600618 419782 600854
rect 419866 600618 420102 600854
rect 419546 564938 419782 565174
rect 419866 564938 420102 565174
rect 419546 564618 419782 564854
rect 419866 564618 420102 564854
rect 419546 528938 419782 529174
rect 419866 528938 420102 529174
rect 419546 528618 419782 528854
rect 419866 528618 420102 528854
rect 419546 492938 419782 493174
rect 419866 492938 420102 493174
rect 419546 492618 419782 492854
rect 419866 492618 420102 492854
rect 419546 456938 419782 457174
rect 419866 456938 420102 457174
rect 419546 456618 419782 456854
rect 419866 456618 420102 456854
rect 419546 420938 419782 421174
rect 419866 420938 420102 421174
rect 419546 420618 419782 420854
rect 419866 420618 420102 420854
rect 419546 384938 419782 385174
rect 419866 384938 420102 385174
rect 419546 384618 419782 384854
rect 419866 384618 420102 384854
rect 419546 348938 419782 349174
rect 419866 348938 420102 349174
rect 419546 348618 419782 348854
rect 419866 348618 420102 348854
rect 419546 312938 419782 313174
rect 419866 312938 420102 313174
rect 419546 312618 419782 312854
rect 419866 312618 420102 312854
rect 419546 276938 419782 277174
rect 419866 276938 420102 277174
rect 419546 276618 419782 276854
rect 419866 276618 420102 276854
rect 419546 240938 419782 241174
rect 419866 240938 420102 241174
rect 419546 240618 419782 240854
rect 419866 240618 420102 240854
rect 419546 204938 419782 205174
rect 419866 204938 420102 205174
rect 419546 204618 419782 204854
rect 419866 204618 420102 204854
rect 419546 168938 419782 169174
rect 419866 168938 420102 169174
rect 419546 168618 419782 168854
rect 419866 168618 420102 168854
rect 419546 132938 419782 133174
rect 419866 132938 420102 133174
rect 419546 132618 419782 132854
rect 419866 132618 420102 132854
rect 419546 96938 419782 97174
rect 419866 96938 420102 97174
rect 419546 96618 419782 96854
rect 419866 96618 420102 96854
rect 419546 60938 419782 61174
rect 419866 60938 420102 61174
rect 419546 60618 419782 60854
rect 419866 60618 420102 60854
rect 419546 24938 419782 25174
rect 419866 24938 420102 25174
rect 419546 24618 419782 24854
rect 419866 24618 420102 24854
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 676658 423502 676894
rect 423586 676658 423822 676894
rect 423266 676338 423502 676574
rect 423586 676338 423822 676574
rect 423266 640658 423502 640894
rect 423586 640658 423822 640894
rect 423266 640338 423502 640574
rect 423586 640338 423822 640574
rect 423266 604658 423502 604894
rect 423586 604658 423822 604894
rect 423266 604338 423502 604574
rect 423586 604338 423822 604574
rect 423266 568658 423502 568894
rect 423586 568658 423822 568894
rect 423266 568338 423502 568574
rect 423586 568338 423822 568574
rect 423266 532658 423502 532894
rect 423586 532658 423822 532894
rect 423266 532338 423502 532574
rect 423586 532338 423822 532574
rect 423266 496658 423502 496894
rect 423586 496658 423822 496894
rect 423266 496338 423502 496574
rect 423586 496338 423822 496574
rect 423266 460658 423502 460894
rect 423586 460658 423822 460894
rect 423266 460338 423502 460574
rect 423586 460338 423822 460574
rect 423266 424658 423502 424894
rect 423586 424658 423822 424894
rect 423266 424338 423502 424574
rect 423586 424338 423822 424574
rect 423266 388658 423502 388894
rect 423586 388658 423822 388894
rect 423266 388338 423502 388574
rect 423586 388338 423822 388574
rect 423266 352658 423502 352894
rect 423586 352658 423822 352894
rect 423266 352338 423502 352574
rect 423586 352338 423822 352574
rect 423266 316658 423502 316894
rect 423586 316658 423822 316894
rect 423266 316338 423502 316574
rect 423586 316338 423822 316574
rect 423266 280658 423502 280894
rect 423586 280658 423822 280894
rect 423266 280338 423502 280574
rect 423586 280338 423822 280574
rect 423266 244658 423502 244894
rect 423586 244658 423822 244894
rect 423266 244338 423502 244574
rect 423586 244338 423822 244574
rect 423266 208658 423502 208894
rect 423586 208658 423822 208894
rect 423266 208338 423502 208574
rect 423586 208338 423822 208574
rect 423266 172658 423502 172894
rect 423586 172658 423822 172894
rect 423266 172338 423502 172574
rect 423586 172338 423822 172574
rect 423266 136658 423502 136894
rect 423586 136658 423822 136894
rect 423266 136338 423502 136574
rect 423586 136338 423822 136574
rect 423266 100658 423502 100894
rect 423586 100658 423822 100894
rect 423266 100338 423502 100574
rect 423586 100338 423822 100574
rect 423266 64658 423502 64894
rect 423586 64658 423822 64894
rect 423266 64338 423502 64574
rect 423586 64338 423822 64574
rect 423266 28658 423502 28894
rect 423586 28658 423822 28894
rect 423266 28338 423502 28574
rect 423586 28338 423822 28574
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 426986 680378 427222 680614
rect 427306 680378 427542 680614
rect 426986 680058 427222 680294
rect 427306 680058 427542 680294
rect 426986 644378 427222 644614
rect 427306 644378 427542 644614
rect 426986 644058 427222 644294
rect 427306 644058 427542 644294
rect 426986 608378 427222 608614
rect 427306 608378 427542 608614
rect 426986 608058 427222 608294
rect 427306 608058 427542 608294
rect 426986 572378 427222 572614
rect 427306 572378 427542 572614
rect 426986 572058 427222 572294
rect 427306 572058 427542 572294
rect 426986 536378 427222 536614
rect 427306 536378 427542 536614
rect 426986 536058 427222 536294
rect 427306 536058 427542 536294
rect 426986 500378 427222 500614
rect 427306 500378 427542 500614
rect 426986 500058 427222 500294
rect 427306 500058 427542 500294
rect 426986 464378 427222 464614
rect 427306 464378 427542 464614
rect 426986 464058 427222 464294
rect 427306 464058 427542 464294
rect 426986 428378 427222 428614
rect 427306 428378 427542 428614
rect 426986 428058 427222 428294
rect 427306 428058 427542 428294
rect 426986 392378 427222 392614
rect 427306 392378 427542 392614
rect 426986 392058 427222 392294
rect 427306 392058 427542 392294
rect 426986 356378 427222 356614
rect 427306 356378 427542 356614
rect 426986 356058 427222 356294
rect 427306 356058 427542 356294
rect 426986 320378 427222 320614
rect 427306 320378 427542 320614
rect 426986 320058 427222 320294
rect 427306 320058 427542 320294
rect 426986 284378 427222 284614
rect 427306 284378 427542 284614
rect 426986 284058 427222 284294
rect 427306 284058 427542 284294
rect 426986 248378 427222 248614
rect 427306 248378 427542 248614
rect 426986 248058 427222 248294
rect 427306 248058 427542 248294
rect 426986 212378 427222 212614
rect 427306 212378 427542 212614
rect 426986 212058 427222 212294
rect 427306 212058 427542 212294
rect 426986 176378 427222 176614
rect 427306 176378 427542 176614
rect 426986 176058 427222 176294
rect 427306 176058 427542 176294
rect 426986 140378 427222 140614
rect 427306 140378 427542 140614
rect 426986 140058 427222 140294
rect 427306 140058 427542 140294
rect 426986 104378 427222 104614
rect 427306 104378 427542 104614
rect 426986 104058 427222 104294
rect 427306 104058 427542 104294
rect 426986 68378 427222 68614
rect 427306 68378 427542 68614
rect 426986 68058 427222 68294
rect 427306 68058 427542 68294
rect 426986 32378 427222 32614
rect 427306 32378 427542 32614
rect 426986 32058 427222 32294
rect 427306 32058 427542 32294
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 433826 687218 434062 687454
rect 434146 687218 434382 687454
rect 433826 686898 434062 687134
rect 434146 686898 434382 687134
rect 433826 651218 434062 651454
rect 434146 651218 434382 651454
rect 433826 650898 434062 651134
rect 434146 650898 434382 651134
rect 433826 615218 434062 615454
rect 434146 615218 434382 615454
rect 433826 614898 434062 615134
rect 434146 614898 434382 615134
rect 433826 579218 434062 579454
rect 434146 579218 434382 579454
rect 433826 578898 434062 579134
rect 434146 578898 434382 579134
rect 433826 543218 434062 543454
rect 434146 543218 434382 543454
rect 433826 542898 434062 543134
rect 434146 542898 434382 543134
rect 433826 507218 434062 507454
rect 434146 507218 434382 507454
rect 433826 506898 434062 507134
rect 434146 506898 434382 507134
rect 433826 471218 434062 471454
rect 434146 471218 434382 471454
rect 433826 470898 434062 471134
rect 434146 470898 434382 471134
rect 433826 435218 434062 435454
rect 434146 435218 434382 435454
rect 433826 434898 434062 435134
rect 434146 434898 434382 435134
rect 433826 399218 434062 399454
rect 434146 399218 434382 399454
rect 433826 398898 434062 399134
rect 434146 398898 434382 399134
rect 433826 363218 434062 363454
rect 434146 363218 434382 363454
rect 433826 362898 434062 363134
rect 434146 362898 434382 363134
rect 433826 327218 434062 327454
rect 434146 327218 434382 327454
rect 433826 326898 434062 327134
rect 434146 326898 434382 327134
rect 433826 291218 434062 291454
rect 434146 291218 434382 291454
rect 433826 290898 434062 291134
rect 434146 290898 434382 291134
rect 433826 255218 434062 255454
rect 434146 255218 434382 255454
rect 433826 254898 434062 255134
rect 434146 254898 434382 255134
rect 433826 219218 434062 219454
rect 434146 219218 434382 219454
rect 433826 218898 434062 219134
rect 434146 218898 434382 219134
rect 433826 183218 434062 183454
rect 434146 183218 434382 183454
rect 433826 182898 434062 183134
rect 434146 182898 434382 183134
rect 433826 147218 434062 147454
rect 434146 147218 434382 147454
rect 433826 146898 434062 147134
rect 434146 146898 434382 147134
rect 433826 111218 434062 111454
rect 434146 111218 434382 111454
rect 433826 110898 434062 111134
rect 434146 110898 434382 111134
rect 433826 75218 434062 75454
rect 434146 75218 434382 75454
rect 433826 74898 434062 75134
rect 434146 74898 434382 75134
rect 433826 39218 434062 39454
rect 434146 39218 434382 39454
rect 433826 38898 434062 39134
rect 434146 38898 434382 39134
rect 433826 3218 434062 3454
rect 434146 3218 434382 3454
rect 433826 2898 434062 3134
rect 434146 2898 434382 3134
rect 433826 -582 434062 -346
rect 434146 -582 434382 -346
rect 433826 -902 434062 -666
rect 434146 -902 434382 -666
rect 437546 690938 437782 691174
rect 437866 690938 438102 691174
rect 437546 690618 437782 690854
rect 437866 690618 438102 690854
rect 437546 654938 437782 655174
rect 437866 654938 438102 655174
rect 437546 654618 437782 654854
rect 437866 654618 438102 654854
rect 437546 618938 437782 619174
rect 437866 618938 438102 619174
rect 437546 618618 437782 618854
rect 437866 618618 438102 618854
rect 437546 582938 437782 583174
rect 437866 582938 438102 583174
rect 437546 582618 437782 582854
rect 437866 582618 438102 582854
rect 437546 546938 437782 547174
rect 437866 546938 438102 547174
rect 437546 546618 437782 546854
rect 437866 546618 438102 546854
rect 437546 510938 437782 511174
rect 437866 510938 438102 511174
rect 437546 510618 437782 510854
rect 437866 510618 438102 510854
rect 437546 474938 437782 475174
rect 437866 474938 438102 475174
rect 437546 474618 437782 474854
rect 437866 474618 438102 474854
rect 437546 438938 437782 439174
rect 437866 438938 438102 439174
rect 437546 438618 437782 438854
rect 437866 438618 438102 438854
rect 437546 402938 437782 403174
rect 437866 402938 438102 403174
rect 437546 402618 437782 402854
rect 437866 402618 438102 402854
rect 437546 366938 437782 367174
rect 437866 366938 438102 367174
rect 437546 366618 437782 366854
rect 437866 366618 438102 366854
rect 437546 330938 437782 331174
rect 437866 330938 438102 331174
rect 437546 330618 437782 330854
rect 437866 330618 438102 330854
rect 437546 294938 437782 295174
rect 437866 294938 438102 295174
rect 437546 294618 437782 294854
rect 437866 294618 438102 294854
rect 437546 258938 437782 259174
rect 437866 258938 438102 259174
rect 437546 258618 437782 258854
rect 437866 258618 438102 258854
rect 437546 222938 437782 223174
rect 437866 222938 438102 223174
rect 437546 222618 437782 222854
rect 437866 222618 438102 222854
rect 437546 186938 437782 187174
rect 437866 186938 438102 187174
rect 437546 186618 437782 186854
rect 437866 186618 438102 186854
rect 437546 150938 437782 151174
rect 437866 150938 438102 151174
rect 437546 150618 437782 150854
rect 437866 150618 438102 150854
rect 437546 114938 437782 115174
rect 437866 114938 438102 115174
rect 437546 114618 437782 114854
rect 437866 114618 438102 114854
rect 437546 78938 437782 79174
rect 437866 78938 438102 79174
rect 437546 78618 437782 78854
rect 437866 78618 438102 78854
rect 437546 42938 437782 43174
rect 437866 42938 438102 43174
rect 437546 42618 437782 42854
rect 437866 42618 438102 42854
rect 437546 6938 437782 7174
rect 437866 6938 438102 7174
rect 437546 6618 437782 6854
rect 437866 6618 438102 6854
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 694658 441502 694894
rect 441586 694658 441822 694894
rect 441266 694338 441502 694574
rect 441586 694338 441822 694574
rect 441266 658658 441502 658894
rect 441586 658658 441822 658894
rect 441266 658338 441502 658574
rect 441586 658338 441822 658574
rect 441266 622658 441502 622894
rect 441586 622658 441822 622894
rect 441266 622338 441502 622574
rect 441586 622338 441822 622574
rect 441266 586658 441502 586894
rect 441586 586658 441822 586894
rect 441266 586338 441502 586574
rect 441586 586338 441822 586574
rect 441266 550658 441502 550894
rect 441586 550658 441822 550894
rect 441266 550338 441502 550574
rect 441586 550338 441822 550574
rect 441266 514658 441502 514894
rect 441586 514658 441822 514894
rect 441266 514338 441502 514574
rect 441586 514338 441822 514574
rect 441266 478658 441502 478894
rect 441586 478658 441822 478894
rect 441266 478338 441502 478574
rect 441586 478338 441822 478574
rect 441266 442658 441502 442894
rect 441586 442658 441822 442894
rect 441266 442338 441502 442574
rect 441586 442338 441822 442574
rect 441266 406658 441502 406894
rect 441586 406658 441822 406894
rect 441266 406338 441502 406574
rect 441586 406338 441822 406574
rect 441266 370658 441502 370894
rect 441586 370658 441822 370894
rect 441266 370338 441502 370574
rect 441586 370338 441822 370574
rect 441266 334658 441502 334894
rect 441586 334658 441822 334894
rect 441266 334338 441502 334574
rect 441586 334338 441822 334574
rect 441266 298658 441502 298894
rect 441586 298658 441822 298894
rect 441266 298338 441502 298574
rect 441586 298338 441822 298574
rect 441266 262658 441502 262894
rect 441586 262658 441822 262894
rect 441266 262338 441502 262574
rect 441586 262338 441822 262574
rect 441266 226658 441502 226894
rect 441586 226658 441822 226894
rect 441266 226338 441502 226574
rect 441586 226338 441822 226574
rect 441266 190658 441502 190894
rect 441586 190658 441822 190894
rect 441266 190338 441502 190574
rect 441586 190338 441822 190574
rect 441266 154658 441502 154894
rect 441586 154658 441822 154894
rect 441266 154338 441502 154574
rect 441586 154338 441822 154574
rect 441266 118658 441502 118894
rect 441586 118658 441822 118894
rect 441266 118338 441502 118574
rect 441586 118338 441822 118574
rect 441266 82658 441502 82894
rect 441586 82658 441822 82894
rect 441266 82338 441502 82574
rect 441586 82338 441822 82574
rect 441266 46658 441502 46894
rect 441586 46658 441822 46894
rect 441266 46338 441502 46574
rect 441586 46338 441822 46574
rect 441266 10658 441502 10894
rect 441586 10658 441822 10894
rect 441266 10338 441502 10574
rect 441586 10338 441822 10574
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 444986 698378 445222 698614
rect 445306 698378 445542 698614
rect 444986 698058 445222 698294
rect 445306 698058 445542 698294
rect 444986 662378 445222 662614
rect 445306 662378 445542 662614
rect 444986 662058 445222 662294
rect 445306 662058 445542 662294
rect 444986 626378 445222 626614
rect 445306 626378 445542 626614
rect 444986 626058 445222 626294
rect 445306 626058 445542 626294
rect 444986 590378 445222 590614
rect 445306 590378 445542 590614
rect 444986 590058 445222 590294
rect 445306 590058 445542 590294
rect 444986 554378 445222 554614
rect 445306 554378 445542 554614
rect 444986 554058 445222 554294
rect 445306 554058 445542 554294
rect 444986 518378 445222 518614
rect 445306 518378 445542 518614
rect 444986 518058 445222 518294
rect 445306 518058 445542 518294
rect 444986 482378 445222 482614
rect 445306 482378 445542 482614
rect 444986 482058 445222 482294
rect 445306 482058 445542 482294
rect 444986 446378 445222 446614
rect 445306 446378 445542 446614
rect 444986 446058 445222 446294
rect 445306 446058 445542 446294
rect 444986 410378 445222 410614
rect 445306 410378 445542 410614
rect 444986 410058 445222 410294
rect 445306 410058 445542 410294
rect 444986 374378 445222 374614
rect 445306 374378 445542 374614
rect 444986 374058 445222 374294
rect 445306 374058 445542 374294
rect 444986 338378 445222 338614
rect 445306 338378 445542 338614
rect 444986 338058 445222 338294
rect 445306 338058 445542 338294
rect 444986 302378 445222 302614
rect 445306 302378 445542 302614
rect 444986 302058 445222 302294
rect 445306 302058 445542 302294
rect 444986 266378 445222 266614
rect 445306 266378 445542 266614
rect 444986 266058 445222 266294
rect 445306 266058 445542 266294
rect 444986 230378 445222 230614
rect 445306 230378 445542 230614
rect 444986 230058 445222 230294
rect 445306 230058 445542 230294
rect 444986 194378 445222 194614
rect 445306 194378 445542 194614
rect 444986 194058 445222 194294
rect 445306 194058 445542 194294
rect 444986 158378 445222 158614
rect 445306 158378 445542 158614
rect 444986 158058 445222 158294
rect 445306 158058 445542 158294
rect 444986 122378 445222 122614
rect 445306 122378 445542 122614
rect 444986 122058 445222 122294
rect 445306 122058 445542 122294
rect 444986 86378 445222 86614
rect 445306 86378 445542 86614
rect 444986 86058 445222 86294
rect 445306 86058 445542 86294
rect 444986 50378 445222 50614
rect 445306 50378 445542 50614
rect 444986 50058 445222 50294
rect 445306 50058 445542 50294
rect 444986 14378 445222 14614
rect 445306 14378 445542 14614
rect 444986 14058 445222 14294
rect 445306 14058 445542 14294
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 451826 669218 452062 669454
rect 452146 669218 452382 669454
rect 451826 668898 452062 669134
rect 452146 668898 452382 669134
rect 451826 633218 452062 633454
rect 452146 633218 452382 633454
rect 451826 632898 452062 633134
rect 452146 632898 452382 633134
rect 451826 597218 452062 597454
rect 452146 597218 452382 597454
rect 451826 596898 452062 597134
rect 452146 596898 452382 597134
rect 451826 561218 452062 561454
rect 452146 561218 452382 561454
rect 451826 560898 452062 561134
rect 452146 560898 452382 561134
rect 451826 525218 452062 525454
rect 452146 525218 452382 525454
rect 451826 524898 452062 525134
rect 452146 524898 452382 525134
rect 451826 489218 452062 489454
rect 452146 489218 452382 489454
rect 451826 488898 452062 489134
rect 452146 488898 452382 489134
rect 451826 453218 452062 453454
rect 452146 453218 452382 453454
rect 451826 452898 452062 453134
rect 452146 452898 452382 453134
rect 451826 417218 452062 417454
rect 452146 417218 452382 417454
rect 451826 416898 452062 417134
rect 452146 416898 452382 417134
rect 451826 381218 452062 381454
rect 452146 381218 452382 381454
rect 451826 380898 452062 381134
rect 452146 380898 452382 381134
rect 451826 345218 452062 345454
rect 452146 345218 452382 345454
rect 451826 344898 452062 345134
rect 452146 344898 452382 345134
rect 451826 309218 452062 309454
rect 452146 309218 452382 309454
rect 451826 308898 452062 309134
rect 452146 308898 452382 309134
rect 451826 273218 452062 273454
rect 452146 273218 452382 273454
rect 451826 272898 452062 273134
rect 452146 272898 452382 273134
rect 451826 237218 452062 237454
rect 452146 237218 452382 237454
rect 451826 236898 452062 237134
rect 452146 236898 452382 237134
rect 451826 201218 452062 201454
rect 452146 201218 452382 201454
rect 451826 200898 452062 201134
rect 452146 200898 452382 201134
rect 451826 165218 452062 165454
rect 452146 165218 452382 165454
rect 451826 164898 452062 165134
rect 452146 164898 452382 165134
rect 451826 129218 452062 129454
rect 452146 129218 452382 129454
rect 451826 128898 452062 129134
rect 452146 128898 452382 129134
rect 451826 93218 452062 93454
rect 452146 93218 452382 93454
rect 451826 92898 452062 93134
rect 452146 92898 452382 93134
rect 451826 57218 452062 57454
rect 452146 57218 452382 57454
rect 451826 56898 452062 57134
rect 452146 56898 452382 57134
rect 451826 21218 452062 21454
rect 452146 21218 452382 21454
rect 451826 20898 452062 21134
rect 452146 20898 452382 21134
rect 451826 -1542 452062 -1306
rect 452146 -1542 452382 -1306
rect 451826 -1862 452062 -1626
rect 452146 -1862 452382 -1626
rect 455546 672938 455782 673174
rect 455866 672938 456102 673174
rect 455546 672618 455782 672854
rect 455866 672618 456102 672854
rect 455546 636938 455782 637174
rect 455866 636938 456102 637174
rect 455546 636618 455782 636854
rect 455866 636618 456102 636854
rect 455546 600938 455782 601174
rect 455866 600938 456102 601174
rect 455546 600618 455782 600854
rect 455866 600618 456102 600854
rect 455546 564938 455782 565174
rect 455866 564938 456102 565174
rect 455546 564618 455782 564854
rect 455866 564618 456102 564854
rect 455546 528938 455782 529174
rect 455866 528938 456102 529174
rect 455546 528618 455782 528854
rect 455866 528618 456102 528854
rect 455546 492938 455782 493174
rect 455866 492938 456102 493174
rect 455546 492618 455782 492854
rect 455866 492618 456102 492854
rect 455546 456938 455782 457174
rect 455866 456938 456102 457174
rect 455546 456618 455782 456854
rect 455866 456618 456102 456854
rect 455546 420938 455782 421174
rect 455866 420938 456102 421174
rect 455546 420618 455782 420854
rect 455866 420618 456102 420854
rect 455546 384938 455782 385174
rect 455866 384938 456102 385174
rect 455546 384618 455782 384854
rect 455866 384618 456102 384854
rect 455546 348938 455782 349174
rect 455866 348938 456102 349174
rect 455546 348618 455782 348854
rect 455866 348618 456102 348854
rect 455546 312938 455782 313174
rect 455866 312938 456102 313174
rect 455546 312618 455782 312854
rect 455866 312618 456102 312854
rect 455546 276938 455782 277174
rect 455866 276938 456102 277174
rect 455546 276618 455782 276854
rect 455866 276618 456102 276854
rect 455546 240938 455782 241174
rect 455866 240938 456102 241174
rect 455546 240618 455782 240854
rect 455866 240618 456102 240854
rect 455546 204938 455782 205174
rect 455866 204938 456102 205174
rect 455546 204618 455782 204854
rect 455866 204618 456102 204854
rect 455546 168938 455782 169174
rect 455866 168938 456102 169174
rect 455546 168618 455782 168854
rect 455866 168618 456102 168854
rect 455546 132938 455782 133174
rect 455866 132938 456102 133174
rect 455546 132618 455782 132854
rect 455866 132618 456102 132854
rect 455546 96938 455782 97174
rect 455866 96938 456102 97174
rect 455546 96618 455782 96854
rect 455866 96618 456102 96854
rect 455546 60938 455782 61174
rect 455866 60938 456102 61174
rect 455546 60618 455782 60854
rect 455866 60618 456102 60854
rect 455546 24938 455782 25174
rect 455866 24938 456102 25174
rect 455546 24618 455782 24854
rect 455866 24618 456102 24854
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 676658 459502 676894
rect 459586 676658 459822 676894
rect 459266 676338 459502 676574
rect 459586 676338 459822 676574
rect 459266 640658 459502 640894
rect 459586 640658 459822 640894
rect 459266 640338 459502 640574
rect 459586 640338 459822 640574
rect 459266 604658 459502 604894
rect 459586 604658 459822 604894
rect 459266 604338 459502 604574
rect 459586 604338 459822 604574
rect 459266 568658 459502 568894
rect 459586 568658 459822 568894
rect 459266 568338 459502 568574
rect 459586 568338 459822 568574
rect 459266 532658 459502 532894
rect 459586 532658 459822 532894
rect 459266 532338 459502 532574
rect 459586 532338 459822 532574
rect 459266 496658 459502 496894
rect 459586 496658 459822 496894
rect 459266 496338 459502 496574
rect 459586 496338 459822 496574
rect 459266 460658 459502 460894
rect 459586 460658 459822 460894
rect 459266 460338 459502 460574
rect 459586 460338 459822 460574
rect 459266 424658 459502 424894
rect 459586 424658 459822 424894
rect 459266 424338 459502 424574
rect 459586 424338 459822 424574
rect 459266 388658 459502 388894
rect 459586 388658 459822 388894
rect 459266 388338 459502 388574
rect 459586 388338 459822 388574
rect 459266 352658 459502 352894
rect 459586 352658 459822 352894
rect 459266 352338 459502 352574
rect 459586 352338 459822 352574
rect 459266 316658 459502 316894
rect 459586 316658 459822 316894
rect 459266 316338 459502 316574
rect 459586 316338 459822 316574
rect 459266 280658 459502 280894
rect 459586 280658 459822 280894
rect 459266 280338 459502 280574
rect 459586 280338 459822 280574
rect 459266 244658 459502 244894
rect 459586 244658 459822 244894
rect 459266 244338 459502 244574
rect 459586 244338 459822 244574
rect 459266 208658 459502 208894
rect 459586 208658 459822 208894
rect 459266 208338 459502 208574
rect 459586 208338 459822 208574
rect 459266 172658 459502 172894
rect 459586 172658 459822 172894
rect 459266 172338 459502 172574
rect 459586 172338 459822 172574
rect 459266 136658 459502 136894
rect 459586 136658 459822 136894
rect 459266 136338 459502 136574
rect 459586 136338 459822 136574
rect 459266 100658 459502 100894
rect 459586 100658 459822 100894
rect 459266 100338 459502 100574
rect 459586 100338 459822 100574
rect 459266 64658 459502 64894
rect 459586 64658 459822 64894
rect 459266 64338 459502 64574
rect 459586 64338 459822 64574
rect 459266 28658 459502 28894
rect 459586 28658 459822 28894
rect 459266 28338 459502 28574
rect 459586 28338 459822 28574
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 462986 680378 463222 680614
rect 463306 680378 463542 680614
rect 462986 680058 463222 680294
rect 463306 680058 463542 680294
rect 462986 644378 463222 644614
rect 463306 644378 463542 644614
rect 462986 644058 463222 644294
rect 463306 644058 463542 644294
rect 462986 608378 463222 608614
rect 463306 608378 463542 608614
rect 462986 608058 463222 608294
rect 463306 608058 463542 608294
rect 462986 572378 463222 572614
rect 463306 572378 463542 572614
rect 462986 572058 463222 572294
rect 463306 572058 463542 572294
rect 462986 536378 463222 536614
rect 463306 536378 463542 536614
rect 462986 536058 463222 536294
rect 463306 536058 463542 536294
rect 462986 500378 463222 500614
rect 463306 500378 463542 500614
rect 462986 500058 463222 500294
rect 463306 500058 463542 500294
rect 462986 464378 463222 464614
rect 463306 464378 463542 464614
rect 462986 464058 463222 464294
rect 463306 464058 463542 464294
rect 462986 428378 463222 428614
rect 463306 428378 463542 428614
rect 462986 428058 463222 428294
rect 463306 428058 463542 428294
rect 462986 392378 463222 392614
rect 463306 392378 463542 392614
rect 462986 392058 463222 392294
rect 463306 392058 463542 392294
rect 462986 356378 463222 356614
rect 463306 356378 463542 356614
rect 462986 356058 463222 356294
rect 463306 356058 463542 356294
rect 462986 320378 463222 320614
rect 463306 320378 463542 320614
rect 462986 320058 463222 320294
rect 463306 320058 463542 320294
rect 462986 284378 463222 284614
rect 463306 284378 463542 284614
rect 462986 284058 463222 284294
rect 463306 284058 463542 284294
rect 462986 248378 463222 248614
rect 463306 248378 463542 248614
rect 462986 248058 463222 248294
rect 463306 248058 463542 248294
rect 462986 212378 463222 212614
rect 463306 212378 463542 212614
rect 462986 212058 463222 212294
rect 463306 212058 463542 212294
rect 462986 176378 463222 176614
rect 463306 176378 463542 176614
rect 462986 176058 463222 176294
rect 463306 176058 463542 176294
rect 462986 140378 463222 140614
rect 463306 140378 463542 140614
rect 462986 140058 463222 140294
rect 463306 140058 463542 140294
rect 462986 104378 463222 104614
rect 463306 104378 463542 104614
rect 462986 104058 463222 104294
rect 463306 104058 463542 104294
rect 462986 68378 463222 68614
rect 463306 68378 463542 68614
rect 462986 68058 463222 68294
rect 463306 68058 463542 68294
rect 462986 32378 463222 32614
rect 463306 32378 463542 32614
rect 462986 32058 463222 32294
rect 463306 32058 463542 32294
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 469826 687218 470062 687454
rect 470146 687218 470382 687454
rect 469826 686898 470062 687134
rect 470146 686898 470382 687134
rect 469826 651218 470062 651454
rect 470146 651218 470382 651454
rect 469826 650898 470062 651134
rect 470146 650898 470382 651134
rect 469826 615218 470062 615454
rect 470146 615218 470382 615454
rect 469826 614898 470062 615134
rect 470146 614898 470382 615134
rect 469826 579218 470062 579454
rect 470146 579218 470382 579454
rect 469826 578898 470062 579134
rect 470146 578898 470382 579134
rect 469826 543218 470062 543454
rect 470146 543218 470382 543454
rect 469826 542898 470062 543134
rect 470146 542898 470382 543134
rect 469826 507218 470062 507454
rect 470146 507218 470382 507454
rect 469826 506898 470062 507134
rect 470146 506898 470382 507134
rect 469826 471218 470062 471454
rect 470146 471218 470382 471454
rect 469826 470898 470062 471134
rect 470146 470898 470382 471134
rect 469826 435218 470062 435454
rect 470146 435218 470382 435454
rect 469826 434898 470062 435134
rect 470146 434898 470382 435134
rect 469826 399218 470062 399454
rect 470146 399218 470382 399454
rect 469826 398898 470062 399134
rect 470146 398898 470382 399134
rect 469826 363218 470062 363454
rect 470146 363218 470382 363454
rect 469826 362898 470062 363134
rect 470146 362898 470382 363134
rect 469826 327218 470062 327454
rect 470146 327218 470382 327454
rect 469826 326898 470062 327134
rect 470146 326898 470382 327134
rect 469826 291218 470062 291454
rect 470146 291218 470382 291454
rect 469826 290898 470062 291134
rect 470146 290898 470382 291134
rect 469826 255218 470062 255454
rect 470146 255218 470382 255454
rect 469826 254898 470062 255134
rect 470146 254898 470382 255134
rect 469826 219218 470062 219454
rect 470146 219218 470382 219454
rect 469826 218898 470062 219134
rect 470146 218898 470382 219134
rect 469826 183218 470062 183454
rect 470146 183218 470382 183454
rect 469826 182898 470062 183134
rect 470146 182898 470382 183134
rect 469826 147218 470062 147454
rect 470146 147218 470382 147454
rect 469826 146898 470062 147134
rect 470146 146898 470382 147134
rect 469826 111218 470062 111454
rect 470146 111218 470382 111454
rect 469826 110898 470062 111134
rect 470146 110898 470382 111134
rect 469826 75218 470062 75454
rect 470146 75218 470382 75454
rect 469826 74898 470062 75134
rect 470146 74898 470382 75134
rect 469826 39218 470062 39454
rect 470146 39218 470382 39454
rect 469826 38898 470062 39134
rect 470146 38898 470382 39134
rect 469826 3218 470062 3454
rect 470146 3218 470382 3454
rect 469826 2898 470062 3134
rect 470146 2898 470382 3134
rect 469826 -582 470062 -346
rect 470146 -582 470382 -346
rect 469826 -902 470062 -666
rect 470146 -902 470382 -666
rect 473546 690938 473782 691174
rect 473866 690938 474102 691174
rect 473546 690618 473782 690854
rect 473866 690618 474102 690854
rect 473546 654938 473782 655174
rect 473866 654938 474102 655174
rect 473546 654618 473782 654854
rect 473866 654618 474102 654854
rect 473546 618938 473782 619174
rect 473866 618938 474102 619174
rect 473546 618618 473782 618854
rect 473866 618618 474102 618854
rect 473546 582938 473782 583174
rect 473866 582938 474102 583174
rect 473546 582618 473782 582854
rect 473866 582618 474102 582854
rect 473546 546938 473782 547174
rect 473866 546938 474102 547174
rect 473546 546618 473782 546854
rect 473866 546618 474102 546854
rect 473546 510938 473782 511174
rect 473866 510938 474102 511174
rect 473546 510618 473782 510854
rect 473866 510618 474102 510854
rect 473546 474938 473782 475174
rect 473866 474938 474102 475174
rect 473546 474618 473782 474854
rect 473866 474618 474102 474854
rect 473546 438938 473782 439174
rect 473866 438938 474102 439174
rect 473546 438618 473782 438854
rect 473866 438618 474102 438854
rect 473546 402938 473782 403174
rect 473866 402938 474102 403174
rect 473546 402618 473782 402854
rect 473866 402618 474102 402854
rect 473546 366938 473782 367174
rect 473866 366938 474102 367174
rect 473546 366618 473782 366854
rect 473866 366618 474102 366854
rect 473546 330938 473782 331174
rect 473866 330938 474102 331174
rect 473546 330618 473782 330854
rect 473866 330618 474102 330854
rect 473546 294938 473782 295174
rect 473866 294938 474102 295174
rect 473546 294618 473782 294854
rect 473866 294618 474102 294854
rect 473546 258938 473782 259174
rect 473866 258938 474102 259174
rect 473546 258618 473782 258854
rect 473866 258618 474102 258854
rect 473546 222938 473782 223174
rect 473866 222938 474102 223174
rect 473546 222618 473782 222854
rect 473866 222618 474102 222854
rect 473546 186938 473782 187174
rect 473866 186938 474102 187174
rect 473546 186618 473782 186854
rect 473866 186618 474102 186854
rect 473546 150938 473782 151174
rect 473866 150938 474102 151174
rect 473546 150618 473782 150854
rect 473866 150618 474102 150854
rect 473546 114938 473782 115174
rect 473866 114938 474102 115174
rect 473546 114618 473782 114854
rect 473866 114618 474102 114854
rect 473546 78938 473782 79174
rect 473866 78938 474102 79174
rect 473546 78618 473782 78854
rect 473866 78618 474102 78854
rect 473546 42938 473782 43174
rect 473866 42938 474102 43174
rect 473546 42618 473782 42854
rect 473866 42618 474102 42854
rect 473546 6938 473782 7174
rect 473866 6938 474102 7174
rect 473546 6618 473782 6854
rect 473866 6618 474102 6854
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 694658 477502 694894
rect 477586 694658 477822 694894
rect 477266 694338 477502 694574
rect 477586 694338 477822 694574
rect 477266 658658 477502 658894
rect 477586 658658 477822 658894
rect 477266 658338 477502 658574
rect 477586 658338 477822 658574
rect 477266 622658 477502 622894
rect 477586 622658 477822 622894
rect 477266 622338 477502 622574
rect 477586 622338 477822 622574
rect 477266 586658 477502 586894
rect 477586 586658 477822 586894
rect 477266 586338 477502 586574
rect 477586 586338 477822 586574
rect 477266 550658 477502 550894
rect 477586 550658 477822 550894
rect 477266 550338 477502 550574
rect 477586 550338 477822 550574
rect 477266 514658 477502 514894
rect 477586 514658 477822 514894
rect 477266 514338 477502 514574
rect 477586 514338 477822 514574
rect 477266 478658 477502 478894
rect 477586 478658 477822 478894
rect 477266 478338 477502 478574
rect 477586 478338 477822 478574
rect 477266 442658 477502 442894
rect 477586 442658 477822 442894
rect 477266 442338 477502 442574
rect 477586 442338 477822 442574
rect 477266 406658 477502 406894
rect 477586 406658 477822 406894
rect 477266 406338 477502 406574
rect 477586 406338 477822 406574
rect 477266 370658 477502 370894
rect 477586 370658 477822 370894
rect 477266 370338 477502 370574
rect 477586 370338 477822 370574
rect 477266 334658 477502 334894
rect 477586 334658 477822 334894
rect 477266 334338 477502 334574
rect 477586 334338 477822 334574
rect 477266 298658 477502 298894
rect 477586 298658 477822 298894
rect 477266 298338 477502 298574
rect 477586 298338 477822 298574
rect 477266 262658 477502 262894
rect 477586 262658 477822 262894
rect 477266 262338 477502 262574
rect 477586 262338 477822 262574
rect 477266 226658 477502 226894
rect 477586 226658 477822 226894
rect 477266 226338 477502 226574
rect 477586 226338 477822 226574
rect 477266 190658 477502 190894
rect 477586 190658 477822 190894
rect 477266 190338 477502 190574
rect 477586 190338 477822 190574
rect 477266 154658 477502 154894
rect 477586 154658 477822 154894
rect 477266 154338 477502 154574
rect 477586 154338 477822 154574
rect 477266 118658 477502 118894
rect 477586 118658 477822 118894
rect 477266 118338 477502 118574
rect 477586 118338 477822 118574
rect 477266 82658 477502 82894
rect 477586 82658 477822 82894
rect 477266 82338 477502 82574
rect 477586 82338 477822 82574
rect 477266 46658 477502 46894
rect 477586 46658 477822 46894
rect 477266 46338 477502 46574
rect 477586 46338 477822 46574
rect 477266 10658 477502 10894
rect 477586 10658 477822 10894
rect 477266 10338 477502 10574
rect 477586 10338 477822 10574
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 480986 698378 481222 698614
rect 481306 698378 481542 698614
rect 480986 698058 481222 698294
rect 481306 698058 481542 698294
rect 480986 662378 481222 662614
rect 481306 662378 481542 662614
rect 480986 662058 481222 662294
rect 481306 662058 481542 662294
rect 480986 626378 481222 626614
rect 481306 626378 481542 626614
rect 480986 626058 481222 626294
rect 481306 626058 481542 626294
rect 480986 590378 481222 590614
rect 481306 590378 481542 590614
rect 480986 590058 481222 590294
rect 481306 590058 481542 590294
rect 480986 554378 481222 554614
rect 481306 554378 481542 554614
rect 480986 554058 481222 554294
rect 481306 554058 481542 554294
rect 480986 518378 481222 518614
rect 481306 518378 481542 518614
rect 480986 518058 481222 518294
rect 481306 518058 481542 518294
rect 480986 482378 481222 482614
rect 481306 482378 481542 482614
rect 480986 482058 481222 482294
rect 481306 482058 481542 482294
rect 480986 446378 481222 446614
rect 481306 446378 481542 446614
rect 480986 446058 481222 446294
rect 481306 446058 481542 446294
rect 480986 410378 481222 410614
rect 481306 410378 481542 410614
rect 480986 410058 481222 410294
rect 481306 410058 481542 410294
rect 480986 374378 481222 374614
rect 481306 374378 481542 374614
rect 480986 374058 481222 374294
rect 481306 374058 481542 374294
rect 480986 338378 481222 338614
rect 481306 338378 481542 338614
rect 480986 338058 481222 338294
rect 481306 338058 481542 338294
rect 480986 302378 481222 302614
rect 481306 302378 481542 302614
rect 480986 302058 481222 302294
rect 481306 302058 481542 302294
rect 480986 266378 481222 266614
rect 481306 266378 481542 266614
rect 480986 266058 481222 266294
rect 481306 266058 481542 266294
rect 480986 230378 481222 230614
rect 481306 230378 481542 230614
rect 480986 230058 481222 230294
rect 481306 230058 481542 230294
rect 480986 194378 481222 194614
rect 481306 194378 481542 194614
rect 480986 194058 481222 194294
rect 481306 194058 481542 194294
rect 480986 158378 481222 158614
rect 481306 158378 481542 158614
rect 480986 158058 481222 158294
rect 481306 158058 481542 158294
rect 480986 122378 481222 122614
rect 481306 122378 481542 122614
rect 480986 122058 481222 122294
rect 481306 122058 481542 122294
rect 480986 86378 481222 86614
rect 481306 86378 481542 86614
rect 480986 86058 481222 86294
rect 481306 86058 481542 86294
rect 480986 50378 481222 50614
rect 481306 50378 481542 50614
rect 480986 50058 481222 50294
rect 481306 50058 481542 50294
rect 480986 14378 481222 14614
rect 481306 14378 481542 14614
rect 480986 14058 481222 14294
rect 481306 14058 481542 14294
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 487826 669218 488062 669454
rect 488146 669218 488382 669454
rect 487826 668898 488062 669134
rect 488146 668898 488382 669134
rect 487826 633218 488062 633454
rect 488146 633218 488382 633454
rect 487826 632898 488062 633134
rect 488146 632898 488382 633134
rect 487826 597218 488062 597454
rect 488146 597218 488382 597454
rect 487826 596898 488062 597134
rect 488146 596898 488382 597134
rect 487826 561218 488062 561454
rect 488146 561218 488382 561454
rect 487826 560898 488062 561134
rect 488146 560898 488382 561134
rect 487826 525218 488062 525454
rect 488146 525218 488382 525454
rect 487826 524898 488062 525134
rect 488146 524898 488382 525134
rect 487826 489218 488062 489454
rect 488146 489218 488382 489454
rect 487826 488898 488062 489134
rect 488146 488898 488382 489134
rect 487826 453218 488062 453454
rect 488146 453218 488382 453454
rect 487826 452898 488062 453134
rect 488146 452898 488382 453134
rect 487826 417218 488062 417454
rect 488146 417218 488382 417454
rect 487826 416898 488062 417134
rect 488146 416898 488382 417134
rect 487826 381218 488062 381454
rect 488146 381218 488382 381454
rect 487826 380898 488062 381134
rect 488146 380898 488382 381134
rect 487826 345218 488062 345454
rect 488146 345218 488382 345454
rect 487826 344898 488062 345134
rect 488146 344898 488382 345134
rect 487826 309218 488062 309454
rect 488146 309218 488382 309454
rect 487826 308898 488062 309134
rect 488146 308898 488382 309134
rect 487826 273218 488062 273454
rect 488146 273218 488382 273454
rect 487826 272898 488062 273134
rect 488146 272898 488382 273134
rect 487826 237218 488062 237454
rect 488146 237218 488382 237454
rect 487826 236898 488062 237134
rect 488146 236898 488382 237134
rect 487826 201218 488062 201454
rect 488146 201218 488382 201454
rect 487826 200898 488062 201134
rect 488146 200898 488382 201134
rect 487826 165218 488062 165454
rect 488146 165218 488382 165454
rect 487826 164898 488062 165134
rect 488146 164898 488382 165134
rect 487826 129218 488062 129454
rect 488146 129218 488382 129454
rect 487826 128898 488062 129134
rect 488146 128898 488382 129134
rect 487826 93218 488062 93454
rect 488146 93218 488382 93454
rect 487826 92898 488062 93134
rect 488146 92898 488382 93134
rect 487826 57218 488062 57454
rect 488146 57218 488382 57454
rect 487826 56898 488062 57134
rect 488146 56898 488382 57134
rect 487826 21218 488062 21454
rect 488146 21218 488382 21454
rect 487826 20898 488062 21134
rect 488146 20898 488382 21134
rect 487826 -1542 488062 -1306
rect 488146 -1542 488382 -1306
rect 487826 -1862 488062 -1626
rect 488146 -1862 488382 -1626
rect 491546 672938 491782 673174
rect 491866 672938 492102 673174
rect 491546 672618 491782 672854
rect 491866 672618 492102 672854
rect 491546 636938 491782 637174
rect 491866 636938 492102 637174
rect 491546 636618 491782 636854
rect 491866 636618 492102 636854
rect 491546 600938 491782 601174
rect 491866 600938 492102 601174
rect 491546 600618 491782 600854
rect 491866 600618 492102 600854
rect 491546 564938 491782 565174
rect 491866 564938 492102 565174
rect 491546 564618 491782 564854
rect 491866 564618 492102 564854
rect 491546 528938 491782 529174
rect 491866 528938 492102 529174
rect 491546 528618 491782 528854
rect 491866 528618 492102 528854
rect 491546 492938 491782 493174
rect 491866 492938 492102 493174
rect 491546 492618 491782 492854
rect 491866 492618 492102 492854
rect 491546 456938 491782 457174
rect 491866 456938 492102 457174
rect 491546 456618 491782 456854
rect 491866 456618 492102 456854
rect 491546 420938 491782 421174
rect 491866 420938 492102 421174
rect 491546 420618 491782 420854
rect 491866 420618 492102 420854
rect 491546 384938 491782 385174
rect 491866 384938 492102 385174
rect 491546 384618 491782 384854
rect 491866 384618 492102 384854
rect 491546 348938 491782 349174
rect 491866 348938 492102 349174
rect 491546 348618 491782 348854
rect 491866 348618 492102 348854
rect 491546 312938 491782 313174
rect 491866 312938 492102 313174
rect 491546 312618 491782 312854
rect 491866 312618 492102 312854
rect 491546 276938 491782 277174
rect 491866 276938 492102 277174
rect 491546 276618 491782 276854
rect 491866 276618 492102 276854
rect 491546 240938 491782 241174
rect 491866 240938 492102 241174
rect 491546 240618 491782 240854
rect 491866 240618 492102 240854
rect 491546 204938 491782 205174
rect 491866 204938 492102 205174
rect 491546 204618 491782 204854
rect 491866 204618 492102 204854
rect 491546 168938 491782 169174
rect 491866 168938 492102 169174
rect 491546 168618 491782 168854
rect 491866 168618 492102 168854
rect 491546 132938 491782 133174
rect 491866 132938 492102 133174
rect 491546 132618 491782 132854
rect 491866 132618 492102 132854
rect 491546 96938 491782 97174
rect 491866 96938 492102 97174
rect 491546 96618 491782 96854
rect 491866 96618 492102 96854
rect 491546 60938 491782 61174
rect 491866 60938 492102 61174
rect 491546 60618 491782 60854
rect 491866 60618 492102 60854
rect 491546 24938 491782 25174
rect 491866 24938 492102 25174
rect 491546 24618 491782 24854
rect 491866 24618 492102 24854
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 676658 495502 676894
rect 495586 676658 495822 676894
rect 495266 676338 495502 676574
rect 495586 676338 495822 676574
rect 495266 640658 495502 640894
rect 495586 640658 495822 640894
rect 495266 640338 495502 640574
rect 495586 640338 495822 640574
rect 495266 604658 495502 604894
rect 495586 604658 495822 604894
rect 495266 604338 495502 604574
rect 495586 604338 495822 604574
rect 495266 568658 495502 568894
rect 495586 568658 495822 568894
rect 495266 568338 495502 568574
rect 495586 568338 495822 568574
rect 495266 532658 495502 532894
rect 495586 532658 495822 532894
rect 495266 532338 495502 532574
rect 495586 532338 495822 532574
rect 495266 496658 495502 496894
rect 495586 496658 495822 496894
rect 495266 496338 495502 496574
rect 495586 496338 495822 496574
rect 495266 460658 495502 460894
rect 495586 460658 495822 460894
rect 495266 460338 495502 460574
rect 495586 460338 495822 460574
rect 495266 424658 495502 424894
rect 495586 424658 495822 424894
rect 495266 424338 495502 424574
rect 495586 424338 495822 424574
rect 495266 388658 495502 388894
rect 495586 388658 495822 388894
rect 495266 388338 495502 388574
rect 495586 388338 495822 388574
rect 495266 352658 495502 352894
rect 495586 352658 495822 352894
rect 495266 352338 495502 352574
rect 495586 352338 495822 352574
rect 495266 316658 495502 316894
rect 495586 316658 495822 316894
rect 495266 316338 495502 316574
rect 495586 316338 495822 316574
rect 495266 280658 495502 280894
rect 495586 280658 495822 280894
rect 495266 280338 495502 280574
rect 495586 280338 495822 280574
rect 495266 244658 495502 244894
rect 495586 244658 495822 244894
rect 495266 244338 495502 244574
rect 495586 244338 495822 244574
rect 495266 208658 495502 208894
rect 495586 208658 495822 208894
rect 495266 208338 495502 208574
rect 495586 208338 495822 208574
rect 495266 172658 495502 172894
rect 495586 172658 495822 172894
rect 495266 172338 495502 172574
rect 495586 172338 495822 172574
rect 495266 136658 495502 136894
rect 495586 136658 495822 136894
rect 495266 136338 495502 136574
rect 495586 136338 495822 136574
rect 495266 100658 495502 100894
rect 495586 100658 495822 100894
rect 495266 100338 495502 100574
rect 495586 100338 495822 100574
rect 495266 64658 495502 64894
rect 495586 64658 495822 64894
rect 495266 64338 495502 64574
rect 495586 64338 495822 64574
rect 495266 28658 495502 28894
rect 495586 28658 495822 28894
rect 495266 28338 495502 28574
rect 495586 28338 495822 28574
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 498986 680378 499222 680614
rect 499306 680378 499542 680614
rect 498986 680058 499222 680294
rect 499306 680058 499542 680294
rect 498986 644378 499222 644614
rect 499306 644378 499542 644614
rect 498986 644058 499222 644294
rect 499306 644058 499542 644294
rect 498986 608378 499222 608614
rect 499306 608378 499542 608614
rect 498986 608058 499222 608294
rect 499306 608058 499542 608294
rect 498986 572378 499222 572614
rect 499306 572378 499542 572614
rect 498986 572058 499222 572294
rect 499306 572058 499542 572294
rect 498986 536378 499222 536614
rect 499306 536378 499542 536614
rect 498986 536058 499222 536294
rect 499306 536058 499542 536294
rect 498986 500378 499222 500614
rect 499306 500378 499542 500614
rect 498986 500058 499222 500294
rect 499306 500058 499542 500294
rect 498986 464378 499222 464614
rect 499306 464378 499542 464614
rect 498986 464058 499222 464294
rect 499306 464058 499542 464294
rect 498986 428378 499222 428614
rect 499306 428378 499542 428614
rect 498986 428058 499222 428294
rect 499306 428058 499542 428294
rect 498986 392378 499222 392614
rect 499306 392378 499542 392614
rect 498986 392058 499222 392294
rect 499306 392058 499542 392294
rect 498986 356378 499222 356614
rect 499306 356378 499542 356614
rect 498986 356058 499222 356294
rect 499306 356058 499542 356294
rect 498986 320378 499222 320614
rect 499306 320378 499542 320614
rect 498986 320058 499222 320294
rect 499306 320058 499542 320294
rect 498986 284378 499222 284614
rect 499306 284378 499542 284614
rect 498986 284058 499222 284294
rect 499306 284058 499542 284294
rect 498986 248378 499222 248614
rect 499306 248378 499542 248614
rect 498986 248058 499222 248294
rect 499306 248058 499542 248294
rect 498986 212378 499222 212614
rect 499306 212378 499542 212614
rect 498986 212058 499222 212294
rect 499306 212058 499542 212294
rect 498986 176378 499222 176614
rect 499306 176378 499542 176614
rect 498986 176058 499222 176294
rect 499306 176058 499542 176294
rect 498986 140378 499222 140614
rect 499306 140378 499542 140614
rect 498986 140058 499222 140294
rect 499306 140058 499542 140294
rect 498986 104378 499222 104614
rect 499306 104378 499542 104614
rect 498986 104058 499222 104294
rect 499306 104058 499542 104294
rect 498986 68378 499222 68614
rect 499306 68378 499542 68614
rect 498986 68058 499222 68294
rect 499306 68058 499542 68294
rect 498986 32378 499222 32614
rect 499306 32378 499542 32614
rect 498986 32058 499222 32294
rect 499306 32058 499542 32294
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 505826 687218 506062 687454
rect 506146 687218 506382 687454
rect 505826 686898 506062 687134
rect 506146 686898 506382 687134
rect 505826 651218 506062 651454
rect 506146 651218 506382 651454
rect 505826 650898 506062 651134
rect 506146 650898 506382 651134
rect 505826 615218 506062 615454
rect 506146 615218 506382 615454
rect 505826 614898 506062 615134
rect 506146 614898 506382 615134
rect 505826 579218 506062 579454
rect 506146 579218 506382 579454
rect 505826 578898 506062 579134
rect 506146 578898 506382 579134
rect 505826 543218 506062 543454
rect 506146 543218 506382 543454
rect 505826 542898 506062 543134
rect 506146 542898 506382 543134
rect 505826 507218 506062 507454
rect 506146 507218 506382 507454
rect 505826 506898 506062 507134
rect 506146 506898 506382 507134
rect 505826 471218 506062 471454
rect 506146 471218 506382 471454
rect 505826 470898 506062 471134
rect 506146 470898 506382 471134
rect 505826 435218 506062 435454
rect 506146 435218 506382 435454
rect 505826 434898 506062 435134
rect 506146 434898 506382 435134
rect 505826 399218 506062 399454
rect 506146 399218 506382 399454
rect 505826 398898 506062 399134
rect 506146 398898 506382 399134
rect 505826 363218 506062 363454
rect 506146 363218 506382 363454
rect 505826 362898 506062 363134
rect 506146 362898 506382 363134
rect 505826 327218 506062 327454
rect 506146 327218 506382 327454
rect 505826 326898 506062 327134
rect 506146 326898 506382 327134
rect 505826 291218 506062 291454
rect 506146 291218 506382 291454
rect 505826 290898 506062 291134
rect 506146 290898 506382 291134
rect 505826 255218 506062 255454
rect 506146 255218 506382 255454
rect 505826 254898 506062 255134
rect 506146 254898 506382 255134
rect 505826 219218 506062 219454
rect 506146 219218 506382 219454
rect 505826 218898 506062 219134
rect 506146 218898 506382 219134
rect 505826 183218 506062 183454
rect 506146 183218 506382 183454
rect 505826 182898 506062 183134
rect 506146 182898 506382 183134
rect 505826 147218 506062 147454
rect 506146 147218 506382 147454
rect 505826 146898 506062 147134
rect 506146 146898 506382 147134
rect 505826 111218 506062 111454
rect 506146 111218 506382 111454
rect 505826 110898 506062 111134
rect 506146 110898 506382 111134
rect 505826 75218 506062 75454
rect 506146 75218 506382 75454
rect 505826 74898 506062 75134
rect 506146 74898 506382 75134
rect 505826 39218 506062 39454
rect 506146 39218 506382 39454
rect 505826 38898 506062 39134
rect 506146 38898 506382 39134
rect 505826 3218 506062 3454
rect 506146 3218 506382 3454
rect 505826 2898 506062 3134
rect 506146 2898 506382 3134
rect 505826 -582 506062 -346
rect 506146 -582 506382 -346
rect 505826 -902 506062 -666
rect 506146 -902 506382 -666
rect 509546 690938 509782 691174
rect 509866 690938 510102 691174
rect 509546 690618 509782 690854
rect 509866 690618 510102 690854
rect 509546 654938 509782 655174
rect 509866 654938 510102 655174
rect 509546 654618 509782 654854
rect 509866 654618 510102 654854
rect 509546 618938 509782 619174
rect 509866 618938 510102 619174
rect 509546 618618 509782 618854
rect 509866 618618 510102 618854
rect 509546 582938 509782 583174
rect 509866 582938 510102 583174
rect 509546 582618 509782 582854
rect 509866 582618 510102 582854
rect 509546 546938 509782 547174
rect 509866 546938 510102 547174
rect 509546 546618 509782 546854
rect 509866 546618 510102 546854
rect 509546 510938 509782 511174
rect 509866 510938 510102 511174
rect 509546 510618 509782 510854
rect 509866 510618 510102 510854
rect 509546 474938 509782 475174
rect 509866 474938 510102 475174
rect 509546 474618 509782 474854
rect 509866 474618 510102 474854
rect 509546 438938 509782 439174
rect 509866 438938 510102 439174
rect 509546 438618 509782 438854
rect 509866 438618 510102 438854
rect 509546 402938 509782 403174
rect 509866 402938 510102 403174
rect 509546 402618 509782 402854
rect 509866 402618 510102 402854
rect 509546 366938 509782 367174
rect 509866 366938 510102 367174
rect 509546 366618 509782 366854
rect 509866 366618 510102 366854
rect 509546 330938 509782 331174
rect 509866 330938 510102 331174
rect 509546 330618 509782 330854
rect 509866 330618 510102 330854
rect 509546 294938 509782 295174
rect 509866 294938 510102 295174
rect 509546 294618 509782 294854
rect 509866 294618 510102 294854
rect 509546 258938 509782 259174
rect 509866 258938 510102 259174
rect 509546 258618 509782 258854
rect 509866 258618 510102 258854
rect 509546 222938 509782 223174
rect 509866 222938 510102 223174
rect 509546 222618 509782 222854
rect 509866 222618 510102 222854
rect 509546 186938 509782 187174
rect 509866 186938 510102 187174
rect 509546 186618 509782 186854
rect 509866 186618 510102 186854
rect 509546 150938 509782 151174
rect 509866 150938 510102 151174
rect 509546 150618 509782 150854
rect 509866 150618 510102 150854
rect 509546 114938 509782 115174
rect 509866 114938 510102 115174
rect 509546 114618 509782 114854
rect 509866 114618 510102 114854
rect 509546 78938 509782 79174
rect 509866 78938 510102 79174
rect 509546 78618 509782 78854
rect 509866 78618 510102 78854
rect 509546 42938 509782 43174
rect 509866 42938 510102 43174
rect 509546 42618 509782 42854
rect 509866 42618 510102 42854
rect 509546 6938 509782 7174
rect 509866 6938 510102 7174
rect 509546 6618 509782 6854
rect 509866 6618 510102 6854
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 694658 513502 694894
rect 513586 694658 513822 694894
rect 513266 694338 513502 694574
rect 513586 694338 513822 694574
rect 513266 658658 513502 658894
rect 513586 658658 513822 658894
rect 513266 658338 513502 658574
rect 513586 658338 513822 658574
rect 513266 622658 513502 622894
rect 513586 622658 513822 622894
rect 513266 622338 513502 622574
rect 513586 622338 513822 622574
rect 513266 586658 513502 586894
rect 513586 586658 513822 586894
rect 513266 586338 513502 586574
rect 513586 586338 513822 586574
rect 513266 550658 513502 550894
rect 513586 550658 513822 550894
rect 513266 550338 513502 550574
rect 513586 550338 513822 550574
rect 513266 514658 513502 514894
rect 513586 514658 513822 514894
rect 513266 514338 513502 514574
rect 513586 514338 513822 514574
rect 513266 478658 513502 478894
rect 513586 478658 513822 478894
rect 513266 478338 513502 478574
rect 513586 478338 513822 478574
rect 513266 442658 513502 442894
rect 513586 442658 513822 442894
rect 513266 442338 513502 442574
rect 513586 442338 513822 442574
rect 513266 406658 513502 406894
rect 513586 406658 513822 406894
rect 513266 406338 513502 406574
rect 513586 406338 513822 406574
rect 513266 370658 513502 370894
rect 513586 370658 513822 370894
rect 513266 370338 513502 370574
rect 513586 370338 513822 370574
rect 513266 334658 513502 334894
rect 513586 334658 513822 334894
rect 513266 334338 513502 334574
rect 513586 334338 513822 334574
rect 513266 298658 513502 298894
rect 513586 298658 513822 298894
rect 513266 298338 513502 298574
rect 513586 298338 513822 298574
rect 513266 262658 513502 262894
rect 513586 262658 513822 262894
rect 513266 262338 513502 262574
rect 513586 262338 513822 262574
rect 513266 226658 513502 226894
rect 513586 226658 513822 226894
rect 513266 226338 513502 226574
rect 513586 226338 513822 226574
rect 513266 190658 513502 190894
rect 513586 190658 513822 190894
rect 513266 190338 513502 190574
rect 513586 190338 513822 190574
rect 513266 154658 513502 154894
rect 513586 154658 513822 154894
rect 513266 154338 513502 154574
rect 513586 154338 513822 154574
rect 513266 118658 513502 118894
rect 513586 118658 513822 118894
rect 513266 118338 513502 118574
rect 513586 118338 513822 118574
rect 513266 82658 513502 82894
rect 513586 82658 513822 82894
rect 513266 82338 513502 82574
rect 513586 82338 513822 82574
rect 513266 46658 513502 46894
rect 513586 46658 513822 46894
rect 513266 46338 513502 46574
rect 513586 46338 513822 46574
rect 513266 10658 513502 10894
rect 513586 10658 513822 10894
rect 513266 10338 513502 10574
rect 513586 10338 513822 10574
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 516986 698378 517222 698614
rect 517306 698378 517542 698614
rect 516986 698058 517222 698294
rect 517306 698058 517542 698294
rect 516986 662378 517222 662614
rect 517306 662378 517542 662614
rect 516986 662058 517222 662294
rect 517306 662058 517542 662294
rect 516986 626378 517222 626614
rect 517306 626378 517542 626614
rect 516986 626058 517222 626294
rect 517306 626058 517542 626294
rect 516986 590378 517222 590614
rect 517306 590378 517542 590614
rect 516986 590058 517222 590294
rect 517306 590058 517542 590294
rect 516986 554378 517222 554614
rect 517306 554378 517542 554614
rect 516986 554058 517222 554294
rect 517306 554058 517542 554294
rect 516986 518378 517222 518614
rect 517306 518378 517542 518614
rect 516986 518058 517222 518294
rect 517306 518058 517542 518294
rect 516986 482378 517222 482614
rect 517306 482378 517542 482614
rect 516986 482058 517222 482294
rect 517306 482058 517542 482294
rect 516986 446378 517222 446614
rect 517306 446378 517542 446614
rect 516986 446058 517222 446294
rect 517306 446058 517542 446294
rect 516986 410378 517222 410614
rect 517306 410378 517542 410614
rect 516986 410058 517222 410294
rect 517306 410058 517542 410294
rect 516986 374378 517222 374614
rect 517306 374378 517542 374614
rect 516986 374058 517222 374294
rect 517306 374058 517542 374294
rect 516986 338378 517222 338614
rect 517306 338378 517542 338614
rect 516986 338058 517222 338294
rect 517306 338058 517542 338294
rect 516986 302378 517222 302614
rect 517306 302378 517542 302614
rect 516986 302058 517222 302294
rect 517306 302058 517542 302294
rect 516986 266378 517222 266614
rect 517306 266378 517542 266614
rect 516986 266058 517222 266294
rect 517306 266058 517542 266294
rect 516986 230378 517222 230614
rect 517306 230378 517542 230614
rect 516986 230058 517222 230294
rect 517306 230058 517542 230294
rect 516986 194378 517222 194614
rect 517306 194378 517542 194614
rect 516986 194058 517222 194294
rect 517306 194058 517542 194294
rect 516986 158378 517222 158614
rect 517306 158378 517542 158614
rect 516986 158058 517222 158294
rect 517306 158058 517542 158294
rect 516986 122378 517222 122614
rect 517306 122378 517542 122614
rect 516986 122058 517222 122294
rect 517306 122058 517542 122294
rect 516986 86378 517222 86614
rect 517306 86378 517542 86614
rect 516986 86058 517222 86294
rect 517306 86058 517542 86294
rect 516986 50378 517222 50614
rect 517306 50378 517542 50614
rect 516986 50058 517222 50294
rect 517306 50058 517542 50294
rect 516986 14378 517222 14614
rect 517306 14378 517542 14614
rect 516986 14058 517222 14294
rect 517306 14058 517542 14294
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 523826 669218 524062 669454
rect 524146 669218 524382 669454
rect 523826 668898 524062 669134
rect 524146 668898 524382 669134
rect 523826 633218 524062 633454
rect 524146 633218 524382 633454
rect 523826 632898 524062 633134
rect 524146 632898 524382 633134
rect 523826 597218 524062 597454
rect 524146 597218 524382 597454
rect 523826 596898 524062 597134
rect 524146 596898 524382 597134
rect 523826 561218 524062 561454
rect 524146 561218 524382 561454
rect 523826 560898 524062 561134
rect 524146 560898 524382 561134
rect 523826 525218 524062 525454
rect 524146 525218 524382 525454
rect 523826 524898 524062 525134
rect 524146 524898 524382 525134
rect 523826 489218 524062 489454
rect 524146 489218 524382 489454
rect 523826 488898 524062 489134
rect 524146 488898 524382 489134
rect 523826 453218 524062 453454
rect 524146 453218 524382 453454
rect 523826 452898 524062 453134
rect 524146 452898 524382 453134
rect 523826 417218 524062 417454
rect 524146 417218 524382 417454
rect 523826 416898 524062 417134
rect 524146 416898 524382 417134
rect 523826 381218 524062 381454
rect 524146 381218 524382 381454
rect 523826 380898 524062 381134
rect 524146 380898 524382 381134
rect 523826 345218 524062 345454
rect 524146 345218 524382 345454
rect 523826 344898 524062 345134
rect 524146 344898 524382 345134
rect 523826 309218 524062 309454
rect 524146 309218 524382 309454
rect 523826 308898 524062 309134
rect 524146 308898 524382 309134
rect 523826 273218 524062 273454
rect 524146 273218 524382 273454
rect 523826 272898 524062 273134
rect 524146 272898 524382 273134
rect 523826 237218 524062 237454
rect 524146 237218 524382 237454
rect 523826 236898 524062 237134
rect 524146 236898 524382 237134
rect 523826 201218 524062 201454
rect 524146 201218 524382 201454
rect 523826 200898 524062 201134
rect 524146 200898 524382 201134
rect 523826 165218 524062 165454
rect 524146 165218 524382 165454
rect 523826 164898 524062 165134
rect 524146 164898 524382 165134
rect 523826 129218 524062 129454
rect 524146 129218 524382 129454
rect 523826 128898 524062 129134
rect 524146 128898 524382 129134
rect 523826 93218 524062 93454
rect 524146 93218 524382 93454
rect 523826 92898 524062 93134
rect 524146 92898 524382 93134
rect 523826 57218 524062 57454
rect 524146 57218 524382 57454
rect 523826 56898 524062 57134
rect 524146 56898 524382 57134
rect 523826 21218 524062 21454
rect 524146 21218 524382 21454
rect 523826 20898 524062 21134
rect 524146 20898 524382 21134
rect 523826 -1542 524062 -1306
rect 524146 -1542 524382 -1306
rect 523826 -1862 524062 -1626
rect 524146 -1862 524382 -1626
rect 527546 672938 527782 673174
rect 527866 672938 528102 673174
rect 527546 672618 527782 672854
rect 527866 672618 528102 672854
rect 527546 636938 527782 637174
rect 527866 636938 528102 637174
rect 527546 636618 527782 636854
rect 527866 636618 528102 636854
rect 527546 600938 527782 601174
rect 527866 600938 528102 601174
rect 527546 600618 527782 600854
rect 527866 600618 528102 600854
rect 527546 564938 527782 565174
rect 527866 564938 528102 565174
rect 527546 564618 527782 564854
rect 527866 564618 528102 564854
rect 527546 528938 527782 529174
rect 527866 528938 528102 529174
rect 527546 528618 527782 528854
rect 527866 528618 528102 528854
rect 527546 492938 527782 493174
rect 527866 492938 528102 493174
rect 527546 492618 527782 492854
rect 527866 492618 528102 492854
rect 527546 456938 527782 457174
rect 527866 456938 528102 457174
rect 527546 456618 527782 456854
rect 527866 456618 528102 456854
rect 527546 420938 527782 421174
rect 527866 420938 528102 421174
rect 527546 420618 527782 420854
rect 527866 420618 528102 420854
rect 527546 384938 527782 385174
rect 527866 384938 528102 385174
rect 527546 384618 527782 384854
rect 527866 384618 528102 384854
rect 527546 348938 527782 349174
rect 527866 348938 528102 349174
rect 527546 348618 527782 348854
rect 527866 348618 528102 348854
rect 527546 312938 527782 313174
rect 527866 312938 528102 313174
rect 527546 312618 527782 312854
rect 527866 312618 528102 312854
rect 527546 276938 527782 277174
rect 527866 276938 528102 277174
rect 527546 276618 527782 276854
rect 527866 276618 528102 276854
rect 527546 240938 527782 241174
rect 527866 240938 528102 241174
rect 527546 240618 527782 240854
rect 527866 240618 528102 240854
rect 527546 204938 527782 205174
rect 527866 204938 528102 205174
rect 527546 204618 527782 204854
rect 527866 204618 528102 204854
rect 527546 168938 527782 169174
rect 527866 168938 528102 169174
rect 527546 168618 527782 168854
rect 527866 168618 528102 168854
rect 527546 132938 527782 133174
rect 527866 132938 528102 133174
rect 527546 132618 527782 132854
rect 527866 132618 528102 132854
rect 527546 96938 527782 97174
rect 527866 96938 528102 97174
rect 527546 96618 527782 96854
rect 527866 96618 528102 96854
rect 527546 60938 527782 61174
rect 527866 60938 528102 61174
rect 527546 60618 527782 60854
rect 527866 60618 528102 60854
rect 527546 24938 527782 25174
rect 527866 24938 528102 25174
rect 527546 24618 527782 24854
rect 527866 24618 528102 24854
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 676658 531502 676894
rect 531586 676658 531822 676894
rect 531266 676338 531502 676574
rect 531586 676338 531822 676574
rect 531266 640658 531502 640894
rect 531586 640658 531822 640894
rect 531266 640338 531502 640574
rect 531586 640338 531822 640574
rect 531266 604658 531502 604894
rect 531586 604658 531822 604894
rect 531266 604338 531502 604574
rect 531586 604338 531822 604574
rect 531266 568658 531502 568894
rect 531586 568658 531822 568894
rect 531266 568338 531502 568574
rect 531586 568338 531822 568574
rect 531266 532658 531502 532894
rect 531586 532658 531822 532894
rect 531266 532338 531502 532574
rect 531586 532338 531822 532574
rect 531266 496658 531502 496894
rect 531586 496658 531822 496894
rect 531266 496338 531502 496574
rect 531586 496338 531822 496574
rect 531266 460658 531502 460894
rect 531586 460658 531822 460894
rect 531266 460338 531502 460574
rect 531586 460338 531822 460574
rect 531266 424658 531502 424894
rect 531586 424658 531822 424894
rect 531266 424338 531502 424574
rect 531586 424338 531822 424574
rect 531266 388658 531502 388894
rect 531586 388658 531822 388894
rect 531266 388338 531502 388574
rect 531586 388338 531822 388574
rect 531266 352658 531502 352894
rect 531586 352658 531822 352894
rect 531266 352338 531502 352574
rect 531586 352338 531822 352574
rect 531266 316658 531502 316894
rect 531586 316658 531822 316894
rect 531266 316338 531502 316574
rect 531586 316338 531822 316574
rect 531266 280658 531502 280894
rect 531586 280658 531822 280894
rect 531266 280338 531502 280574
rect 531586 280338 531822 280574
rect 531266 244658 531502 244894
rect 531586 244658 531822 244894
rect 531266 244338 531502 244574
rect 531586 244338 531822 244574
rect 531266 208658 531502 208894
rect 531586 208658 531822 208894
rect 531266 208338 531502 208574
rect 531586 208338 531822 208574
rect 531266 172658 531502 172894
rect 531586 172658 531822 172894
rect 531266 172338 531502 172574
rect 531586 172338 531822 172574
rect 531266 136658 531502 136894
rect 531586 136658 531822 136894
rect 531266 136338 531502 136574
rect 531586 136338 531822 136574
rect 531266 100658 531502 100894
rect 531586 100658 531822 100894
rect 531266 100338 531502 100574
rect 531586 100338 531822 100574
rect 531266 64658 531502 64894
rect 531586 64658 531822 64894
rect 531266 64338 531502 64574
rect 531586 64338 531822 64574
rect 531266 28658 531502 28894
rect 531586 28658 531822 28894
rect 531266 28338 531502 28574
rect 531586 28338 531822 28574
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 534986 680378 535222 680614
rect 535306 680378 535542 680614
rect 534986 680058 535222 680294
rect 535306 680058 535542 680294
rect 534986 644378 535222 644614
rect 535306 644378 535542 644614
rect 534986 644058 535222 644294
rect 535306 644058 535542 644294
rect 534986 608378 535222 608614
rect 535306 608378 535542 608614
rect 534986 608058 535222 608294
rect 535306 608058 535542 608294
rect 534986 572378 535222 572614
rect 535306 572378 535542 572614
rect 534986 572058 535222 572294
rect 535306 572058 535542 572294
rect 534986 536378 535222 536614
rect 535306 536378 535542 536614
rect 534986 536058 535222 536294
rect 535306 536058 535542 536294
rect 534986 500378 535222 500614
rect 535306 500378 535542 500614
rect 534986 500058 535222 500294
rect 535306 500058 535542 500294
rect 534986 464378 535222 464614
rect 535306 464378 535542 464614
rect 534986 464058 535222 464294
rect 535306 464058 535542 464294
rect 534986 428378 535222 428614
rect 535306 428378 535542 428614
rect 534986 428058 535222 428294
rect 535306 428058 535542 428294
rect 534986 392378 535222 392614
rect 535306 392378 535542 392614
rect 534986 392058 535222 392294
rect 535306 392058 535542 392294
rect 534986 356378 535222 356614
rect 535306 356378 535542 356614
rect 534986 356058 535222 356294
rect 535306 356058 535542 356294
rect 534986 320378 535222 320614
rect 535306 320378 535542 320614
rect 534986 320058 535222 320294
rect 535306 320058 535542 320294
rect 534986 284378 535222 284614
rect 535306 284378 535542 284614
rect 534986 284058 535222 284294
rect 535306 284058 535542 284294
rect 534986 248378 535222 248614
rect 535306 248378 535542 248614
rect 534986 248058 535222 248294
rect 535306 248058 535542 248294
rect 534986 212378 535222 212614
rect 535306 212378 535542 212614
rect 534986 212058 535222 212294
rect 535306 212058 535542 212294
rect 534986 176378 535222 176614
rect 535306 176378 535542 176614
rect 534986 176058 535222 176294
rect 535306 176058 535542 176294
rect 534986 140378 535222 140614
rect 535306 140378 535542 140614
rect 534986 140058 535222 140294
rect 535306 140058 535542 140294
rect 534986 104378 535222 104614
rect 535306 104378 535542 104614
rect 534986 104058 535222 104294
rect 535306 104058 535542 104294
rect 534986 68378 535222 68614
rect 535306 68378 535542 68614
rect 534986 68058 535222 68294
rect 535306 68058 535542 68294
rect 534986 32378 535222 32614
rect 535306 32378 535542 32614
rect 534986 32058 535222 32294
rect 535306 32058 535542 32294
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 541826 687218 542062 687454
rect 542146 687218 542382 687454
rect 541826 686898 542062 687134
rect 542146 686898 542382 687134
rect 541826 651218 542062 651454
rect 542146 651218 542382 651454
rect 541826 650898 542062 651134
rect 542146 650898 542382 651134
rect 541826 615218 542062 615454
rect 542146 615218 542382 615454
rect 541826 614898 542062 615134
rect 542146 614898 542382 615134
rect 541826 579218 542062 579454
rect 542146 579218 542382 579454
rect 541826 578898 542062 579134
rect 542146 578898 542382 579134
rect 541826 543218 542062 543454
rect 542146 543218 542382 543454
rect 541826 542898 542062 543134
rect 542146 542898 542382 543134
rect 541826 507218 542062 507454
rect 542146 507218 542382 507454
rect 541826 506898 542062 507134
rect 542146 506898 542382 507134
rect 541826 471218 542062 471454
rect 542146 471218 542382 471454
rect 541826 470898 542062 471134
rect 542146 470898 542382 471134
rect 541826 435218 542062 435454
rect 542146 435218 542382 435454
rect 541826 434898 542062 435134
rect 542146 434898 542382 435134
rect 541826 399218 542062 399454
rect 542146 399218 542382 399454
rect 541826 398898 542062 399134
rect 542146 398898 542382 399134
rect 541826 363218 542062 363454
rect 542146 363218 542382 363454
rect 541826 362898 542062 363134
rect 542146 362898 542382 363134
rect 541826 327218 542062 327454
rect 542146 327218 542382 327454
rect 541826 326898 542062 327134
rect 542146 326898 542382 327134
rect 541826 291218 542062 291454
rect 542146 291218 542382 291454
rect 541826 290898 542062 291134
rect 542146 290898 542382 291134
rect 541826 255218 542062 255454
rect 542146 255218 542382 255454
rect 541826 254898 542062 255134
rect 542146 254898 542382 255134
rect 541826 219218 542062 219454
rect 542146 219218 542382 219454
rect 541826 218898 542062 219134
rect 542146 218898 542382 219134
rect 541826 183218 542062 183454
rect 542146 183218 542382 183454
rect 541826 182898 542062 183134
rect 542146 182898 542382 183134
rect 541826 147218 542062 147454
rect 542146 147218 542382 147454
rect 541826 146898 542062 147134
rect 542146 146898 542382 147134
rect 541826 111218 542062 111454
rect 542146 111218 542382 111454
rect 541826 110898 542062 111134
rect 542146 110898 542382 111134
rect 541826 75218 542062 75454
rect 542146 75218 542382 75454
rect 541826 74898 542062 75134
rect 542146 74898 542382 75134
rect 541826 39218 542062 39454
rect 542146 39218 542382 39454
rect 541826 38898 542062 39134
rect 542146 38898 542382 39134
rect 541826 3218 542062 3454
rect 542146 3218 542382 3454
rect 541826 2898 542062 3134
rect 542146 2898 542382 3134
rect 541826 -582 542062 -346
rect 542146 -582 542382 -346
rect 541826 -902 542062 -666
rect 542146 -902 542382 -666
rect 545546 690938 545782 691174
rect 545866 690938 546102 691174
rect 545546 690618 545782 690854
rect 545866 690618 546102 690854
rect 545546 654938 545782 655174
rect 545866 654938 546102 655174
rect 545546 654618 545782 654854
rect 545866 654618 546102 654854
rect 545546 618938 545782 619174
rect 545866 618938 546102 619174
rect 545546 618618 545782 618854
rect 545866 618618 546102 618854
rect 545546 582938 545782 583174
rect 545866 582938 546102 583174
rect 545546 582618 545782 582854
rect 545866 582618 546102 582854
rect 545546 546938 545782 547174
rect 545866 546938 546102 547174
rect 545546 546618 545782 546854
rect 545866 546618 546102 546854
rect 545546 510938 545782 511174
rect 545866 510938 546102 511174
rect 545546 510618 545782 510854
rect 545866 510618 546102 510854
rect 545546 474938 545782 475174
rect 545866 474938 546102 475174
rect 545546 474618 545782 474854
rect 545866 474618 546102 474854
rect 545546 438938 545782 439174
rect 545866 438938 546102 439174
rect 545546 438618 545782 438854
rect 545866 438618 546102 438854
rect 545546 402938 545782 403174
rect 545866 402938 546102 403174
rect 545546 402618 545782 402854
rect 545866 402618 546102 402854
rect 545546 366938 545782 367174
rect 545866 366938 546102 367174
rect 545546 366618 545782 366854
rect 545866 366618 546102 366854
rect 545546 330938 545782 331174
rect 545866 330938 546102 331174
rect 545546 330618 545782 330854
rect 545866 330618 546102 330854
rect 545546 294938 545782 295174
rect 545866 294938 546102 295174
rect 545546 294618 545782 294854
rect 545866 294618 546102 294854
rect 545546 258938 545782 259174
rect 545866 258938 546102 259174
rect 545546 258618 545782 258854
rect 545866 258618 546102 258854
rect 545546 222938 545782 223174
rect 545866 222938 546102 223174
rect 545546 222618 545782 222854
rect 545866 222618 546102 222854
rect 545546 186938 545782 187174
rect 545866 186938 546102 187174
rect 545546 186618 545782 186854
rect 545866 186618 546102 186854
rect 545546 150938 545782 151174
rect 545866 150938 546102 151174
rect 545546 150618 545782 150854
rect 545866 150618 546102 150854
rect 545546 114938 545782 115174
rect 545866 114938 546102 115174
rect 545546 114618 545782 114854
rect 545866 114618 546102 114854
rect 545546 78938 545782 79174
rect 545866 78938 546102 79174
rect 545546 78618 545782 78854
rect 545866 78618 546102 78854
rect 545546 42938 545782 43174
rect 545866 42938 546102 43174
rect 545546 42618 545782 42854
rect 545866 42618 546102 42854
rect 545546 6938 545782 7174
rect 545866 6938 546102 7174
rect 545546 6618 545782 6854
rect 545866 6618 546102 6854
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 694658 549502 694894
rect 549586 694658 549822 694894
rect 549266 694338 549502 694574
rect 549586 694338 549822 694574
rect 549266 658658 549502 658894
rect 549586 658658 549822 658894
rect 549266 658338 549502 658574
rect 549586 658338 549822 658574
rect 549266 622658 549502 622894
rect 549586 622658 549822 622894
rect 549266 622338 549502 622574
rect 549586 622338 549822 622574
rect 549266 586658 549502 586894
rect 549586 586658 549822 586894
rect 549266 586338 549502 586574
rect 549586 586338 549822 586574
rect 549266 550658 549502 550894
rect 549586 550658 549822 550894
rect 549266 550338 549502 550574
rect 549586 550338 549822 550574
rect 549266 514658 549502 514894
rect 549586 514658 549822 514894
rect 549266 514338 549502 514574
rect 549586 514338 549822 514574
rect 549266 478658 549502 478894
rect 549586 478658 549822 478894
rect 549266 478338 549502 478574
rect 549586 478338 549822 478574
rect 549266 442658 549502 442894
rect 549586 442658 549822 442894
rect 549266 442338 549502 442574
rect 549586 442338 549822 442574
rect 549266 406658 549502 406894
rect 549586 406658 549822 406894
rect 549266 406338 549502 406574
rect 549586 406338 549822 406574
rect 549266 370658 549502 370894
rect 549586 370658 549822 370894
rect 549266 370338 549502 370574
rect 549586 370338 549822 370574
rect 549266 334658 549502 334894
rect 549586 334658 549822 334894
rect 549266 334338 549502 334574
rect 549586 334338 549822 334574
rect 549266 298658 549502 298894
rect 549586 298658 549822 298894
rect 549266 298338 549502 298574
rect 549586 298338 549822 298574
rect 549266 262658 549502 262894
rect 549586 262658 549822 262894
rect 549266 262338 549502 262574
rect 549586 262338 549822 262574
rect 549266 226658 549502 226894
rect 549586 226658 549822 226894
rect 549266 226338 549502 226574
rect 549586 226338 549822 226574
rect 549266 190658 549502 190894
rect 549586 190658 549822 190894
rect 549266 190338 549502 190574
rect 549586 190338 549822 190574
rect 549266 154658 549502 154894
rect 549586 154658 549822 154894
rect 549266 154338 549502 154574
rect 549586 154338 549822 154574
rect 549266 118658 549502 118894
rect 549586 118658 549822 118894
rect 549266 118338 549502 118574
rect 549586 118338 549822 118574
rect 549266 82658 549502 82894
rect 549586 82658 549822 82894
rect 549266 82338 549502 82574
rect 549586 82338 549822 82574
rect 549266 46658 549502 46894
rect 549586 46658 549822 46894
rect 549266 46338 549502 46574
rect 549586 46338 549822 46574
rect 549266 10658 549502 10894
rect 549586 10658 549822 10894
rect 549266 10338 549502 10574
rect 549586 10338 549822 10574
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 552986 698378 553222 698614
rect 553306 698378 553542 698614
rect 552986 698058 553222 698294
rect 553306 698058 553542 698294
rect 552986 662378 553222 662614
rect 553306 662378 553542 662614
rect 552986 662058 553222 662294
rect 553306 662058 553542 662294
rect 552986 626378 553222 626614
rect 553306 626378 553542 626614
rect 552986 626058 553222 626294
rect 553306 626058 553542 626294
rect 552986 590378 553222 590614
rect 553306 590378 553542 590614
rect 552986 590058 553222 590294
rect 553306 590058 553542 590294
rect 552986 554378 553222 554614
rect 553306 554378 553542 554614
rect 552986 554058 553222 554294
rect 553306 554058 553542 554294
rect 552986 518378 553222 518614
rect 553306 518378 553542 518614
rect 552986 518058 553222 518294
rect 553306 518058 553542 518294
rect 552986 482378 553222 482614
rect 553306 482378 553542 482614
rect 552986 482058 553222 482294
rect 553306 482058 553542 482294
rect 552986 446378 553222 446614
rect 553306 446378 553542 446614
rect 552986 446058 553222 446294
rect 553306 446058 553542 446294
rect 552986 410378 553222 410614
rect 553306 410378 553542 410614
rect 552986 410058 553222 410294
rect 553306 410058 553542 410294
rect 552986 374378 553222 374614
rect 553306 374378 553542 374614
rect 552986 374058 553222 374294
rect 553306 374058 553542 374294
rect 552986 338378 553222 338614
rect 553306 338378 553542 338614
rect 552986 338058 553222 338294
rect 553306 338058 553542 338294
rect 552986 302378 553222 302614
rect 553306 302378 553542 302614
rect 552986 302058 553222 302294
rect 553306 302058 553542 302294
rect 552986 266378 553222 266614
rect 553306 266378 553542 266614
rect 552986 266058 553222 266294
rect 553306 266058 553542 266294
rect 552986 230378 553222 230614
rect 553306 230378 553542 230614
rect 552986 230058 553222 230294
rect 553306 230058 553542 230294
rect 552986 194378 553222 194614
rect 553306 194378 553542 194614
rect 552986 194058 553222 194294
rect 553306 194058 553542 194294
rect 552986 158378 553222 158614
rect 553306 158378 553542 158614
rect 552986 158058 553222 158294
rect 553306 158058 553542 158294
rect 552986 122378 553222 122614
rect 553306 122378 553542 122614
rect 552986 122058 553222 122294
rect 553306 122058 553542 122294
rect 552986 86378 553222 86614
rect 553306 86378 553542 86614
rect 552986 86058 553222 86294
rect 553306 86058 553542 86294
rect 552986 50378 553222 50614
rect 553306 50378 553542 50614
rect 552986 50058 553222 50294
rect 553306 50058 553542 50294
rect 552986 14378 553222 14614
rect 553306 14378 553542 14614
rect 552986 14058 553222 14294
rect 553306 14058 553542 14294
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect 559826 669218 560062 669454
rect 560146 669218 560382 669454
rect 559826 668898 560062 669134
rect 560146 668898 560382 669134
rect 559826 633218 560062 633454
rect 560146 633218 560382 633454
rect 559826 632898 560062 633134
rect 560146 632898 560382 633134
rect 559826 597218 560062 597454
rect 560146 597218 560382 597454
rect 559826 596898 560062 597134
rect 560146 596898 560382 597134
rect 559826 561218 560062 561454
rect 560146 561218 560382 561454
rect 559826 560898 560062 561134
rect 560146 560898 560382 561134
rect 559826 525218 560062 525454
rect 560146 525218 560382 525454
rect 559826 524898 560062 525134
rect 560146 524898 560382 525134
rect 559826 489218 560062 489454
rect 560146 489218 560382 489454
rect 559826 488898 560062 489134
rect 560146 488898 560382 489134
rect 559826 453218 560062 453454
rect 560146 453218 560382 453454
rect 559826 452898 560062 453134
rect 560146 452898 560382 453134
rect 559826 417218 560062 417454
rect 560146 417218 560382 417454
rect 559826 416898 560062 417134
rect 560146 416898 560382 417134
rect 559826 381218 560062 381454
rect 560146 381218 560382 381454
rect 559826 380898 560062 381134
rect 560146 380898 560382 381134
rect 559826 345218 560062 345454
rect 560146 345218 560382 345454
rect 559826 344898 560062 345134
rect 560146 344898 560382 345134
rect 559826 309218 560062 309454
rect 560146 309218 560382 309454
rect 559826 308898 560062 309134
rect 560146 308898 560382 309134
rect 559826 273218 560062 273454
rect 560146 273218 560382 273454
rect 559826 272898 560062 273134
rect 560146 272898 560382 273134
rect 559826 237218 560062 237454
rect 560146 237218 560382 237454
rect 559826 236898 560062 237134
rect 560146 236898 560382 237134
rect 559826 201218 560062 201454
rect 560146 201218 560382 201454
rect 559826 200898 560062 201134
rect 560146 200898 560382 201134
rect 559826 165218 560062 165454
rect 560146 165218 560382 165454
rect 559826 164898 560062 165134
rect 560146 164898 560382 165134
rect 559826 129218 560062 129454
rect 560146 129218 560382 129454
rect 559826 128898 560062 129134
rect 560146 128898 560382 129134
rect 559826 93218 560062 93454
rect 560146 93218 560382 93454
rect 559826 92898 560062 93134
rect 560146 92898 560382 93134
rect 559826 57218 560062 57454
rect 560146 57218 560382 57454
rect 559826 56898 560062 57134
rect 560146 56898 560382 57134
rect 559826 21218 560062 21454
rect 560146 21218 560382 21454
rect 559826 20898 560062 21134
rect 560146 20898 560382 21134
rect 559826 -1542 560062 -1306
rect 560146 -1542 560382 -1306
rect 559826 -1862 560062 -1626
rect 560146 -1862 560382 -1626
rect 563546 672938 563782 673174
rect 563866 672938 564102 673174
rect 563546 672618 563782 672854
rect 563866 672618 564102 672854
rect 563546 636938 563782 637174
rect 563866 636938 564102 637174
rect 563546 636618 563782 636854
rect 563866 636618 564102 636854
rect 563546 600938 563782 601174
rect 563866 600938 564102 601174
rect 563546 600618 563782 600854
rect 563866 600618 564102 600854
rect 563546 564938 563782 565174
rect 563866 564938 564102 565174
rect 563546 564618 563782 564854
rect 563866 564618 564102 564854
rect 563546 528938 563782 529174
rect 563866 528938 564102 529174
rect 563546 528618 563782 528854
rect 563866 528618 564102 528854
rect 563546 492938 563782 493174
rect 563866 492938 564102 493174
rect 563546 492618 563782 492854
rect 563866 492618 564102 492854
rect 563546 456938 563782 457174
rect 563866 456938 564102 457174
rect 563546 456618 563782 456854
rect 563866 456618 564102 456854
rect 563546 420938 563782 421174
rect 563866 420938 564102 421174
rect 563546 420618 563782 420854
rect 563866 420618 564102 420854
rect 563546 384938 563782 385174
rect 563866 384938 564102 385174
rect 563546 384618 563782 384854
rect 563866 384618 564102 384854
rect 563546 348938 563782 349174
rect 563866 348938 564102 349174
rect 563546 348618 563782 348854
rect 563866 348618 564102 348854
rect 563546 312938 563782 313174
rect 563866 312938 564102 313174
rect 563546 312618 563782 312854
rect 563866 312618 564102 312854
rect 563546 276938 563782 277174
rect 563866 276938 564102 277174
rect 563546 276618 563782 276854
rect 563866 276618 564102 276854
rect 563546 240938 563782 241174
rect 563866 240938 564102 241174
rect 563546 240618 563782 240854
rect 563866 240618 564102 240854
rect 563546 204938 563782 205174
rect 563866 204938 564102 205174
rect 563546 204618 563782 204854
rect 563866 204618 564102 204854
rect 563546 168938 563782 169174
rect 563866 168938 564102 169174
rect 563546 168618 563782 168854
rect 563866 168618 564102 168854
rect 563546 132938 563782 133174
rect 563866 132938 564102 133174
rect 563546 132618 563782 132854
rect 563866 132618 564102 132854
rect 563546 96938 563782 97174
rect 563866 96938 564102 97174
rect 563546 96618 563782 96854
rect 563866 96618 564102 96854
rect 563546 60938 563782 61174
rect 563866 60938 564102 61174
rect 563546 60618 563782 60854
rect 563866 60618 564102 60854
rect 563546 24938 563782 25174
rect 563866 24938 564102 25174
rect 563546 24618 563782 24854
rect 563866 24618 564102 24854
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 12986 698614
rect 13222 698378 13306 698614
rect 13542 698378 48986 698614
rect 49222 698378 49306 698614
rect 49542 698378 84986 698614
rect 85222 698378 85306 698614
rect 85542 698378 120986 698614
rect 121222 698378 121306 698614
rect 121542 698378 156986 698614
rect 157222 698378 157306 698614
rect 157542 698378 192986 698614
rect 193222 698378 193306 698614
rect 193542 698378 228986 698614
rect 229222 698378 229306 698614
rect 229542 698378 264986 698614
rect 265222 698378 265306 698614
rect 265542 698378 300986 698614
rect 301222 698378 301306 698614
rect 301542 698378 336986 698614
rect 337222 698378 337306 698614
rect 337542 698378 372986 698614
rect 373222 698378 373306 698614
rect 373542 698378 408986 698614
rect 409222 698378 409306 698614
rect 409542 698378 444986 698614
rect 445222 698378 445306 698614
rect 445542 698378 480986 698614
rect 481222 698378 481306 698614
rect 481542 698378 516986 698614
rect 517222 698378 517306 698614
rect 517542 698378 552986 698614
rect 553222 698378 553306 698614
rect 553542 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 12986 698294
rect 13222 698058 13306 698294
rect 13542 698058 48986 698294
rect 49222 698058 49306 698294
rect 49542 698058 84986 698294
rect 85222 698058 85306 698294
rect 85542 698058 120986 698294
rect 121222 698058 121306 698294
rect 121542 698058 156986 698294
rect 157222 698058 157306 698294
rect 157542 698058 192986 698294
rect 193222 698058 193306 698294
rect 193542 698058 228986 698294
rect 229222 698058 229306 698294
rect 229542 698058 264986 698294
rect 265222 698058 265306 698294
rect 265542 698058 300986 698294
rect 301222 698058 301306 698294
rect 301542 698058 336986 698294
rect 337222 698058 337306 698294
rect 337542 698058 372986 698294
rect 373222 698058 373306 698294
rect 373542 698058 408986 698294
rect 409222 698058 409306 698294
rect 409542 698058 444986 698294
rect 445222 698058 445306 698294
rect 445542 698058 480986 698294
rect 481222 698058 481306 698294
rect 481542 698058 516986 698294
rect 517222 698058 517306 698294
rect 517542 698058 552986 698294
rect 553222 698058 553306 698294
rect 553542 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 9266 694894
rect 9502 694658 9586 694894
rect 9822 694658 45266 694894
rect 45502 694658 45586 694894
rect 45822 694658 81266 694894
rect 81502 694658 81586 694894
rect 81822 694658 117266 694894
rect 117502 694658 117586 694894
rect 117822 694658 153266 694894
rect 153502 694658 153586 694894
rect 153822 694658 189266 694894
rect 189502 694658 189586 694894
rect 189822 694658 225266 694894
rect 225502 694658 225586 694894
rect 225822 694658 261266 694894
rect 261502 694658 261586 694894
rect 261822 694658 297266 694894
rect 297502 694658 297586 694894
rect 297822 694658 333266 694894
rect 333502 694658 333586 694894
rect 333822 694658 369266 694894
rect 369502 694658 369586 694894
rect 369822 694658 405266 694894
rect 405502 694658 405586 694894
rect 405822 694658 441266 694894
rect 441502 694658 441586 694894
rect 441822 694658 477266 694894
rect 477502 694658 477586 694894
rect 477822 694658 513266 694894
rect 513502 694658 513586 694894
rect 513822 694658 549266 694894
rect 549502 694658 549586 694894
rect 549822 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 9266 694574
rect 9502 694338 9586 694574
rect 9822 694338 45266 694574
rect 45502 694338 45586 694574
rect 45822 694338 81266 694574
rect 81502 694338 81586 694574
rect 81822 694338 117266 694574
rect 117502 694338 117586 694574
rect 117822 694338 153266 694574
rect 153502 694338 153586 694574
rect 153822 694338 189266 694574
rect 189502 694338 189586 694574
rect 189822 694338 225266 694574
rect 225502 694338 225586 694574
rect 225822 694338 261266 694574
rect 261502 694338 261586 694574
rect 261822 694338 297266 694574
rect 297502 694338 297586 694574
rect 297822 694338 333266 694574
rect 333502 694338 333586 694574
rect 333822 694338 369266 694574
rect 369502 694338 369586 694574
rect 369822 694338 405266 694574
rect 405502 694338 405586 694574
rect 405822 694338 441266 694574
rect 441502 694338 441586 694574
rect 441822 694338 477266 694574
rect 477502 694338 477586 694574
rect 477822 694338 513266 694574
rect 513502 694338 513586 694574
rect 513822 694338 549266 694574
rect 549502 694338 549586 694574
rect 549822 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 5546 691174
rect 5782 690938 5866 691174
rect 6102 690938 41546 691174
rect 41782 690938 41866 691174
rect 42102 690938 77546 691174
rect 77782 690938 77866 691174
rect 78102 690938 113546 691174
rect 113782 690938 113866 691174
rect 114102 690938 149546 691174
rect 149782 690938 149866 691174
rect 150102 690938 185546 691174
rect 185782 690938 185866 691174
rect 186102 690938 221546 691174
rect 221782 690938 221866 691174
rect 222102 690938 257546 691174
rect 257782 690938 257866 691174
rect 258102 690938 293546 691174
rect 293782 690938 293866 691174
rect 294102 690938 329546 691174
rect 329782 690938 329866 691174
rect 330102 690938 365546 691174
rect 365782 690938 365866 691174
rect 366102 690938 401546 691174
rect 401782 690938 401866 691174
rect 402102 690938 437546 691174
rect 437782 690938 437866 691174
rect 438102 690938 473546 691174
rect 473782 690938 473866 691174
rect 474102 690938 509546 691174
rect 509782 690938 509866 691174
rect 510102 690938 545546 691174
rect 545782 690938 545866 691174
rect 546102 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 5546 690854
rect 5782 690618 5866 690854
rect 6102 690618 41546 690854
rect 41782 690618 41866 690854
rect 42102 690618 77546 690854
rect 77782 690618 77866 690854
rect 78102 690618 113546 690854
rect 113782 690618 113866 690854
rect 114102 690618 149546 690854
rect 149782 690618 149866 690854
rect 150102 690618 185546 690854
rect 185782 690618 185866 690854
rect 186102 690618 221546 690854
rect 221782 690618 221866 690854
rect 222102 690618 257546 690854
rect 257782 690618 257866 690854
rect 258102 690618 293546 690854
rect 293782 690618 293866 690854
rect 294102 690618 329546 690854
rect 329782 690618 329866 690854
rect 330102 690618 365546 690854
rect 365782 690618 365866 690854
rect 366102 690618 401546 690854
rect 401782 690618 401866 690854
rect 402102 690618 437546 690854
rect 437782 690618 437866 690854
rect 438102 690618 473546 690854
rect 473782 690618 473866 690854
rect 474102 690618 509546 690854
rect 509782 690618 509866 690854
rect 510102 690618 545546 690854
rect 545782 690618 545866 690854
rect 546102 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 1826 687454
rect 2062 687218 2146 687454
rect 2382 687218 37826 687454
rect 38062 687218 38146 687454
rect 38382 687218 73826 687454
rect 74062 687218 74146 687454
rect 74382 687218 109826 687454
rect 110062 687218 110146 687454
rect 110382 687218 145826 687454
rect 146062 687218 146146 687454
rect 146382 687218 181826 687454
rect 182062 687218 182146 687454
rect 182382 687218 217826 687454
rect 218062 687218 218146 687454
rect 218382 687218 253826 687454
rect 254062 687218 254146 687454
rect 254382 687218 289826 687454
rect 290062 687218 290146 687454
rect 290382 687218 325826 687454
rect 326062 687218 326146 687454
rect 326382 687218 361826 687454
rect 362062 687218 362146 687454
rect 362382 687218 397826 687454
rect 398062 687218 398146 687454
rect 398382 687218 433826 687454
rect 434062 687218 434146 687454
rect 434382 687218 469826 687454
rect 470062 687218 470146 687454
rect 470382 687218 505826 687454
rect 506062 687218 506146 687454
rect 506382 687218 541826 687454
rect 542062 687218 542146 687454
rect 542382 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 1826 687134
rect 2062 686898 2146 687134
rect 2382 686898 37826 687134
rect 38062 686898 38146 687134
rect 38382 686898 73826 687134
rect 74062 686898 74146 687134
rect 74382 686898 109826 687134
rect 110062 686898 110146 687134
rect 110382 686898 145826 687134
rect 146062 686898 146146 687134
rect 146382 686898 181826 687134
rect 182062 686898 182146 687134
rect 182382 686898 217826 687134
rect 218062 686898 218146 687134
rect 218382 686898 253826 687134
rect 254062 686898 254146 687134
rect 254382 686898 289826 687134
rect 290062 686898 290146 687134
rect 290382 686898 325826 687134
rect 326062 686898 326146 687134
rect 326382 686898 361826 687134
rect 362062 686898 362146 687134
rect 362382 686898 397826 687134
rect 398062 686898 398146 687134
rect 398382 686898 433826 687134
rect 434062 686898 434146 687134
rect 434382 686898 469826 687134
rect 470062 686898 470146 687134
rect 470382 686898 505826 687134
rect 506062 686898 506146 687134
rect 506382 686898 541826 687134
rect 542062 686898 542146 687134
rect 542382 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 30986 680614
rect 31222 680378 31306 680614
rect 31542 680378 66986 680614
rect 67222 680378 67306 680614
rect 67542 680378 102986 680614
rect 103222 680378 103306 680614
rect 103542 680378 138986 680614
rect 139222 680378 139306 680614
rect 139542 680378 174986 680614
rect 175222 680378 175306 680614
rect 175542 680378 210986 680614
rect 211222 680378 211306 680614
rect 211542 680378 246986 680614
rect 247222 680378 247306 680614
rect 247542 680378 282986 680614
rect 283222 680378 283306 680614
rect 283542 680378 318986 680614
rect 319222 680378 319306 680614
rect 319542 680378 354986 680614
rect 355222 680378 355306 680614
rect 355542 680378 390986 680614
rect 391222 680378 391306 680614
rect 391542 680378 426986 680614
rect 427222 680378 427306 680614
rect 427542 680378 462986 680614
rect 463222 680378 463306 680614
rect 463542 680378 498986 680614
rect 499222 680378 499306 680614
rect 499542 680378 534986 680614
rect 535222 680378 535306 680614
rect 535542 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 30986 680294
rect 31222 680058 31306 680294
rect 31542 680058 66986 680294
rect 67222 680058 67306 680294
rect 67542 680058 102986 680294
rect 103222 680058 103306 680294
rect 103542 680058 138986 680294
rect 139222 680058 139306 680294
rect 139542 680058 174986 680294
rect 175222 680058 175306 680294
rect 175542 680058 210986 680294
rect 211222 680058 211306 680294
rect 211542 680058 246986 680294
rect 247222 680058 247306 680294
rect 247542 680058 282986 680294
rect 283222 680058 283306 680294
rect 283542 680058 318986 680294
rect 319222 680058 319306 680294
rect 319542 680058 354986 680294
rect 355222 680058 355306 680294
rect 355542 680058 390986 680294
rect 391222 680058 391306 680294
rect 391542 680058 426986 680294
rect 427222 680058 427306 680294
rect 427542 680058 462986 680294
rect 463222 680058 463306 680294
rect 463542 680058 498986 680294
rect 499222 680058 499306 680294
rect 499542 680058 534986 680294
rect 535222 680058 535306 680294
rect 535542 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 27266 676894
rect 27502 676658 27586 676894
rect 27822 676658 63266 676894
rect 63502 676658 63586 676894
rect 63822 676658 99266 676894
rect 99502 676658 99586 676894
rect 99822 676658 135266 676894
rect 135502 676658 135586 676894
rect 135822 676658 171266 676894
rect 171502 676658 171586 676894
rect 171822 676658 207266 676894
rect 207502 676658 207586 676894
rect 207822 676658 243266 676894
rect 243502 676658 243586 676894
rect 243822 676658 279266 676894
rect 279502 676658 279586 676894
rect 279822 676658 315266 676894
rect 315502 676658 315586 676894
rect 315822 676658 351266 676894
rect 351502 676658 351586 676894
rect 351822 676658 387266 676894
rect 387502 676658 387586 676894
rect 387822 676658 423266 676894
rect 423502 676658 423586 676894
rect 423822 676658 459266 676894
rect 459502 676658 459586 676894
rect 459822 676658 495266 676894
rect 495502 676658 495586 676894
rect 495822 676658 531266 676894
rect 531502 676658 531586 676894
rect 531822 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 27266 676574
rect 27502 676338 27586 676574
rect 27822 676338 63266 676574
rect 63502 676338 63586 676574
rect 63822 676338 99266 676574
rect 99502 676338 99586 676574
rect 99822 676338 135266 676574
rect 135502 676338 135586 676574
rect 135822 676338 171266 676574
rect 171502 676338 171586 676574
rect 171822 676338 207266 676574
rect 207502 676338 207586 676574
rect 207822 676338 243266 676574
rect 243502 676338 243586 676574
rect 243822 676338 279266 676574
rect 279502 676338 279586 676574
rect 279822 676338 315266 676574
rect 315502 676338 315586 676574
rect 315822 676338 351266 676574
rect 351502 676338 351586 676574
rect 351822 676338 387266 676574
rect 387502 676338 387586 676574
rect 387822 676338 423266 676574
rect 423502 676338 423586 676574
rect 423822 676338 459266 676574
rect 459502 676338 459586 676574
rect 459822 676338 495266 676574
rect 495502 676338 495586 676574
rect 495822 676338 531266 676574
rect 531502 676338 531586 676574
rect 531822 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 23546 673174
rect 23782 672938 23866 673174
rect 24102 672938 59546 673174
rect 59782 672938 59866 673174
rect 60102 672938 95546 673174
rect 95782 672938 95866 673174
rect 96102 672938 131546 673174
rect 131782 672938 131866 673174
rect 132102 672938 167546 673174
rect 167782 672938 167866 673174
rect 168102 672938 203546 673174
rect 203782 672938 203866 673174
rect 204102 672938 239546 673174
rect 239782 672938 239866 673174
rect 240102 672938 275546 673174
rect 275782 672938 275866 673174
rect 276102 672938 311546 673174
rect 311782 672938 311866 673174
rect 312102 672938 347546 673174
rect 347782 672938 347866 673174
rect 348102 672938 383546 673174
rect 383782 672938 383866 673174
rect 384102 672938 419546 673174
rect 419782 672938 419866 673174
rect 420102 672938 455546 673174
rect 455782 672938 455866 673174
rect 456102 672938 491546 673174
rect 491782 672938 491866 673174
rect 492102 672938 527546 673174
rect 527782 672938 527866 673174
rect 528102 672938 563546 673174
rect 563782 672938 563866 673174
rect 564102 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 23546 672854
rect 23782 672618 23866 672854
rect 24102 672618 59546 672854
rect 59782 672618 59866 672854
rect 60102 672618 95546 672854
rect 95782 672618 95866 672854
rect 96102 672618 131546 672854
rect 131782 672618 131866 672854
rect 132102 672618 167546 672854
rect 167782 672618 167866 672854
rect 168102 672618 203546 672854
rect 203782 672618 203866 672854
rect 204102 672618 239546 672854
rect 239782 672618 239866 672854
rect 240102 672618 275546 672854
rect 275782 672618 275866 672854
rect 276102 672618 311546 672854
rect 311782 672618 311866 672854
rect 312102 672618 347546 672854
rect 347782 672618 347866 672854
rect 348102 672618 383546 672854
rect 383782 672618 383866 672854
rect 384102 672618 419546 672854
rect 419782 672618 419866 672854
rect 420102 672618 455546 672854
rect 455782 672618 455866 672854
rect 456102 672618 491546 672854
rect 491782 672618 491866 672854
rect 492102 672618 527546 672854
rect 527782 672618 527866 672854
rect 528102 672618 563546 672854
rect 563782 672618 563866 672854
rect 564102 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 19826 669454
rect 20062 669218 20146 669454
rect 20382 669218 55826 669454
rect 56062 669218 56146 669454
rect 56382 669218 91826 669454
rect 92062 669218 92146 669454
rect 92382 669218 127826 669454
rect 128062 669218 128146 669454
rect 128382 669218 163826 669454
rect 164062 669218 164146 669454
rect 164382 669218 199826 669454
rect 200062 669218 200146 669454
rect 200382 669218 235826 669454
rect 236062 669218 236146 669454
rect 236382 669218 271826 669454
rect 272062 669218 272146 669454
rect 272382 669218 307826 669454
rect 308062 669218 308146 669454
rect 308382 669218 343826 669454
rect 344062 669218 344146 669454
rect 344382 669218 379826 669454
rect 380062 669218 380146 669454
rect 380382 669218 415826 669454
rect 416062 669218 416146 669454
rect 416382 669218 451826 669454
rect 452062 669218 452146 669454
rect 452382 669218 487826 669454
rect 488062 669218 488146 669454
rect 488382 669218 523826 669454
rect 524062 669218 524146 669454
rect 524382 669218 559826 669454
rect 560062 669218 560146 669454
rect 560382 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 19826 669134
rect 20062 668898 20146 669134
rect 20382 668898 55826 669134
rect 56062 668898 56146 669134
rect 56382 668898 91826 669134
rect 92062 668898 92146 669134
rect 92382 668898 127826 669134
rect 128062 668898 128146 669134
rect 128382 668898 163826 669134
rect 164062 668898 164146 669134
rect 164382 668898 199826 669134
rect 200062 668898 200146 669134
rect 200382 668898 235826 669134
rect 236062 668898 236146 669134
rect 236382 668898 271826 669134
rect 272062 668898 272146 669134
rect 272382 668898 307826 669134
rect 308062 668898 308146 669134
rect 308382 668898 343826 669134
rect 344062 668898 344146 669134
rect 344382 668898 379826 669134
rect 380062 668898 380146 669134
rect 380382 668898 415826 669134
rect 416062 668898 416146 669134
rect 416382 668898 451826 669134
rect 452062 668898 452146 669134
rect 452382 668898 487826 669134
rect 488062 668898 488146 669134
rect 488382 668898 523826 669134
rect 524062 668898 524146 669134
rect 524382 668898 559826 669134
rect 560062 668898 560146 669134
rect 560382 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 12986 662614
rect 13222 662378 13306 662614
rect 13542 662378 48986 662614
rect 49222 662378 49306 662614
rect 49542 662378 84986 662614
rect 85222 662378 85306 662614
rect 85542 662378 120986 662614
rect 121222 662378 121306 662614
rect 121542 662378 156986 662614
rect 157222 662378 157306 662614
rect 157542 662378 192986 662614
rect 193222 662378 193306 662614
rect 193542 662378 228986 662614
rect 229222 662378 229306 662614
rect 229542 662378 264986 662614
rect 265222 662378 265306 662614
rect 265542 662378 300986 662614
rect 301222 662378 301306 662614
rect 301542 662378 336986 662614
rect 337222 662378 337306 662614
rect 337542 662378 372986 662614
rect 373222 662378 373306 662614
rect 373542 662378 408986 662614
rect 409222 662378 409306 662614
rect 409542 662378 444986 662614
rect 445222 662378 445306 662614
rect 445542 662378 480986 662614
rect 481222 662378 481306 662614
rect 481542 662378 516986 662614
rect 517222 662378 517306 662614
rect 517542 662378 552986 662614
rect 553222 662378 553306 662614
rect 553542 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 12986 662294
rect 13222 662058 13306 662294
rect 13542 662058 48986 662294
rect 49222 662058 49306 662294
rect 49542 662058 84986 662294
rect 85222 662058 85306 662294
rect 85542 662058 120986 662294
rect 121222 662058 121306 662294
rect 121542 662058 156986 662294
rect 157222 662058 157306 662294
rect 157542 662058 192986 662294
rect 193222 662058 193306 662294
rect 193542 662058 228986 662294
rect 229222 662058 229306 662294
rect 229542 662058 264986 662294
rect 265222 662058 265306 662294
rect 265542 662058 300986 662294
rect 301222 662058 301306 662294
rect 301542 662058 336986 662294
rect 337222 662058 337306 662294
rect 337542 662058 372986 662294
rect 373222 662058 373306 662294
rect 373542 662058 408986 662294
rect 409222 662058 409306 662294
rect 409542 662058 444986 662294
rect 445222 662058 445306 662294
rect 445542 662058 480986 662294
rect 481222 662058 481306 662294
rect 481542 662058 516986 662294
rect 517222 662058 517306 662294
rect 517542 662058 552986 662294
rect 553222 662058 553306 662294
rect 553542 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 9266 658894
rect 9502 658658 9586 658894
rect 9822 658658 45266 658894
rect 45502 658658 45586 658894
rect 45822 658658 81266 658894
rect 81502 658658 81586 658894
rect 81822 658658 117266 658894
rect 117502 658658 117586 658894
rect 117822 658658 153266 658894
rect 153502 658658 153586 658894
rect 153822 658658 189266 658894
rect 189502 658658 189586 658894
rect 189822 658658 225266 658894
rect 225502 658658 225586 658894
rect 225822 658658 261266 658894
rect 261502 658658 261586 658894
rect 261822 658658 297266 658894
rect 297502 658658 297586 658894
rect 297822 658658 333266 658894
rect 333502 658658 333586 658894
rect 333822 658658 369266 658894
rect 369502 658658 369586 658894
rect 369822 658658 405266 658894
rect 405502 658658 405586 658894
rect 405822 658658 441266 658894
rect 441502 658658 441586 658894
rect 441822 658658 477266 658894
rect 477502 658658 477586 658894
rect 477822 658658 513266 658894
rect 513502 658658 513586 658894
rect 513822 658658 549266 658894
rect 549502 658658 549586 658894
rect 549822 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 9266 658574
rect 9502 658338 9586 658574
rect 9822 658338 45266 658574
rect 45502 658338 45586 658574
rect 45822 658338 81266 658574
rect 81502 658338 81586 658574
rect 81822 658338 117266 658574
rect 117502 658338 117586 658574
rect 117822 658338 153266 658574
rect 153502 658338 153586 658574
rect 153822 658338 189266 658574
rect 189502 658338 189586 658574
rect 189822 658338 225266 658574
rect 225502 658338 225586 658574
rect 225822 658338 261266 658574
rect 261502 658338 261586 658574
rect 261822 658338 297266 658574
rect 297502 658338 297586 658574
rect 297822 658338 333266 658574
rect 333502 658338 333586 658574
rect 333822 658338 369266 658574
rect 369502 658338 369586 658574
rect 369822 658338 405266 658574
rect 405502 658338 405586 658574
rect 405822 658338 441266 658574
rect 441502 658338 441586 658574
rect 441822 658338 477266 658574
rect 477502 658338 477586 658574
rect 477822 658338 513266 658574
rect 513502 658338 513586 658574
rect 513822 658338 549266 658574
rect 549502 658338 549586 658574
rect 549822 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 5546 655174
rect 5782 654938 5866 655174
rect 6102 654938 41546 655174
rect 41782 654938 41866 655174
rect 42102 654938 77546 655174
rect 77782 654938 77866 655174
rect 78102 654938 113546 655174
rect 113782 654938 113866 655174
rect 114102 654938 149546 655174
rect 149782 654938 149866 655174
rect 150102 654938 185546 655174
rect 185782 654938 185866 655174
rect 186102 654938 221546 655174
rect 221782 654938 221866 655174
rect 222102 654938 257546 655174
rect 257782 654938 257866 655174
rect 258102 654938 293546 655174
rect 293782 654938 293866 655174
rect 294102 654938 329546 655174
rect 329782 654938 329866 655174
rect 330102 654938 365546 655174
rect 365782 654938 365866 655174
rect 366102 654938 401546 655174
rect 401782 654938 401866 655174
rect 402102 654938 437546 655174
rect 437782 654938 437866 655174
rect 438102 654938 473546 655174
rect 473782 654938 473866 655174
rect 474102 654938 509546 655174
rect 509782 654938 509866 655174
rect 510102 654938 545546 655174
rect 545782 654938 545866 655174
rect 546102 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 5546 654854
rect 5782 654618 5866 654854
rect 6102 654618 41546 654854
rect 41782 654618 41866 654854
rect 42102 654618 77546 654854
rect 77782 654618 77866 654854
rect 78102 654618 113546 654854
rect 113782 654618 113866 654854
rect 114102 654618 149546 654854
rect 149782 654618 149866 654854
rect 150102 654618 185546 654854
rect 185782 654618 185866 654854
rect 186102 654618 221546 654854
rect 221782 654618 221866 654854
rect 222102 654618 257546 654854
rect 257782 654618 257866 654854
rect 258102 654618 293546 654854
rect 293782 654618 293866 654854
rect 294102 654618 329546 654854
rect 329782 654618 329866 654854
rect 330102 654618 365546 654854
rect 365782 654618 365866 654854
rect 366102 654618 401546 654854
rect 401782 654618 401866 654854
rect 402102 654618 437546 654854
rect 437782 654618 437866 654854
rect 438102 654618 473546 654854
rect 473782 654618 473866 654854
rect 474102 654618 509546 654854
rect 509782 654618 509866 654854
rect 510102 654618 545546 654854
rect 545782 654618 545866 654854
rect 546102 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 1826 651454
rect 2062 651218 2146 651454
rect 2382 651218 37826 651454
rect 38062 651218 38146 651454
rect 38382 651218 73826 651454
rect 74062 651218 74146 651454
rect 74382 651218 109826 651454
rect 110062 651218 110146 651454
rect 110382 651218 145826 651454
rect 146062 651218 146146 651454
rect 146382 651218 181826 651454
rect 182062 651218 182146 651454
rect 182382 651218 217826 651454
rect 218062 651218 218146 651454
rect 218382 651218 253826 651454
rect 254062 651218 254146 651454
rect 254382 651218 289826 651454
rect 290062 651218 290146 651454
rect 290382 651218 325826 651454
rect 326062 651218 326146 651454
rect 326382 651218 361826 651454
rect 362062 651218 362146 651454
rect 362382 651218 397826 651454
rect 398062 651218 398146 651454
rect 398382 651218 433826 651454
rect 434062 651218 434146 651454
rect 434382 651218 469826 651454
rect 470062 651218 470146 651454
rect 470382 651218 505826 651454
rect 506062 651218 506146 651454
rect 506382 651218 541826 651454
rect 542062 651218 542146 651454
rect 542382 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 1826 651134
rect 2062 650898 2146 651134
rect 2382 650898 37826 651134
rect 38062 650898 38146 651134
rect 38382 650898 73826 651134
rect 74062 650898 74146 651134
rect 74382 650898 109826 651134
rect 110062 650898 110146 651134
rect 110382 650898 145826 651134
rect 146062 650898 146146 651134
rect 146382 650898 181826 651134
rect 182062 650898 182146 651134
rect 182382 650898 217826 651134
rect 218062 650898 218146 651134
rect 218382 650898 253826 651134
rect 254062 650898 254146 651134
rect 254382 650898 289826 651134
rect 290062 650898 290146 651134
rect 290382 650898 325826 651134
rect 326062 650898 326146 651134
rect 326382 650898 361826 651134
rect 362062 650898 362146 651134
rect 362382 650898 397826 651134
rect 398062 650898 398146 651134
rect 398382 650898 433826 651134
rect 434062 650898 434146 651134
rect 434382 650898 469826 651134
rect 470062 650898 470146 651134
rect 470382 650898 505826 651134
rect 506062 650898 506146 651134
rect 506382 650898 541826 651134
rect 542062 650898 542146 651134
rect 542382 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 30986 644614
rect 31222 644378 31306 644614
rect 31542 644378 66986 644614
rect 67222 644378 67306 644614
rect 67542 644378 102986 644614
rect 103222 644378 103306 644614
rect 103542 644378 138986 644614
rect 139222 644378 139306 644614
rect 139542 644378 174986 644614
rect 175222 644378 175306 644614
rect 175542 644378 210986 644614
rect 211222 644378 211306 644614
rect 211542 644378 246986 644614
rect 247222 644378 247306 644614
rect 247542 644378 282986 644614
rect 283222 644378 283306 644614
rect 283542 644378 318986 644614
rect 319222 644378 319306 644614
rect 319542 644378 354986 644614
rect 355222 644378 355306 644614
rect 355542 644378 390986 644614
rect 391222 644378 391306 644614
rect 391542 644378 426986 644614
rect 427222 644378 427306 644614
rect 427542 644378 462986 644614
rect 463222 644378 463306 644614
rect 463542 644378 498986 644614
rect 499222 644378 499306 644614
rect 499542 644378 534986 644614
rect 535222 644378 535306 644614
rect 535542 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 30986 644294
rect 31222 644058 31306 644294
rect 31542 644058 66986 644294
rect 67222 644058 67306 644294
rect 67542 644058 102986 644294
rect 103222 644058 103306 644294
rect 103542 644058 138986 644294
rect 139222 644058 139306 644294
rect 139542 644058 174986 644294
rect 175222 644058 175306 644294
rect 175542 644058 210986 644294
rect 211222 644058 211306 644294
rect 211542 644058 246986 644294
rect 247222 644058 247306 644294
rect 247542 644058 282986 644294
rect 283222 644058 283306 644294
rect 283542 644058 318986 644294
rect 319222 644058 319306 644294
rect 319542 644058 354986 644294
rect 355222 644058 355306 644294
rect 355542 644058 390986 644294
rect 391222 644058 391306 644294
rect 391542 644058 426986 644294
rect 427222 644058 427306 644294
rect 427542 644058 462986 644294
rect 463222 644058 463306 644294
rect 463542 644058 498986 644294
rect 499222 644058 499306 644294
rect 499542 644058 534986 644294
rect 535222 644058 535306 644294
rect 535542 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 27266 640894
rect 27502 640658 27586 640894
rect 27822 640658 63266 640894
rect 63502 640658 63586 640894
rect 63822 640658 99266 640894
rect 99502 640658 99586 640894
rect 99822 640658 135266 640894
rect 135502 640658 135586 640894
rect 135822 640658 171266 640894
rect 171502 640658 171586 640894
rect 171822 640658 207266 640894
rect 207502 640658 207586 640894
rect 207822 640658 243266 640894
rect 243502 640658 243586 640894
rect 243822 640658 279266 640894
rect 279502 640658 279586 640894
rect 279822 640658 315266 640894
rect 315502 640658 315586 640894
rect 315822 640658 351266 640894
rect 351502 640658 351586 640894
rect 351822 640658 387266 640894
rect 387502 640658 387586 640894
rect 387822 640658 423266 640894
rect 423502 640658 423586 640894
rect 423822 640658 459266 640894
rect 459502 640658 459586 640894
rect 459822 640658 495266 640894
rect 495502 640658 495586 640894
rect 495822 640658 531266 640894
rect 531502 640658 531586 640894
rect 531822 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 27266 640574
rect 27502 640338 27586 640574
rect 27822 640338 63266 640574
rect 63502 640338 63586 640574
rect 63822 640338 99266 640574
rect 99502 640338 99586 640574
rect 99822 640338 135266 640574
rect 135502 640338 135586 640574
rect 135822 640338 171266 640574
rect 171502 640338 171586 640574
rect 171822 640338 207266 640574
rect 207502 640338 207586 640574
rect 207822 640338 243266 640574
rect 243502 640338 243586 640574
rect 243822 640338 279266 640574
rect 279502 640338 279586 640574
rect 279822 640338 315266 640574
rect 315502 640338 315586 640574
rect 315822 640338 351266 640574
rect 351502 640338 351586 640574
rect 351822 640338 387266 640574
rect 387502 640338 387586 640574
rect 387822 640338 423266 640574
rect 423502 640338 423586 640574
rect 423822 640338 459266 640574
rect 459502 640338 459586 640574
rect 459822 640338 495266 640574
rect 495502 640338 495586 640574
rect 495822 640338 531266 640574
rect 531502 640338 531586 640574
rect 531822 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 23546 637174
rect 23782 636938 23866 637174
rect 24102 636938 59546 637174
rect 59782 636938 59866 637174
rect 60102 636938 95546 637174
rect 95782 636938 95866 637174
rect 96102 636938 131546 637174
rect 131782 636938 131866 637174
rect 132102 636938 167546 637174
rect 167782 636938 167866 637174
rect 168102 636938 203546 637174
rect 203782 636938 203866 637174
rect 204102 636938 239546 637174
rect 239782 636938 239866 637174
rect 240102 636938 275546 637174
rect 275782 636938 275866 637174
rect 276102 636938 311546 637174
rect 311782 636938 311866 637174
rect 312102 636938 347546 637174
rect 347782 636938 347866 637174
rect 348102 636938 383546 637174
rect 383782 636938 383866 637174
rect 384102 636938 419546 637174
rect 419782 636938 419866 637174
rect 420102 636938 455546 637174
rect 455782 636938 455866 637174
rect 456102 636938 491546 637174
rect 491782 636938 491866 637174
rect 492102 636938 527546 637174
rect 527782 636938 527866 637174
rect 528102 636938 563546 637174
rect 563782 636938 563866 637174
rect 564102 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 23546 636854
rect 23782 636618 23866 636854
rect 24102 636618 59546 636854
rect 59782 636618 59866 636854
rect 60102 636618 95546 636854
rect 95782 636618 95866 636854
rect 96102 636618 131546 636854
rect 131782 636618 131866 636854
rect 132102 636618 167546 636854
rect 167782 636618 167866 636854
rect 168102 636618 203546 636854
rect 203782 636618 203866 636854
rect 204102 636618 239546 636854
rect 239782 636618 239866 636854
rect 240102 636618 275546 636854
rect 275782 636618 275866 636854
rect 276102 636618 311546 636854
rect 311782 636618 311866 636854
rect 312102 636618 347546 636854
rect 347782 636618 347866 636854
rect 348102 636618 383546 636854
rect 383782 636618 383866 636854
rect 384102 636618 419546 636854
rect 419782 636618 419866 636854
rect 420102 636618 455546 636854
rect 455782 636618 455866 636854
rect 456102 636618 491546 636854
rect 491782 636618 491866 636854
rect 492102 636618 527546 636854
rect 527782 636618 527866 636854
rect 528102 636618 563546 636854
rect 563782 636618 563866 636854
rect 564102 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 19826 633454
rect 20062 633218 20146 633454
rect 20382 633218 55826 633454
rect 56062 633218 56146 633454
rect 56382 633218 91826 633454
rect 92062 633218 92146 633454
rect 92382 633218 127826 633454
rect 128062 633218 128146 633454
rect 128382 633218 163826 633454
rect 164062 633218 164146 633454
rect 164382 633218 199826 633454
rect 200062 633218 200146 633454
rect 200382 633218 235826 633454
rect 236062 633218 236146 633454
rect 236382 633218 271826 633454
rect 272062 633218 272146 633454
rect 272382 633218 307826 633454
rect 308062 633218 308146 633454
rect 308382 633218 343826 633454
rect 344062 633218 344146 633454
rect 344382 633218 379826 633454
rect 380062 633218 380146 633454
rect 380382 633218 415826 633454
rect 416062 633218 416146 633454
rect 416382 633218 451826 633454
rect 452062 633218 452146 633454
rect 452382 633218 487826 633454
rect 488062 633218 488146 633454
rect 488382 633218 523826 633454
rect 524062 633218 524146 633454
rect 524382 633218 559826 633454
rect 560062 633218 560146 633454
rect 560382 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 19826 633134
rect 20062 632898 20146 633134
rect 20382 632898 55826 633134
rect 56062 632898 56146 633134
rect 56382 632898 91826 633134
rect 92062 632898 92146 633134
rect 92382 632898 127826 633134
rect 128062 632898 128146 633134
rect 128382 632898 163826 633134
rect 164062 632898 164146 633134
rect 164382 632898 199826 633134
rect 200062 632898 200146 633134
rect 200382 632898 235826 633134
rect 236062 632898 236146 633134
rect 236382 632898 271826 633134
rect 272062 632898 272146 633134
rect 272382 632898 307826 633134
rect 308062 632898 308146 633134
rect 308382 632898 343826 633134
rect 344062 632898 344146 633134
rect 344382 632898 379826 633134
rect 380062 632898 380146 633134
rect 380382 632898 415826 633134
rect 416062 632898 416146 633134
rect 416382 632898 451826 633134
rect 452062 632898 452146 633134
rect 452382 632898 487826 633134
rect 488062 632898 488146 633134
rect 488382 632898 523826 633134
rect 524062 632898 524146 633134
rect 524382 632898 559826 633134
rect 560062 632898 560146 633134
rect 560382 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 12986 626614
rect 13222 626378 13306 626614
rect 13542 626378 48986 626614
rect 49222 626378 49306 626614
rect 49542 626378 84986 626614
rect 85222 626378 85306 626614
rect 85542 626378 120986 626614
rect 121222 626378 121306 626614
rect 121542 626378 156986 626614
rect 157222 626378 157306 626614
rect 157542 626378 192986 626614
rect 193222 626378 193306 626614
rect 193542 626378 228986 626614
rect 229222 626378 229306 626614
rect 229542 626378 264986 626614
rect 265222 626378 265306 626614
rect 265542 626378 300986 626614
rect 301222 626378 301306 626614
rect 301542 626378 336986 626614
rect 337222 626378 337306 626614
rect 337542 626378 372986 626614
rect 373222 626378 373306 626614
rect 373542 626378 408986 626614
rect 409222 626378 409306 626614
rect 409542 626378 444986 626614
rect 445222 626378 445306 626614
rect 445542 626378 480986 626614
rect 481222 626378 481306 626614
rect 481542 626378 516986 626614
rect 517222 626378 517306 626614
rect 517542 626378 552986 626614
rect 553222 626378 553306 626614
rect 553542 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 12986 626294
rect 13222 626058 13306 626294
rect 13542 626058 48986 626294
rect 49222 626058 49306 626294
rect 49542 626058 84986 626294
rect 85222 626058 85306 626294
rect 85542 626058 120986 626294
rect 121222 626058 121306 626294
rect 121542 626058 156986 626294
rect 157222 626058 157306 626294
rect 157542 626058 192986 626294
rect 193222 626058 193306 626294
rect 193542 626058 228986 626294
rect 229222 626058 229306 626294
rect 229542 626058 264986 626294
rect 265222 626058 265306 626294
rect 265542 626058 300986 626294
rect 301222 626058 301306 626294
rect 301542 626058 336986 626294
rect 337222 626058 337306 626294
rect 337542 626058 372986 626294
rect 373222 626058 373306 626294
rect 373542 626058 408986 626294
rect 409222 626058 409306 626294
rect 409542 626058 444986 626294
rect 445222 626058 445306 626294
rect 445542 626058 480986 626294
rect 481222 626058 481306 626294
rect 481542 626058 516986 626294
rect 517222 626058 517306 626294
rect 517542 626058 552986 626294
rect 553222 626058 553306 626294
rect 553542 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 9266 622894
rect 9502 622658 9586 622894
rect 9822 622658 45266 622894
rect 45502 622658 45586 622894
rect 45822 622658 81266 622894
rect 81502 622658 81586 622894
rect 81822 622658 117266 622894
rect 117502 622658 117586 622894
rect 117822 622658 153266 622894
rect 153502 622658 153586 622894
rect 153822 622658 189266 622894
rect 189502 622658 189586 622894
rect 189822 622658 225266 622894
rect 225502 622658 225586 622894
rect 225822 622658 261266 622894
rect 261502 622658 261586 622894
rect 261822 622658 297266 622894
rect 297502 622658 297586 622894
rect 297822 622658 333266 622894
rect 333502 622658 333586 622894
rect 333822 622658 369266 622894
rect 369502 622658 369586 622894
rect 369822 622658 405266 622894
rect 405502 622658 405586 622894
rect 405822 622658 441266 622894
rect 441502 622658 441586 622894
rect 441822 622658 477266 622894
rect 477502 622658 477586 622894
rect 477822 622658 513266 622894
rect 513502 622658 513586 622894
rect 513822 622658 549266 622894
rect 549502 622658 549586 622894
rect 549822 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 9266 622574
rect 9502 622338 9586 622574
rect 9822 622338 45266 622574
rect 45502 622338 45586 622574
rect 45822 622338 81266 622574
rect 81502 622338 81586 622574
rect 81822 622338 117266 622574
rect 117502 622338 117586 622574
rect 117822 622338 153266 622574
rect 153502 622338 153586 622574
rect 153822 622338 189266 622574
rect 189502 622338 189586 622574
rect 189822 622338 225266 622574
rect 225502 622338 225586 622574
rect 225822 622338 261266 622574
rect 261502 622338 261586 622574
rect 261822 622338 297266 622574
rect 297502 622338 297586 622574
rect 297822 622338 333266 622574
rect 333502 622338 333586 622574
rect 333822 622338 369266 622574
rect 369502 622338 369586 622574
rect 369822 622338 405266 622574
rect 405502 622338 405586 622574
rect 405822 622338 441266 622574
rect 441502 622338 441586 622574
rect 441822 622338 477266 622574
rect 477502 622338 477586 622574
rect 477822 622338 513266 622574
rect 513502 622338 513586 622574
rect 513822 622338 549266 622574
rect 549502 622338 549586 622574
rect 549822 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 5546 619174
rect 5782 618938 5866 619174
rect 6102 618938 41546 619174
rect 41782 618938 41866 619174
rect 42102 618938 77546 619174
rect 77782 618938 77866 619174
rect 78102 618938 113546 619174
rect 113782 618938 113866 619174
rect 114102 618938 149546 619174
rect 149782 618938 149866 619174
rect 150102 618938 185546 619174
rect 185782 618938 185866 619174
rect 186102 618938 221546 619174
rect 221782 618938 221866 619174
rect 222102 618938 257546 619174
rect 257782 618938 257866 619174
rect 258102 618938 293546 619174
rect 293782 618938 293866 619174
rect 294102 618938 329546 619174
rect 329782 618938 329866 619174
rect 330102 618938 365546 619174
rect 365782 618938 365866 619174
rect 366102 618938 401546 619174
rect 401782 618938 401866 619174
rect 402102 618938 437546 619174
rect 437782 618938 437866 619174
rect 438102 618938 473546 619174
rect 473782 618938 473866 619174
rect 474102 618938 509546 619174
rect 509782 618938 509866 619174
rect 510102 618938 545546 619174
rect 545782 618938 545866 619174
rect 546102 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 5546 618854
rect 5782 618618 5866 618854
rect 6102 618618 41546 618854
rect 41782 618618 41866 618854
rect 42102 618618 77546 618854
rect 77782 618618 77866 618854
rect 78102 618618 113546 618854
rect 113782 618618 113866 618854
rect 114102 618618 149546 618854
rect 149782 618618 149866 618854
rect 150102 618618 185546 618854
rect 185782 618618 185866 618854
rect 186102 618618 221546 618854
rect 221782 618618 221866 618854
rect 222102 618618 257546 618854
rect 257782 618618 257866 618854
rect 258102 618618 293546 618854
rect 293782 618618 293866 618854
rect 294102 618618 329546 618854
rect 329782 618618 329866 618854
rect 330102 618618 365546 618854
rect 365782 618618 365866 618854
rect 366102 618618 401546 618854
rect 401782 618618 401866 618854
rect 402102 618618 437546 618854
rect 437782 618618 437866 618854
rect 438102 618618 473546 618854
rect 473782 618618 473866 618854
rect 474102 618618 509546 618854
rect 509782 618618 509866 618854
rect 510102 618618 545546 618854
rect 545782 618618 545866 618854
rect 546102 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 1826 615454
rect 2062 615218 2146 615454
rect 2382 615218 37826 615454
rect 38062 615218 38146 615454
rect 38382 615218 73826 615454
rect 74062 615218 74146 615454
rect 74382 615218 109826 615454
rect 110062 615218 110146 615454
rect 110382 615218 145826 615454
rect 146062 615218 146146 615454
rect 146382 615218 181826 615454
rect 182062 615218 182146 615454
rect 182382 615218 217826 615454
rect 218062 615218 218146 615454
rect 218382 615218 253826 615454
rect 254062 615218 254146 615454
rect 254382 615218 289826 615454
rect 290062 615218 290146 615454
rect 290382 615218 325826 615454
rect 326062 615218 326146 615454
rect 326382 615218 361826 615454
rect 362062 615218 362146 615454
rect 362382 615218 397826 615454
rect 398062 615218 398146 615454
rect 398382 615218 433826 615454
rect 434062 615218 434146 615454
rect 434382 615218 469826 615454
rect 470062 615218 470146 615454
rect 470382 615218 505826 615454
rect 506062 615218 506146 615454
rect 506382 615218 541826 615454
rect 542062 615218 542146 615454
rect 542382 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 1826 615134
rect 2062 614898 2146 615134
rect 2382 614898 37826 615134
rect 38062 614898 38146 615134
rect 38382 614898 73826 615134
rect 74062 614898 74146 615134
rect 74382 614898 109826 615134
rect 110062 614898 110146 615134
rect 110382 614898 145826 615134
rect 146062 614898 146146 615134
rect 146382 614898 181826 615134
rect 182062 614898 182146 615134
rect 182382 614898 217826 615134
rect 218062 614898 218146 615134
rect 218382 614898 253826 615134
rect 254062 614898 254146 615134
rect 254382 614898 289826 615134
rect 290062 614898 290146 615134
rect 290382 614898 325826 615134
rect 326062 614898 326146 615134
rect 326382 614898 361826 615134
rect 362062 614898 362146 615134
rect 362382 614898 397826 615134
rect 398062 614898 398146 615134
rect 398382 614898 433826 615134
rect 434062 614898 434146 615134
rect 434382 614898 469826 615134
rect 470062 614898 470146 615134
rect 470382 614898 505826 615134
rect 506062 614898 506146 615134
rect 506382 614898 541826 615134
rect 542062 614898 542146 615134
rect 542382 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 30986 608614
rect 31222 608378 31306 608614
rect 31542 608378 66986 608614
rect 67222 608378 67306 608614
rect 67542 608378 102986 608614
rect 103222 608378 103306 608614
rect 103542 608378 138986 608614
rect 139222 608378 139306 608614
rect 139542 608378 174986 608614
rect 175222 608378 175306 608614
rect 175542 608378 210986 608614
rect 211222 608378 211306 608614
rect 211542 608378 246986 608614
rect 247222 608378 247306 608614
rect 247542 608378 282986 608614
rect 283222 608378 283306 608614
rect 283542 608378 318986 608614
rect 319222 608378 319306 608614
rect 319542 608378 354986 608614
rect 355222 608378 355306 608614
rect 355542 608378 390986 608614
rect 391222 608378 391306 608614
rect 391542 608378 426986 608614
rect 427222 608378 427306 608614
rect 427542 608378 462986 608614
rect 463222 608378 463306 608614
rect 463542 608378 498986 608614
rect 499222 608378 499306 608614
rect 499542 608378 534986 608614
rect 535222 608378 535306 608614
rect 535542 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 30986 608294
rect 31222 608058 31306 608294
rect 31542 608058 66986 608294
rect 67222 608058 67306 608294
rect 67542 608058 102986 608294
rect 103222 608058 103306 608294
rect 103542 608058 138986 608294
rect 139222 608058 139306 608294
rect 139542 608058 174986 608294
rect 175222 608058 175306 608294
rect 175542 608058 210986 608294
rect 211222 608058 211306 608294
rect 211542 608058 246986 608294
rect 247222 608058 247306 608294
rect 247542 608058 282986 608294
rect 283222 608058 283306 608294
rect 283542 608058 318986 608294
rect 319222 608058 319306 608294
rect 319542 608058 354986 608294
rect 355222 608058 355306 608294
rect 355542 608058 390986 608294
rect 391222 608058 391306 608294
rect 391542 608058 426986 608294
rect 427222 608058 427306 608294
rect 427542 608058 462986 608294
rect 463222 608058 463306 608294
rect 463542 608058 498986 608294
rect 499222 608058 499306 608294
rect 499542 608058 534986 608294
rect 535222 608058 535306 608294
rect 535542 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 27266 604894
rect 27502 604658 27586 604894
rect 27822 604658 63266 604894
rect 63502 604658 63586 604894
rect 63822 604658 99266 604894
rect 99502 604658 99586 604894
rect 99822 604658 135266 604894
rect 135502 604658 135586 604894
rect 135822 604658 171266 604894
rect 171502 604658 171586 604894
rect 171822 604658 207266 604894
rect 207502 604658 207586 604894
rect 207822 604658 243266 604894
rect 243502 604658 243586 604894
rect 243822 604658 279266 604894
rect 279502 604658 279586 604894
rect 279822 604658 315266 604894
rect 315502 604658 315586 604894
rect 315822 604658 351266 604894
rect 351502 604658 351586 604894
rect 351822 604658 387266 604894
rect 387502 604658 387586 604894
rect 387822 604658 423266 604894
rect 423502 604658 423586 604894
rect 423822 604658 459266 604894
rect 459502 604658 459586 604894
rect 459822 604658 495266 604894
rect 495502 604658 495586 604894
rect 495822 604658 531266 604894
rect 531502 604658 531586 604894
rect 531822 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 27266 604574
rect 27502 604338 27586 604574
rect 27822 604338 63266 604574
rect 63502 604338 63586 604574
rect 63822 604338 99266 604574
rect 99502 604338 99586 604574
rect 99822 604338 135266 604574
rect 135502 604338 135586 604574
rect 135822 604338 171266 604574
rect 171502 604338 171586 604574
rect 171822 604338 207266 604574
rect 207502 604338 207586 604574
rect 207822 604338 243266 604574
rect 243502 604338 243586 604574
rect 243822 604338 279266 604574
rect 279502 604338 279586 604574
rect 279822 604338 315266 604574
rect 315502 604338 315586 604574
rect 315822 604338 351266 604574
rect 351502 604338 351586 604574
rect 351822 604338 387266 604574
rect 387502 604338 387586 604574
rect 387822 604338 423266 604574
rect 423502 604338 423586 604574
rect 423822 604338 459266 604574
rect 459502 604338 459586 604574
rect 459822 604338 495266 604574
rect 495502 604338 495586 604574
rect 495822 604338 531266 604574
rect 531502 604338 531586 604574
rect 531822 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 23546 601174
rect 23782 600938 23866 601174
rect 24102 600938 59546 601174
rect 59782 600938 59866 601174
rect 60102 600938 95546 601174
rect 95782 600938 95866 601174
rect 96102 600938 131546 601174
rect 131782 600938 131866 601174
rect 132102 600938 167546 601174
rect 167782 600938 167866 601174
rect 168102 600938 203546 601174
rect 203782 600938 203866 601174
rect 204102 600938 239546 601174
rect 239782 600938 239866 601174
rect 240102 600938 275546 601174
rect 275782 600938 275866 601174
rect 276102 600938 311546 601174
rect 311782 600938 311866 601174
rect 312102 600938 347546 601174
rect 347782 600938 347866 601174
rect 348102 600938 383546 601174
rect 383782 600938 383866 601174
rect 384102 600938 419546 601174
rect 419782 600938 419866 601174
rect 420102 600938 455546 601174
rect 455782 600938 455866 601174
rect 456102 600938 491546 601174
rect 491782 600938 491866 601174
rect 492102 600938 527546 601174
rect 527782 600938 527866 601174
rect 528102 600938 563546 601174
rect 563782 600938 563866 601174
rect 564102 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 23546 600854
rect 23782 600618 23866 600854
rect 24102 600618 59546 600854
rect 59782 600618 59866 600854
rect 60102 600618 95546 600854
rect 95782 600618 95866 600854
rect 96102 600618 131546 600854
rect 131782 600618 131866 600854
rect 132102 600618 167546 600854
rect 167782 600618 167866 600854
rect 168102 600618 203546 600854
rect 203782 600618 203866 600854
rect 204102 600618 239546 600854
rect 239782 600618 239866 600854
rect 240102 600618 275546 600854
rect 275782 600618 275866 600854
rect 276102 600618 311546 600854
rect 311782 600618 311866 600854
rect 312102 600618 347546 600854
rect 347782 600618 347866 600854
rect 348102 600618 383546 600854
rect 383782 600618 383866 600854
rect 384102 600618 419546 600854
rect 419782 600618 419866 600854
rect 420102 600618 455546 600854
rect 455782 600618 455866 600854
rect 456102 600618 491546 600854
rect 491782 600618 491866 600854
rect 492102 600618 527546 600854
rect 527782 600618 527866 600854
rect 528102 600618 563546 600854
rect 563782 600618 563866 600854
rect 564102 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 19826 597454
rect 20062 597218 20146 597454
rect 20382 597218 55826 597454
rect 56062 597218 56146 597454
rect 56382 597218 91826 597454
rect 92062 597218 92146 597454
rect 92382 597218 127826 597454
rect 128062 597218 128146 597454
rect 128382 597218 163826 597454
rect 164062 597218 164146 597454
rect 164382 597218 199826 597454
rect 200062 597218 200146 597454
rect 200382 597218 235826 597454
rect 236062 597218 236146 597454
rect 236382 597218 271826 597454
rect 272062 597218 272146 597454
rect 272382 597218 307826 597454
rect 308062 597218 308146 597454
rect 308382 597218 343826 597454
rect 344062 597218 344146 597454
rect 344382 597218 379826 597454
rect 380062 597218 380146 597454
rect 380382 597218 415826 597454
rect 416062 597218 416146 597454
rect 416382 597218 451826 597454
rect 452062 597218 452146 597454
rect 452382 597218 487826 597454
rect 488062 597218 488146 597454
rect 488382 597218 523826 597454
rect 524062 597218 524146 597454
rect 524382 597218 559826 597454
rect 560062 597218 560146 597454
rect 560382 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 19826 597134
rect 20062 596898 20146 597134
rect 20382 596898 55826 597134
rect 56062 596898 56146 597134
rect 56382 596898 91826 597134
rect 92062 596898 92146 597134
rect 92382 596898 127826 597134
rect 128062 596898 128146 597134
rect 128382 596898 163826 597134
rect 164062 596898 164146 597134
rect 164382 596898 199826 597134
rect 200062 596898 200146 597134
rect 200382 596898 235826 597134
rect 236062 596898 236146 597134
rect 236382 596898 271826 597134
rect 272062 596898 272146 597134
rect 272382 596898 307826 597134
rect 308062 596898 308146 597134
rect 308382 596898 343826 597134
rect 344062 596898 344146 597134
rect 344382 596898 379826 597134
rect 380062 596898 380146 597134
rect 380382 596898 415826 597134
rect 416062 596898 416146 597134
rect 416382 596898 451826 597134
rect 452062 596898 452146 597134
rect 452382 596898 487826 597134
rect 488062 596898 488146 597134
rect 488382 596898 523826 597134
rect 524062 596898 524146 597134
rect 524382 596898 559826 597134
rect 560062 596898 560146 597134
rect 560382 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 12986 590614
rect 13222 590378 13306 590614
rect 13542 590378 48986 590614
rect 49222 590378 49306 590614
rect 49542 590378 84986 590614
rect 85222 590378 85306 590614
rect 85542 590378 120986 590614
rect 121222 590378 121306 590614
rect 121542 590378 156986 590614
rect 157222 590378 157306 590614
rect 157542 590378 192986 590614
rect 193222 590378 193306 590614
rect 193542 590378 228986 590614
rect 229222 590378 229306 590614
rect 229542 590378 264986 590614
rect 265222 590378 265306 590614
rect 265542 590378 300986 590614
rect 301222 590378 301306 590614
rect 301542 590378 336986 590614
rect 337222 590378 337306 590614
rect 337542 590378 372986 590614
rect 373222 590378 373306 590614
rect 373542 590378 408986 590614
rect 409222 590378 409306 590614
rect 409542 590378 444986 590614
rect 445222 590378 445306 590614
rect 445542 590378 480986 590614
rect 481222 590378 481306 590614
rect 481542 590378 516986 590614
rect 517222 590378 517306 590614
rect 517542 590378 552986 590614
rect 553222 590378 553306 590614
rect 553542 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 12986 590294
rect 13222 590058 13306 590294
rect 13542 590058 48986 590294
rect 49222 590058 49306 590294
rect 49542 590058 84986 590294
rect 85222 590058 85306 590294
rect 85542 590058 120986 590294
rect 121222 590058 121306 590294
rect 121542 590058 156986 590294
rect 157222 590058 157306 590294
rect 157542 590058 192986 590294
rect 193222 590058 193306 590294
rect 193542 590058 228986 590294
rect 229222 590058 229306 590294
rect 229542 590058 264986 590294
rect 265222 590058 265306 590294
rect 265542 590058 300986 590294
rect 301222 590058 301306 590294
rect 301542 590058 336986 590294
rect 337222 590058 337306 590294
rect 337542 590058 372986 590294
rect 373222 590058 373306 590294
rect 373542 590058 408986 590294
rect 409222 590058 409306 590294
rect 409542 590058 444986 590294
rect 445222 590058 445306 590294
rect 445542 590058 480986 590294
rect 481222 590058 481306 590294
rect 481542 590058 516986 590294
rect 517222 590058 517306 590294
rect 517542 590058 552986 590294
rect 553222 590058 553306 590294
rect 553542 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 9266 586894
rect 9502 586658 9586 586894
rect 9822 586658 45266 586894
rect 45502 586658 45586 586894
rect 45822 586658 81266 586894
rect 81502 586658 81586 586894
rect 81822 586658 117266 586894
rect 117502 586658 117586 586894
rect 117822 586658 153266 586894
rect 153502 586658 153586 586894
rect 153822 586658 189266 586894
rect 189502 586658 189586 586894
rect 189822 586658 225266 586894
rect 225502 586658 225586 586894
rect 225822 586658 261266 586894
rect 261502 586658 261586 586894
rect 261822 586658 297266 586894
rect 297502 586658 297586 586894
rect 297822 586658 333266 586894
rect 333502 586658 333586 586894
rect 333822 586658 369266 586894
rect 369502 586658 369586 586894
rect 369822 586658 405266 586894
rect 405502 586658 405586 586894
rect 405822 586658 441266 586894
rect 441502 586658 441586 586894
rect 441822 586658 477266 586894
rect 477502 586658 477586 586894
rect 477822 586658 513266 586894
rect 513502 586658 513586 586894
rect 513822 586658 549266 586894
rect 549502 586658 549586 586894
rect 549822 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 9266 586574
rect 9502 586338 9586 586574
rect 9822 586338 45266 586574
rect 45502 586338 45586 586574
rect 45822 586338 81266 586574
rect 81502 586338 81586 586574
rect 81822 586338 117266 586574
rect 117502 586338 117586 586574
rect 117822 586338 153266 586574
rect 153502 586338 153586 586574
rect 153822 586338 189266 586574
rect 189502 586338 189586 586574
rect 189822 586338 225266 586574
rect 225502 586338 225586 586574
rect 225822 586338 261266 586574
rect 261502 586338 261586 586574
rect 261822 586338 297266 586574
rect 297502 586338 297586 586574
rect 297822 586338 333266 586574
rect 333502 586338 333586 586574
rect 333822 586338 369266 586574
rect 369502 586338 369586 586574
rect 369822 586338 405266 586574
rect 405502 586338 405586 586574
rect 405822 586338 441266 586574
rect 441502 586338 441586 586574
rect 441822 586338 477266 586574
rect 477502 586338 477586 586574
rect 477822 586338 513266 586574
rect 513502 586338 513586 586574
rect 513822 586338 549266 586574
rect 549502 586338 549586 586574
rect 549822 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 5546 583174
rect 5782 582938 5866 583174
rect 6102 582938 41546 583174
rect 41782 582938 41866 583174
rect 42102 582938 77546 583174
rect 77782 582938 77866 583174
rect 78102 582938 113546 583174
rect 113782 582938 113866 583174
rect 114102 582938 149546 583174
rect 149782 582938 149866 583174
rect 150102 582938 185546 583174
rect 185782 582938 185866 583174
rect 186102 582938 221546 583174
rect 221782 582938 221866 583174
rect 222102 582938 257546 583174
rect 257782 582938 257866 583174
rect 258102 582938 293546 583174
rect 293782 582938 293866 583174
rect 294102 582938 329546 583174
rect 329782 582938 329866 583174
rect 330102 582938 365546 583174
rect 365782 582938 365866 583174
rect 366102 582938 401546 583174
rect 401782 582938 401866 583174
rect 402102 582938 437546 583174
rect 437782 582938 437866 583174
rect 438102 582938 473546 583174
rect 473782 582938 473866 583174
rect 474102 582938 509546 583174
rect 509782 582938 509866 583174
rect 510102 582938 545546 583174
rect 545782 582938 545866 583174
rect 546102 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 5546 582854
rect 5782 582618 5866 582854
rect 6102 582618 41546 582854
rect 41782 582618 41866 582854
rect 42102 582618 77546 582854
rect 77782 582618 77866 582854
rect 78102 582618 113546 582854
rect 113782 582618 113866 582854
rect 114102 582618 149546 582854
rect 149782 582618 149866 582854
rect 150102 582618 185546 582854
rect 185782 582618 185866 582854
rect 186102 582618 221546 582854
rect 221782 582618 221866 582854
rect 222102 582618 257546 582854
rect 257782 582618 257866 582854
rect 258102 582618 293546 582854
rect 293782 582618 293866 582854
rect 294102 582618 329546 582854
rect 329782 582618 329866 582854
rect 330102 582618 365546 582854
rect 365782 582618 365866 582854
rect 366102 582618 401546 582854
rect 401782 582618 401866 582854
rect 402102 582618 437546 582854
rect 437782 582618 437866 582854
rect 438102 582618 473546 582854
rect 473782 582618 473866 582854
rect 474102 582618 509546 582854
rect 509782 582618 509866 582854
rect 510102 582618 545546 582854
rect 545782 582618 545866 582854
rect 546102 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 1826 579454
rect 2062 579218 2146 579454
rect 2382 579218 37826 579454
rect 38062 579218 38146 579454
rect 38382 579218 73826 579454
rect 74062 579218 74146 579454
rect 74382 579218 109826 579454
rect 110062 579218 110146 579454
rect 110382 579218 145826 579454
rect 146062 579218 146146 579454
rect 146382 579218 181826 579454
rect 182062 579218 182146 579454
rect 182382 579218 217826 579454
rect 218062 579218 218146 579454
rect 218382 579218 253826 579454
rect 254062 579218 254146 579454
rect 254382 579218 289826 579454
rect 290062 579218 290146 579454
rect 290382 579218 325826 579454
rect 326062 579218 326146 579454
rect 326382 579218 361826 579454
rect 362062 579218 362146 579454
rect 362382 579218 397826 579454
rect 398062 579218 398146 579454
rect 398382 579218 433826 579454
rect 434062 579218 434146 579454
rect 434382 579218 469826 579454
rect 470062 579218 470146 579454
rect 470382 579218 505826 579454
rect 506062 579218 506146 579454
rect 506382 579218 541826 579454
rect 542062 579218 542146 579454
rect 542382 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 1826 579134
rect 2062 578898 2146 579134
rect 2382 578898 37826 579134
rect 38062 578898 38146 579134
rect 38382 578898 73826 579134
rect 74062 578898 74146 579134
rect 74382 578898 109826 579134
rect 110062 578898 110146 579134
rect 110382 578898 145826 579134
rect 146062 578898 146146 579134
rect 146382 578898 181826 579134
rect 182062 578898 182146 579134
rect 182382 578898 217826 579134
rect 218062 578898 218146 579134
rect 218382 578898 253826 579134
rect 254062 578898 254146 579134
rect 254382 578898 289826 579134
rect 290062 578898 290146 579134
rect 290382 578898 325826 579134
rect 326062 578898 326146 579134
rect 326382 578898 361826 579134
rect 362062 578898 362146 579134
rect 362382 578898 397826 579134
rect 398062 578898 398146 579134
rect 398382 578898 433826 579134
rect 434062 578898 434146 579134
rect 434382 578898 469826 579134
rect 470062 578898 470146 579134
rect 470382 578898 505826 579134
rect 506062 578898 506146 579134
rect 506382 578898 541826 579134
rect 542062 578898 542146 579134
rect 542382 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 30986 572614
rect 31222 572378 31306 572614
rect 31542 572378 66986 572614
rect 67222 572378 67306 572614
rect 67542 572378 102986 572614
rect 103222 572378 103306 572614
rect 103542 572378 138986 572614
rect 139222 572378 139306 572614
rect 139542 572378 174986 572614
rect 175222 572378 175306 572614
rect 175542 572378 210986 572614
rect 211222 572378 211306 572614
rect 211542 572378 246986 572614
rect 247222 572378 247306 572614
rect 247542 572378 282986 572614
rect 283222 572378 283306 572614
rect 283542 572378 318986 572614
rect 319222 572378 319306 572614
rect 319542 572378 354986 572614
rect 355222 572378 355306 572614
rect 355542 572378 390986 572614
rect 391222 572378 391306 572614
rect 391542 572378 426986 572614
rect 427222 572378 427306 572614
rect 427542 572378 462986 572614
rect 463222 572378 463306 572614
rect 463542 572378 498986 572614
rect 499222 572378 499306 572614
rect 499542 572378 534986 572614
rect 535222 572378 535306 572614
rect 535542 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 30986 572294
rect 31222 572058 31306 572294
rect 31542 572058 66986 572294
rect 67222 572058 67306 572294
rect 67542 572058 102986 572294
rect 103222 572058 103306 572294
rect 103542 572058 138986 572294
rect 139222 572058 139306 572294
rect 139542 572058 174986 572294
rect 175222 572058 175306 572294
rect 175542 572058 210986 572294
rect 211222 572058 211306 572294
rect 211542 572058 246986 572294
rect 247222 572058 247306 572294
rect 247542 572058 282986 572294
rect 283222 572058 283306 572294
rect 283542 572058 318986 572294
rect 319222 572058 319306 572294
rect 319542 572058 354986 572294
rect 355222 572058 355306 572294
rect 355542 572058 390986 572294
rect 391222 572058 391306 572294
rect 391542 572058 426986 572294
rect 427222 572058 427306 572294
rect 427542 572058 462986 572294
rect 463222 572058 463306 572294
rect 463542 572058 498986 572294
rect 499222 572058 499306 572294
rect 499542 572058 534986 572294
rect 535222 572058 535306 572294
rect 535542 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 27266 568894
rect 27502 568658 27586 568894
rect 27822 568658 63266 568894
rect 63502 568658 63586 568894
rect 63822 568658 99266 568894
rect 99502 568658 99586 568894
rect 99822 568658 135266 568894
rect 135502 568658 135586 568894
rect 135822 568658 171266 568894
rect 171502 568658 171586 568894
rect 171822 568658 207266 568894
rect 207502 568658 207586 568894
rect 207822 568658 243266 568894
rect 243502 568658 243586 568894
rect 243822 568658 279266 568894
rect 279502 568658 279586 568894
rect 279822 568658 315266 568894
rect 315502 568658 315586 568894
rect 315822 568658 351266 568894
rect 351502 568658 351586 568894
rect 351822 568658 387266 568894
rect 387502 568658 387586 568894
rect 387822 568658 423266 568894
rect 423502 568658 423586 568894
rect 423822 568658 459266 568894
rect 459502 568658 459586 568894
rect 459822 568658 495266 568894
rect 495502 568658 495586 568894
rect 495822 568658 531266 568894
rect 531502 568658 531586 568894
rect 531822 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 27266 568574
rect 27502 568338 27586 568574
rect 27822 568338 63266 568574
rect 63502 568338 63586 568574
rect 63822 568338 99266 568574
rect 99502 568338 99586 568574
rect 99822 568338 135266 568574
rect 135502 568338 135586 568574
rect 135822 568338 171266 568574
rect 171502 568338 171586 568574
rect 171822 568338 207266 568574
rect 207502 568338 207586 568574
rect 207822 568338 243266 568574
rect 243502 568338 243586 568574
rect 243822 568338 279266 568574
rect 279502 568338 279586 568574
rect 279822 568338 315266 568574
rect 315502 568338 315586 568574
rect 315822 568338 351266 568574
rect 351502 568338 351586 568574
rect 351822 568338 387266 568574
rect 387502 568338 387586 568574
rect 387822 568338 423266 568574
rect 423502 568338 423586 568574
rect 423822 568338 459266 568574
rect 459502 568338 459586 568574
rect 459822 568338 495266 568574
rect 495502 568338 495586 568574
rect 495822 568338 531266 568574
rect 531502 568338 531586 568574
rect 531822 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 23546 565174
rect 23782 564938 23866 565174
rect 24102 564938 59546 565174
rect 59782 564938 59866 565174
rect 60102 564938 95546 565174
rect 95782 564938 95866 565174
rect 96102 564938 131546 565174
rect 131782 564938 131866 565174
rect 132102 564938 167546 565174
rect 167782 564938 167866 565174
rect 168102 564938 203546 565174
rect 203782 564938 203866 565174
rect 204102 564938 239546 565174
rect 239782 564938 239866 565174
rect 240102 564938 275546 565174
rect 275782 564938 275866 565174
rect 276102 564938 311546 565174
rect 311782 564938 311866 565174
rect 312102 564938 347546 565174
rect 347782 564938 347866 565174
rect 348102 564938 383546 565174
rect 383782 564938 383866 565174
rect 384102 564938 419546 565174
rect 419782 564938 419866 565174
rect 420102 564938 455546 565174
rect 455782 564938 455866 565174
rect 456102 564938 491546 565174
rect 491782 564938 491866 565174
rect 492102 564938 527546 565174
rect 527782 564938 527866 565174
rect 528102 564938 563546 565174
rect 563782 564938 563866 565174
rect 564102 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 23546 564854
rect 23782 564618 23866 564854
rect 24102 564618 59546 564854
rect 59782 564618 59866 564854
rect 60102 564618 95546 564854
rect 95782 564618 95866 564854
rect 96102 564618 131546 564854
rect 131782 564618 131866 564854
rect 132102 564618 167546 564854
rect 167782 564618 167866 564854
rect 168102 564618 203546 564854
rect 203782 564618 203866 564854
rect 204102 564618 239546 564854
rect 239782 564618 239866 564854
rect 240102 564618 275546 564854
rect 275782 564618 275866 564854
rect 276102 564618 311546 564854
rect 311782 564618 311866 564854
rect 312102 564618 347546 564854
rect 347782 564618 347866 564854
rect 348102 564618 383546 564854
rect 383782 564618 383866 564854
rect 384102 564618 419546 564854
rect 419782 564618 419866 564854
rect 420102 564618 455546 564854
rect 455782 564618 455866 564854
rect 456102 564618 491546 564854
rect 491782 564618 491866 564854
rect 492102 564618 527546 564854
rect 527782 564618 527866 564854
rect 528102 564618 563546 564854
rect 563782 564618 563866 564854
rect 564102 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 19826 561454
rect 20062 561218 20146 561454
rect 20382 561218 55826 561454
rect 56062 561218 56146 561454
rect 56382 561218 91826 561454
rect 92062 561218 92146 561454
rect 92382 561218 127826 561454
rect 128062 561218 128146 561454
rect 128382 561218 163826 561454
rect 164062 561218 164146 561454
rect 164382 561218 199826 561454
rect 200062 561218 200146 561454
rect 200382 561218 235826 561454
rect 236062 561218 236146 561454
rect 236382 561218 271826 561454
rect 272062 561218 272146 561454
rect 272382 561218 307826 561454
rect 308062 561218 308146 561454
rect 308382 561218 343826 561454
rect 344062 561218 344146 561454
rect 344382 561218 379826 561454
rect 380062 561218 380146 561454
rect 380382 561218 415826 561454
rect 416062 561218 416146 561454
rect 416382 561218 451826 561454
rect 452062 561218 452146 561454
rect 452382 561218 487826 561454
rect 488062 561218 488146 561454
rect 488382 561218 523826 561454
rect 524062 561218 524146 561454
rect 524382 561218 559826 561454
rect 560062 561218 560146 561454
rect 560382 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 19826 561134
rect 20062 560898 20146 561134
rect 20382 560898 55826 561134
rect 56062 560898 56146 561134
rect 56382 560898 91826 561134
rect 92062 560898 92146 561134
rect 92382 560898 127826 561134
rect 128062 560898 128146 561134
rect 128382 560898 163826 561134
rect 164062 560898 164146 561134
rect 164382 560898 199826 561134
rect 200062 560898 200146 561134
rect 200382 560898 235826 561134
rect 236062 560898 236146 561134
rect 236382 560898 271826 561134
rect 272062 560898 272146 561134
rect 272382 560898 307826 561134
rect 308062 560898 308146 561134
rect 308382 560898 343826 561134
rect 344062 560898 344146 561134
rect 344382 560898 379826 561134
rect 380062 560898 380146 561134
rect 380382 560898 415826 561134
rect 416062 560898 416146 561134
rect 416382 560898 451826 561134
rect 452062 560898 452146 561134
rect 452382 560898 487826 561134
rect 488062 560898 488146 561134
rect 488382 560898 523826 561134
rect 524062 560898 524146 561134
rect 524382 560898 559826 561134
rect 560062 560898 560146 561134
rect 560382 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 12986 554614
rect 13222 554378 13306 554614
rect 13542 554378 48986 554614
rect 49222 554378 49306 554614
rect 49542 554378 84986 554614
rect 85222 554378 85306 554614
rect 85542 554378 120986 554614
rect 121222 554378 121306 554614
rect 121542 554378 156986 554614
rect 157222 554378 157306 554614
rect 157542 554378 192986 554614
rect 193222 554378 193306 554614
rect 193542 554378 228986 554614
rect 229222 554378 229306 554614
rect 229542 554378 264986 554614
rect 265222 554378 265306 554614
rect 265542 554378 300986 554614
rect 301222 554378 301306 554614
rect 301542 554378 336986 554614
rect 337222 554378 337306 554614
rect 337542 554378 372986 554614
rect 373222 554378 373306 554614
rect 373542 554378 408986 554614
rect 409222 554378 409306 554614
rect 409542 554378 444986 554614
rect 445222 554378 445306 554614
rect 445542 554378 480986 554614
rect 481222 554378 481306 554614
rect 481542 554378 516986 554614
rect 517222 554378 517306 554614
rect 517542 554378 552986 554614
rect 553222 554378 553306 554614
rect 553542 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 12986 554294
rect 13222 554058 13306 554294
rect 13542 554058 48986 554294
rect 49222 554058 49306 554294
rect 49542 554058 84986 554294
rect 85222 554058 85306 554294
rect 85542 554058 120986 554294
rect 121222 554058 121306 554294
rect 121542 554058 156986 554294
rect 157222 554058 157306 554294
rect 157542 554058 192986 554294
rect 193222 554058 193306 554294
rect 193542 554058 228986 554294
rect 229222 554058 229306 554294
rect 229542 554058 264986 554294
rect 265222 554058 265306 554294
rect 265542 554058 300986 554294
rect 301222 554058 301306 554294
rect 301542 554058 336986 554294
rect 337222 554058 337306 554294
rect 337542 554058 372986 554294
rect 373222 554058 373306 554294
rect 373542 554058 408986 554294
rect 409222 554058 409306 554294
rect 409542 554058 444986 554294
rect 445222 554058 445306 554294
rect 445542 554058 480986 554294
rect 481222 554058 481306 554294
rect 481542 554058 516986 554294
rect 517222 554058 517306 554294
rect 517542 554058 552986 554294
rect 553222 554058 553306 554294
rect 553542 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 9266 550894
rect 9502 550658 9586 550894
rect 9822 550658 45266 550894
rect 45502 550658 45586 550894
rect 45822 550658 81266 550894
rect 81502 550658 81586 550894
rect 81822 550658 117266 550894
rect 117502 550658 117586 550894
rect 117822 550658 153266 550894
rect 153502 550658 153586 550894
rect 153822 550658 189266 550894
rect 189502 550658 189586 550894
rect 189822 550658 225266 550894
rect 225502 550658 225586 550894
rect 225822 550658 261266 550894
rect 261502 550658 261586 550894
rect 261822 550658 297266 550894
rect 297502 550658 297586 550894
rect 297822 550658 333266 550894
rect 333502 550658 333586 550894
rect 333822 550658 369266 550894
rect 369502 550658 369586 550894
rect 369822 550658 405266 550894
rect 405502 550658 405586 550894
rect 405822 550658 441266 550894
rect 441502 550658 441586 550894
rect 441822 550658 477266 550894
rect 477502 550658 477586 550894
rect 477822 550658 513266 550894
rect 513502 550658 513586 550894
rect 513822 550658 549266 550894
rect 549502 550658 549586 550894
rect 549822 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 9266 550574
rect 9502 550338 9586 550574
rect 9822 550338 45266 550574
rect 45502 550338 45586 550574
rect 45822 550338 81266 550574
rect 81502 550338 81586 550574
rect 81822 550338 117266 550574
rect 117502 550338 117586 550574
rect 117822 550338 153266 550574
rect 153502 550338 153586 550574
rect 153822 550338 189266 550574
rect 189502 550338 189586 550574
rect 189822 550338 225266 550574
rect 225502 550338 225586 550574
rect 225822 550338 261266 550574
rect 261502 550338 261586 550574
rect 261822 550338 297266 550574
rect 297502 550338 297586 550574
rect 297822 550338 333266 550574
rect 333502 550338 333586 550574
rect 333822 550338 369266 550574
rect 369502 550338 369586 550574
rect 369822 550338 405266 550574
rect 405502 550338 405586 550574
rect 405822 550338 441266 550574
rect 441502 550338 441586 550574
rect 441822 550338 477266 550574
rect 477502 550338 477586 550574
rect 477822 550338 513266 550574
rect 513502 550338 513586 550574
rect 513822 550338 549266 550574
rect 549502 550338 549586 550574
rect 549822 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 5546 547174
rect 5782 546938 5866 547174
rect 6102 546938 41546 547174
rect 41782 546938 41866 547174
rect 42102 546938 77546 547174
rect 77782 546938 77866 547174
rect 78102 546938 113546 547174
rect 113782 546938 113866 547174
rect 114102 546938 149546 547174
rect 149782 546938 149866 547174
rect 150102 546938 185546 547174
rect 185782 546938 185866 547174
rect 186102 546938 221546 547174
rect 221782 546938 221866 547174
rect 222102 546938 257546 547174
rect 257782 546938 257866 547174
rect 258102 546938 293546 547174
rect 293782 546938 293866 547174
rect 294102 546938 329546 547174
rect 329782 546938 329866 547174
rect 330102 546938 365546 547174
rect 365782 546938 365866 547174
rect 366102 546938 401546 547174
rect 401782 546938 401866 547174
rect 402102 546938 437546 547174
rect 437782 546938 437866 547174
rect 438102 546938 473546 547174
rect 473782 546938 473866 547174
rect 474102 546938 509546 547174
rect 509782 546938 509866 547174
rect 510102 546938 545546 547174
rect 545782 546938 545866 547174
rect 546102 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 5546 546854
rect 5782 546618 5866 546854
rect 6102 546618 41546 546854
rect 41782 546618 41866 546854
rect 42102 546618 77546 546854
rect 77782 546618 77866 546854
rect 78102 546618 113546 546854
rect 113782 546618 113866 546854
rect 114102 546618 149546 546854
rect 149782 546618 149866 546854
rect 150102 546618 185546 546854
rect 185782 546618 185866 546854
rect 186102 546618 221546 546854
rect 221782 546618 221866 546854
rect 222102 546618 257546 546854
rect 257782 546618 257866 546854
rect 258102 546618 293546 546854
rect 293782 546618 293866 546854
rect 294102 546618 329546 546854
rect 329782 546618 329866 546854
rect 330102 546618 365546 546854
rect 365782 546618 365866 546854
rect 366102 546618 401546 546854
rect 401782 546618 401866 546854
rect 402102 546618 437546 546854
rect 437782 546618 437866 546854
rect 438102 546618 473546 546854
rect 473782 546618 473866 546854
rect 474102 546618 509546 546854
rect 509782 546618 509866 546854
rect 510102 546618 545546 546854
rect 545782 546618 545866 546854
rect 546102 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 1826 543454
rect 2062 543218 2146 543454
rect 2382 543218 37826 543454
rect 38062 543218 38146 543454
rect 38382 543218 73826 543454
rect 74062 543218 74146 543454
rect 74382 543218 109826 543454
rect 110062 543218 110146 543454
rect 110382 543218 145826 543454
rect 146062 543218 146146 543454
rect 146382 543218 181826 543454
rect 182062 543218 182146 543454
rect 182382 543218 217826 543454
rect 218062 543218 218146 543454
rect 218382 543218 253826 543454
rect 254062 543218 254146 543454
rect 254382 543218 289826 543454
rect 290062 543218 290146 543454
rect 290382 543218 325826 543454
rect 326062 543218 326146 543454
rect 326382 543218 361826 543454
rect 362062 543218 362146 543454
rect 362382 543218 397826 543454
rect 398062 543218 398146 543454
rect 398382 543218 433826 543454
rect 434062 543218 434146 543454
rect 434382 543218 469826 543454
rect 470062 543218 470146 543454
rect 470382 543218 505826 543454
rect 506062 543218 506146 543454
rect 506382 543218 541826 543454
rect 542062 543218 542146 543454
rect 542382 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 1826 543134
rect 2062 542898 2146 543134
rect 2382 542898 37826 543134
rect 38062 542898 38146 543134
rect 38382 542898 73826 543134
rect 74062 542898 74146 543134
rect 74382 542898 109826 543134
rect 110062 542898 110146 543134
rect 110382 542898 145826 543134
rect 146062 542898 146146 543134
rect 146382 542898 181826 543134
rect 182062 542898 182146 543134
rect 182382 542898 217826 543134
rect 218062 542898 218146 543134
rect 218382 542898 253826 543134
rect 254062 542898 254146 543134
rect 254382 542898 289826 543134
rect 290062 542898 290146 543134
rect 290382 542898 325826 543134
rect 326062 542898 326146 543134
rect 326382 542898 361826 543134
rect 362062 542898 362146 543134
rect 362382 542898 397826 543134
rect 398062 542898 398146 543134
rect 398382 542898 433826 543134
rect 434062 542898 434146 543134
rect 434382 542898 469826 543134
rect 470062 542898 470146 543134
rect 470382 542898 505826 543134
rect 506062 542898 506146 543134
rect 506382 542898 541826 543134
rect 542062 542898 542146 543134
rect 542382 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 30986 536614
rect 31222 536378 31306 536614
rect 31542 536378 66986 536614
rect 67222 536378 67306 536614
rect 67542 536378 102986 536614
rect 103222 536378 103306 536614
rect 103542 536378 138986 536614
rect 139222 536378 139306 536614
rect 139542 536378 174986 536614
rect 175222 536378 175306 536614
rect 175542 536378 210986 536614
rect 211222 536378 211306 536614
rect 211542 536378 246986 536614
rect 247222 536378 247306 536614
rect 247542 536378 282986 536614
rect 283222 536378 283306 536614
rect 283542 536378 318986 536614
rect 319222 536378 319306 536614
rect 319542 536378 354986 536614
rect 355222 536378 355306 536614
rect 355542 536378 390986 536614
rect 391222 536378 391306 536614
rect 391542 536378 426986 536614
rect 427222 536378 427306 536614
rect 427542 536378 462986 536614
rect 463222 536378 463306 536614
rect 463542 536378 498986 536614
rect 499222 536378 499306 536614
rect 499542 536378 534986 536614
rect 535222 536378 535306 536614
rect 535542 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 30986 536294
rect 31222 536058 31306 536294
rect 31542 536058 66986 536294
rect 67222 536058 67306 536294
rect 67542 536058 102986 536294
rect 103222 536058 103306 536294
rect 103542 536058 138986 536294
rect 139222 536058 139306 536294
rect 139542 536058 174986 536294
rect 175222 536058 175306 536294
rect 175542 536058 210986 536294
rect 211222 536058 211306 536294
rect 211542 536058 246986 536294
rect 247222 536058 247306 536294
rect 247542 536058 282986 536294
rect 283222 536058 283306 536294
rect 283542 536058 318986 536294
rect 319222 536058 319306 536294
rect 319542 536058 354986 536294
rect 355222 536058 355306 536294
rect 355542 536058 390986 536294
rect 391222 536058 391306 536294
rect 391542 536058 426986 536294
rect 427222 536058 427306 536294
rect 427542 536058 462986 536294
rect 463222 536058 463306 536294
rect 463542 536058 498986 536294
rect 499222 536058 499306 536294
rect 499542 536058 534986 536294
rect 535222 536058 535306 536294
rect 535542 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 27266 532894
rect 27502 532658 27586 532894
rect 27822 532658 63266 532894
rect 63502 532658 63586 532894
rect 63822 532658 99266 532894
rect 99502 532658 99586 532894
rect 99822 532658 135266 532894
rect 135502 532658 135586 532894
rect 135822 532658 171266 532894
rect 171502 532658 171586 532894
rect 171822 532658 207266 532894
rect 207502 532658 207586 532894
rect 207822 532658 243266 532894
rect 243502 532658 243586 532894
rect 243822 532658 279266 532894
rect 279502 532658 279586 532894
rect 279822 532658 315266 532894
rect 315502 532658 315586 532894
rect 315822 532658 351266 532894
rect 351502 532658 351586 532894
rect 351822 532658 387266 532894
rect 387502 532658 387586 532894
rect 387822 532658 423266 532894
rect 423502 532658 423586 532894
rect 423822 532658 459266 532894
rect 459502 532658 459586 532894
rect 459822 532658 495266 532894
rect 495502 532658 495586 532894
rect 495822 532658 531266 532894
rect 531502 532658 531586 532894
rect 531822 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 27266 532574
rect 27502 532338 27586 532574
rect 27822 532338 63266 532574
rect 63502 532338 63586 532574
rect 63822 532338 99266 532574
rect 99502 532338 99586 532574
rect 99822 532338 135266 532574
rect 135502 532338 135586 532574
rect 135822 532338 171266 532574
rect 171502 532338 171586 532574
rect 171822 532338 207266 532574
rect 207502 532338 207586 532574
rect 207822 532338 243266 532574
rect 243502 532338 243586 532574
rect 243822 532338 279266 532574
rect 279502 532338 279586 532574
rect 279822 532338 315266 532574
rect 315502 532338 315586 532574
rect 315822 532338 351266 532574
rect 351502 532338 351586 532574
rect 351822 532338 387266 532574
rect 387502 532338 387586 532574
rect 387822 532338 423266 532574
rect 423502 532338 423586 532574
rect 423822 532338 459266 532574
rect 459502 532338 459586 532574
rect 459822 532338 495266 532574
rect 495502 532338 495586 532574
rect 495822 532338 531266 532574
rect 531502 532338 531586 532574
rect 531822 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 23546 529174
rect 23782 528938 23866 529174
rect 24102 528938 59546 529174
rect 59782 528938 59866 529174
rect 60102 528938 95546 529174
rect 95782 528938 95866 529174
rect 96102 528938 131546 529174
rect 131782 528938 131866 529174
rect 132102 528938 167546 529174
rect 167782 528938 167866 529174
rect 168102 528938 203546 529174
rect 203782 528938 203866 529174
rect 204102 528938 239546 529174
rect 239782 528938 239866 529174
rect 240102 528938 275546 529174
rect 275782 528938 275866 529174
rect 276102 528938 311546 529174
rect 311782 528938 311866 529174
rect 312102 528938 347546 529174
rect 347782 528938 347866 529174
rect 348102 528938 383546 529174
rect 383782 528938 383866 529174
rect 384102 528938 419546 529174
rect 419782 528938 419866 529174
rect 420102 528938 455546 529174
rect 455782 528938 455866 529174
rect 456102 528938 491546 529174
rect 491782 528938 491866 529174
rect 492102 528938 527546 529174
rect 527782 528938 527866 529174
rect 528102 528938 563546 529174
rect 563782 528938 563866 529174
rect 564102 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 23546 528854
rect 23782 528618 23866 528854
rect 24102 528618 59546 528854
rect 59782 528618 59866 528854
rect 60102 528618 95546 528854
rect 95782 528618 95866 528854
rect 96102 528618 131546 528854
rect 131782 528618 131866 528854
rect 132102 528618 167546 528854
rect 167782 528618 167866 528854
rect 168102 528618 203546 528854
rect 203782 528618 203866 528854
rect 204102 528618 239546 528854
rect 239782 528618 239866 528854
rect 240102 528618 275546 528854
rect 275782 528618 275866 528854
rect 276102 528618 311546 528854
rect 311782 528618 311866 528854
rect 312102 528618 347546 528854
rect 347782 528618 347866 528854
rect 348102 528618 383546 528854
rect 383782 528618 383866 528854
rect 384102 528618 419546 528854
rect 419782 528618 419866 528854
rect 420102 528618 455546 528854
rect 455782 528618 455866 528854
rect 456102 528618 491546 528854
rect 491782 528618 491866 528854
rect 492102 528618 527546 528854
rect 527782 528618 527866 528854
rect 528102 528618 563546 528854
rect 563782 528618 563866 528854
rect 564102 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 19826 525454
rect 20062 525218 20146 525454
rect 20382 525218 55826 525454
rect 56062 525218 56146 525454
rect 56382 525218 91826 525454
rect 92062 525218 92146 525454
rect 92382 525218 127826 525454
rect 128062 525218 128146 525454
rect 128382 525218 163826 525454
rect 164062 525218 164146 525454
rect 164382 525218 199826 525454
rect 200062 525218 200146 525454
rect 200382 525218 235826 525454
rect 236062 525218 236146 525454
rect 236382 525218 271826 525454
rect 272062 525218 272146 525454
rect 272382 525218 307826 525454
rect 308062 525218 308146 525454
rect 308382 525218 343826 525454
rect 344062 525218 344146 525454
rect 344382 525218 379826 525454
rect 380062 525218 380146 525454
rect 380382 525218 415826 525454
rect 416062 525218 416146 525454
rect 416382 525218 451826 525454
rect 452062 525218 452146 525454
rect 452382 525218 487826 525454
rect 488062 525218 488146 525454
rect 488382 525218 523826 525454
rect 524062 525218 524146 525454
rect 524382 525218 559826 525454
rect 560062 525218 560146 525454
rect 560382 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 19826 525134
rect 20062 524898 20146 525134
rect 20382 524898 55826 525134
rect 56062 524898 56146 525134
rect 56382 524898 91826 525134
rect 92062 524898 92146 525134
rect 92382 524898 127826 525134
rect 128062 524898 128146 525134
rect 128382 524898 163826 525134
rect 164062 524898 164146 525134
rect 164382 524898 199826 525134
rect 200062 524898 200146 525134
rect 200382 524898 235826 525134
rect 236062 524898 236146 525134
rect 236382 524898 271826 525134
rect 272062 524898 272146 525134
rect 272382 524898 307826 525134
rect 308062 524898 308146 525134
rect 308382 524898 343826 525134
rect 344062 524898 344146 525134
rect 344382 524898 379826 525134
rect 380062 524898 380146 525134
rect 380382 524898 415826 525134
rect 416062 524898 416146 525134
rect 416382 524898 451826 525134
rect 452062 524898 452146 525134
rect 452382 524898 487826 525134
rect 488062 524898 488146 525134
rect 488382 524898 523826 525134
rect 524062 524898 524146 525134
rect 524382 524898 559826 525134
rect 560062 524898 560146 525134
rect 560382 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 12986 518614
rect 13222 518378 13306 518614
rect 13542 518378 48986 518614
rect 49222 518378 49306 518614
rect 49542 518378 84986 518614
rect 85222 518378 85306 518614
rect 85542 518378 120986 518614
rect 121222 518378 121306 518614
rect 121542 518378 156986 518614
rect 157222 518378 157306 518614
rect 157542 518378 192986 518614
rect 193222 518378 193306 518614
rect 193542 518378 228986 518614
rect 229222 518378 229306 518614
rect 229542 518378 264986 518614
rect 265222 518378 265306 518614
rect 265542 518378 300986 518614
rect 301222 518378 301306 518614
rect 301542 518378 336986 518614
rect 337222 518378 337306 518614
rect 337542 518378 372986 518614
rect 373222 518378 373306 518614
rect 373542 518378 408986 518614
rect 409222 518378 409306 518614
rect 409542 518378 444986 518614
rect 445222 518378 445306 518614
rect 445542 518378 480986 518614
rect 481222 518378 481306 518614
rect 481542 518378 516986 518614
rect 517222 518378 517306 518614
rect 517542 518378 552986 518614
rect 553222 518378 553306 518614
rect 553542 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 12986 518294
rect 13222 518058 13306 518294
rect 13542 518058 48986 518294
rect 49222 518058 49306 518294
rect 49542 518058 84986 518294
rect 85222 518058 85306 518294
rect 85542 518058 120986 518294
rect 121222 518058 121306 518294
rect 121542 518058 156986 518294
rect 157222 518058 157306 518294
rect 157542 518058 192986 518294
rect 193222 518058 193306 518294
rect 193542 518058 228986 518294
rect 229222 518058 229306 518294
rect 229542 518058 264986 518294
rect 265222 518058 265306 518294
rect 265542 518058 300986 518294
rect 301222 518058 301306 518294
rect 301542 518058 336986 518294
rect 337222 518058 337306 518294
rect 337542 518058 372986 518294
rect 373222 518058 373306 518294
rect 373542 518058 408986 518294
rect 409222 518058 409306 518294
rect 409542 518058 444986 518294
rect 445222 518058 445306 518294
rect 445542 518058 480986 518294
rect 481222 518058 481306 518294
rect 481542 518058 516986 518294
rect 517222 518058 517306 518294
rect 517542 518058 552986 518294
rect 553222 518058 553306 518294
rect 553542 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 9266 514894
rect 9502 514658 9586 514894
rect 9822 514658 45266 514894
rect 45502 514658 45586 514894
rect 45822 514658 81266 514894
rect 81502 514658 81586 514894
rect 81822 514658 117266 514894
rect 117502 514658 117586 514894
rect 117822 514658 153266 514894
rect 153502 514658 153586 514894
rect 153822 514658 189266 514894
rect 189502 514658 189586 514894
rect 189822 514658 225266 514894
rect 225502 514658 225586 514894
rect 225822 514658 261266 514894
rect 261502 514658 261586 514894
rect 261822 514658 297266 514894
rect 297502 514658 297586 514894
rect 297822 514658 333266 514894
rect 333502 514658 333586 514894
rect 333822 514658 369266 514894
rect 369502 514658 369586 514894
rect 369822 514658 405266 514894
rect 405502 514658 405586 514894
rect 405822 514658 441266 514894
rect 441502 514658 441586 514894
rect 441822 514658 477266 514894
rect 477502 514658 477586 514894
rect 477822 514658 513266 514894
rect 513502 514658 513586 514894
rect 513822 514658 549266 514894
rect 549502 514658 549586 514894
rect 549822 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 9266 514574
rect 9502 514338 9586 514574
rect 9822 514338 45266 514574
rect 45502 514338 45586 514574
rect 45822 514338 81266 514574
rect 81502 514338 81586 514574
rect 81822 514338 117266 514574
rect 117502 514338 117586 514574
rect 117822 514338 153266 514574
rect 153502 514338 153586 514574
rect 153822 514338 189266 514574
rect 189502 514338 189586 514574
rect 189822 514338 225266 514574
rect 225502 514338 225586 514574
rect 225822 514338 261266 514574
rect 261502 514338 261586 514574
rect 261822 514338 297266 514574
rect 297502 514338 297586 514574
rect 297822 514338 333266 514574
rect 333502 514338 333586 514574
rect 333822 514338 369266 514574
rect 369502 514338 369586 514574
rect 369822 514338 405266 514574
rect 405502 514338 405586 514574
rect 405822 514338 441266 514574
rect 441502 514338 441586 514574
rect 441822 514338 477266 514574
rect 477502 514338 477586 514574
rect 477822 514338 513266 514574
rect 513502 514338 513586 514574
rect 513822 514338 549266 514574
rect 549502 514338 549586 514574
rect 549822 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 5546 511174
rect 5782 510938 5866 511174
rect 6102 510938 41546 511174
rect 41782 510938 41866 511174
rect 42102 510938 77546 511174
rect 77782 510938 77866 511174
rect 78102 510938 113546 511174
rect 113782 510938 113866 511174
rect 114102 510938 149546 511174
rect 149782 510938 149866 511174
rect 150102 510938 185546 511174
rect 185782 510938 185866 511174
rect 186102 510938 221546 511174
rect 221782 510938 221866 511174
rect 222102 510938 257546 511174
rect 257782 510938 257866 511174
rect 258102 510938 293546 511174
rect 293782 510938 293866 511174
rect 294102 510938 329546 511174
rect 329782 510938 329866 511174
rect 330102 510938 365546 511174
rect 365782 510938 365866 511174
rect 366102 510938 401546 511174
rect 401782 510938 401866 511174
rect 402102 510938 437546 511174
rect 437782 510938 437866 511174
rect 438102 510938 473546 511174
rect 473782 510938 473866 511174
rect 474102 510938 509546 511174
rect 509782 510938 509866 511174
rect 510102 510938 545546 511174
rect 545782 510938 545866 511174
rect 546102 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 5546 510854
rect 5782 510618 5866 510854
rect 6102 510618 41546 510854
rect 41782 510618 41866 510854
rect 42102 510618 77546 510854
rect 77782 510618 77866 510854
rect 78102 510618 113546 510854
rect 113782 510618 113866 510854
rect 114102 510618 149546 510854
rect 149782 510618 149866 510854
rect 150102 510618 185546 510854
rect 185782 510618 185866 510854
rect 186102 510618 221546 510854
rect 221782 510618 221866 510854
rect 222102 510618 257546 510854
rect 257782 510618 257866 510854
rect 258102 510618 293546 510854
rect 293782 510618 293866 510854
rect 294102 510618 329546 510854
rect 329782 510618 329866 510854
rect 330102 510618 365546 510854
rect 365782 510618 365866 510854
rect 366102 510618 401546 510854
rect 401782 510618 401866 510854
rect 402102 510618 437546 510854
rect 437782 510618 437866 510854
rect 438102 510618 473546 510854
rect 473782 510618 473866 510854
rect 474102 510618 509546 510854
rect 509782 510618 509866 510854
rect 510102 510618 545546 510854
rect 545782 510618 545866 510854
rect 546102 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 1826 507454
rect 2062 507218 2146 507454
rect 2382 507218 37826 507454
rect 38062 507218 38146 507454
rect 38382 507218 73826 507454
rect 74062 507218 74146 507454
rect 74382 507218 109826 507454
rect 110062 507218 110146 507454
rect 110382 507218 145826 507454
rect 146062 507218 146146 507454
rect 146382 507218 181826 507454
rect 182062 507218 182146 507454
rect 182382 507218 217826 507454
rect 218062 507218 218146 507454
rect 218382 507218 253826 507454
rect 254062 507218 254146 507454
rect 254382 507218 289826 507454
rect 290062 507218 290146 507454
rect 290382 507218 325826 507454
rect 326062 507218 326146 507454
rect 326382 507218 361826 507454
rect 362062 507218 362146 507454
rect 362382 507218 397826 507454
rect 398062 507218 398146 507454
rect 398382 507218 433826 507454
rect 434062 507218 434146 507454
rect 434382 507218 469826 507454
rect 470062 507218 470146 507454
rect 470382 507218 505826 507454
rect 506062 507218 506146 507454
rect 506382 507218 541826 507454
rect 542062 507218 542146 507454
rect 542382 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 1826 507134
rect 2062 506898 2146 507134
rect 2382 506898 37826 507134
rect 38062 506898 38146 507134
rect 38382 506898 73826 507134
rect 74062 506898 74146 507134
rect 74382 506898 109826 507134
rect 110062 506898 110146 507134
rect 110382 506898 145826 507134
rect 146062 506898 146146 507134
rect 146382 506898 181826 507134
rect 182062 506898 182146 507134
rect 182382 506898 217826 507134
rect 218062 506898 218146 507134
rect 218382 506898 253826 507134
rect 254062 506898 254146 507134
rect 254382 506898 289826 507134
rect 290062 506898 290146 507134
rect 290382 506898 325826 507134
rect 326062 506898 326146 507134
rect 326382 506898 361826 507134
rect 362062 506898 362146 507134
rect 362382 506898 397826 507134
rect 398062 506898 398146 507134
rect 398382 506898 433826 507134
rect 434062 506898 434146 507134
rect 434382 506898 469826 507134
rect 470062 506898 470146 507134
rect 470382 506898 505826 507134
rect 506062 506898 506146 507134
rect 506382 506898 541826 507134
rect 542062 506898 542146 507134
rect 542382 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 30986 500614
rect 31222 500378 31306 500614
rect 31542 500378 66986 500614
rect 67222 500378 67306 500614
rect 67542 500378 102986 500614
rect 103222 500378 103306 500614
rect 103542 500378 138986 500614
rect 139222 500378 139306 500614
rect 139542 500378 174986 500614
rect 175222 500378 175306 500614
rect 175542 500378 210986 500614
rect 211222 500378 211306 500614
rect 211542 500378 246986 500614
rect 247222 500378 247306 500614
rect 247542 500378 282986 500614
rect 283222 500378 283306 500614
rect 283542 500378 318986 500614
rect 319222 500378 319306 500614
rect 319542 500378 354986 500614
rect 355222 500378 355306 500614
rect 355542 500378 390986 500614
rect 391222 500378 391306 500614
rect 391542 500378 426986 500614
rect 427222 500378 427306 500614
rect 427542 500378 462986 500614
rect 463222 500378 463306 500614
rect 463542 500378 498986 500614
rect 499222 500378 499306 500614
rect 499542 500378 534986 500614
rect 535222 500378 535306 500614
rect 535542 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 30986 500294
rect 31222 500058 31306 500294
rect 31542 500058 66986 500294
rect 67222 500058 67306 500294
rect 67542 500058 102986 500294
rect 103222 500058 103306 500294
rect 103542 500058 138986 500294
rect 139222 500058 139306 500294
rect 139542 500058 174986 500294
rect 175222 500058 175306 500294
rect 175542 500058 210986 500294
rect 211222 500058 211306 500294
rect 211542 500058 246986 500294
rect 247222 500058 247306 500294
rect 247542 500058 282986 500294
rect 283222 500058 283306 500294
rect 283542 500058 318986 500294
rect 319222 500058 319306 500294
rect 319542 500058 354986 500294
rect 355222 500058 355306 500294
rect 355542 500058 390986 500294
rect 391222 500058 391306 500294
rect 391542 500058 426986 500294
rect 427222 500058 427306 500294
rect 427542 500058 462986 500294
rect 463222 500058 463306 500294
rect 463542 500058 498986 500294
rect 499222 500058 499306 500294
rect 499542 500058 534986 500294
rect 535222 500058 535306 500294
rect 535542 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 27266 496894
rect 27502 496658 27586 496894
rect 27822 496658 63266 496894
rect 63502 496658 63586 496894
rect 63822 496658 99266 496894
rect 99502 496658 99586 496894
rect 99822 496658 135266 496894
rect 135502 496658 135586 496894
rect 135822 496658 171266 496894
rect 171502 496658 171586 496894
rect 171822 496658 207266 496894
rect 207502 496658 207586 496894
rect 207822 496658 243266 496894
rect 243502 496658 243586 496894
rect 243822 496658 279266 496894
rect 279502 496658 279586 496894
rect 279822 496658 315266 496894
rect 315502 496658 315586 496894
rect 315822 496658 351266 496894
rect 351502 496658 351586 496894
rect 351822 496658 387266 496894
rect 387502 496658 387586 496894
rect 387822 496658 423266 496894
rect 423502 496658 423586 496894
rect 423822 496658 459266 496894
rect 459502 496658 459586 496894
rect 459822 496658 495266 496894
rect 495502 496658 495586 496894
rect 495822 496658 531266 496894
rect 531502 496658 531586 496894
rect 531822 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 27266 496574
rect 27502 496338 27586 496574
rect 27822 496338 63266 496574
rect 63502 496338 63586 496574
rect 63822 496338 99266 496574
rect 99502 496338 99586 496574
rect 99822 496338 135266 496574
rect 135502 496338 135586 496574
rect 135822 496338 171266 496574
rect 171502 496338 171586 496574
rect 171822 496338 207266 496574
rect 207502 496338 207586 496574
rect 207822 496338 243266 496574
rect 243502 496338 243586 496574
rect 243822 496338 279266 496574
rect 279502 496338 279586 496574
rect 279822 496338 315266 496574
rect 315502 496338 315586 496574
rect 315822 496338 351266 496574
rect 351502 496338 351586 496574
rect 351822 496338 387266 496574
rect 387502 496338 387586 496574
rect 387822 496338 423266 496574
rect 423502 496338 423586 496574
rect 423822 496338 459266 496574
rect 459502 496338 459586 496574
rect 459822 496338 495266 496574
rect 495502 496338 495586 496574
rect 495822 496338 531266 496574
rect 531502 496338 531586 496574
rect 531822 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 23546 493174
rect 23782 492938 23866 493174
rect 24102 492938 59546 493174
rect 59782 492938 59866 493174
rect 60102 492938 95546 493174
rect 95782 492938 95866 493174
rect 96102 492938 131546 493174
rect 131782 492938 131866 493174
rect 132102 492938 167546 493174
rect 167782 492938 167866 493174
rect 168102 492938 203546 493174
rect 203782 492938 203866 493174
rect 204102 492938 239546 493174
rect 239782 492938 239866 493174
rect 240102 492938 275546 493174
rect 275782 492938 275866 493174
rect 276102 492938 311546 493174
rect 311782 492938 311866 493174
rect 312102 492938 347546 493174
rect 347782 492938 347866 493174
rect 348102 492938 383546 493174
rect 383782 492938 383866 493174
rect 384102 492938 419546 493174
rect 419782 492938 419866 493174
rect 420102 492938 455546 493174
rect 455782 492938 455866 493174
rect 456102 492938 491546 493174
rect 491782 492938 491866 493174
rect 492102 492938 527546 493174
rect 527782 492938 527866 493174
rect 528102 492938 563546 493174
rect 563782 492938 563866 493174
rect 564102 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 23546 492854
rect 23782 492618 23866 492854
rect 24102 492618 59546 492854
rect 59782 492618 59866 492854
rect 60102 492618 95546 492854
rect 95782 492618 95866 492854
rect 96102 492618 131546 492854
rect 131782 492618 131866 492854
rect 132102 492618 167546 492854
rect 167782 492618 167866 492854
rect 168102 492618 203546 492854
rect 203782 492618 203866 492854
rect 204102 492618 239546 492854
rect 239782 492618 239866 492854
rect 240102 492618 275546 492854
rect 275782 492618 275866 492854
rect 276102 492618 311546 492854
rect 311782 492618 311866 492854
rect 312102 492618 347546 492854
rect 347782 492618 347866 492854
rect 348102 492618 383546 492854
rect 383782 492618 383866 492854
rect 384102 492618 419546 492854
rect 419782 492618 419866 492854
rect 420102 492618 455546 492854
rect 455782 492618 455866 492854
rect 456102 492618 491546 492854
rect 491782 492618 491866 492854
rect 492102 492618 527546 492854
rect 527782 492618 527866 492854
rect 528102 492618 563546 492854
rect 563782 492618 563866 492854
rect 564102 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 19826 489454
rect 20062 489218 20146 489454
rect 20382 489218 55826 489454
rect 56062 489218 56146 489454
rect 56382 489218 91826 489454
rect 92062 489218 92146 489454
rect 92382 489218 127826 489454
rect 128062 489218 128146 489454
rect 128382 489218 163826 489454
rect 164062 489218 164146 489454
rect 164382 489218 199826 489454
rect 200062 489218 200146 489454
rect 200382 489218 235826 489454
rect 236062 489218 236146 489454
rect 236382 489218 271826 489454
rect 272062 489218 272146 489454
rect 272382 489218 307826 489454
rect 308062 489218 308146 489454
rect 308382 489218 343826 489454
rect 344062 489218 344146 489454
rect 344382 489218 379826 489454
rect 380062 489218 380146 489454
rect 380382 489218 415826 489454
rect 416062 489218 416146 489454
rect 416382 489218 451826 489454
rect 452062 489218 452146 489454
rect 452382 489218 487826 489454
rect 488062 489218 488146 489454
rect 488382 489218 523826 489454
rect 524062 489218 524146 489454
rect 524382 489218 559826 489454
rect 560062 489218 560146 489454
rect 560382 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 19826 489134
rect 20062 488898 20146 489134
rect 20382 488898 55826 489134
rect 56062 488898 56146 489134
rect 56382 488898 91826 489134
rect 92062 488898 92146 489134
rect 92382 488898 127826 489134
rect 128062 488898 128146 489134
rect 128382 488898 163826 489134
rect 164062 488898 164146 489134
rect 164382 488898 199826 489134
rect 200062 488898 200146 489134
rect 200382 488898 235826 489134
rect 236062 488898 236146 489134
rect 236382 488898 271826 489134
rect 272062 488898 272146 489134
rect 272382 488898 307826 489134
rect 308062 488898 308146 489134
rect 308382 488898 343826 489134
rect 344062 488898 344146 489134
rect 344382 488898 379826 489134
rect 380062 488898 380146 489134
rect 380382 488898 415826 489134
rect 416062 488898 416146 489134
rect 416382 488898 451826 489134
rect 452062 488898 452146 489134
rect 452382 488898 487826 489134
rect 488062 488898 488146 489134
rect 488382 488898 523826 489134
rect 524062 488898 524146 489134
rect 524382 488898 559826 489134
rect 560062 488898 560146 489134
rect 560382 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 12986 482614
rect 13222 482378 13306 482614
rect 13542 482378 48986 482614
rect 49222 482378 49306 482614
rect 49542 482378 372986 482614
rect 373222 482378 373306 482614
rect 373542 482378 408986 482614
rect 409222 482378 409306 482614
rect 409542 482378 444986 482614
rect 445222 482378 445306 482614
rect 445542 482378 480986 482614
rect 481222 482378 481306 482614
rect 481542 482378 516986 482614
rect 517222 482378 517306 482614
rect 517542 482378 552986 482614
rect 553222 482378 553306 482614
rect 553542 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 12986 482294
rect 13222 482058 13306 482294
rect 13542 482058 48986 482294
rect 49222 482058 49306 482294
rect 49542 482058 372986 482294
rect 373222 482058 373306 482294
rect 373542 482058 408986 482294
rect 409222 482058 409306 482294
rect 409542 482058 444986 482294
rect 445222 482058 445306 482294
rect 445542 482058 480986 482294
rect 481222 482058 481306 482294
rect 481542 482058 516986 482294
rect 517222 482058 517306 482294
rect 517542 482058 552986 482294
rect 553222 482058 553306 482294
rect 553542 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 9266 478894
rect 9502 478658 9586 478894
rect 9822 478658 45266 478894
rect 45502 478658 45586 478894
rect 45822 478658 369266 478894
rect 369502 478658 369586 478894
rect 369822 478658 405266 478894
rect 405502 478658 405586 478894
rect 405822 478658 441266 478894
rect 441502 478658 441586 478894
rect 441822 478658 477266 478894
rect 477502 478658 477586 478894
rect 477822 478658 513266 478894
rect 513502 478658 513586 478894
rect 513822 478658 549266 478894
rect 549502 478658 549586 478894
rect 549822 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 9266 478574
rect 9502 478338 9586 478574
rect 9822 478338 45266 478574
rect 45502 478338 45586 478574
rect 45822 478338 369266 478574
rect 369502 478338 369586 478574
rect 369822 478338 405266 478574
rect 405502 478338 405586 478574
rect 405822 478338 441266 478574
rect 441502 478338 441586 478574
rect 441822 478338 477266 478574
rect 477502 478338 477586 478574
rect 477822 478338 513266 478574
rect 513502 478338 513586 478574
rect 513822 478338 549266 478574
rect 549502 478338 549586 478574
rect 549822 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 5546 475174
rect 5782 474938 5866 475174
rect 6102 474938 41546 475174
rect 41782 474938 41866 475174
rect 42102 474938 365546 475174
rect 365782 474938 365866 475174
rect 366102 474938 401546 475174
rect 401782 474938 401866 475174
rect 402102 474938 437546 475174
rect 437782 474938 437866 475174
rect 438102 474938 473546 475174
rect 473782 474938 473866 475174
rect 474102 474938 509546 475174
rect 509782 474938 509866 475174
rect 510102 474938 545546 475174
rect 545782 474938 545866 475174
rect 546102 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 5546 474854
rect 5782 474618 5866 474854
rect 6102 474618 41546 474854
rect 41782 474618 41866 474854
rect 42102 474618 365546 474854
rect 365782 474618 365866 474854
rect 366102 474618 401546 474854
rect 401782 474618 401866 474854
rect 402102 474618 437546 474854
rect 437782 474618 437866 474854
rect 438102 474618 473546 474854
rect 473782 474618 473866 474854
rect 474102 474618 509546 474854
rect 509782 474618 509866 474854
rect 510102 474618 545546 474854
rect 545782 474618 545866 474854
rect 546102 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 1826 471454
rect 2062 471218 2146 471454
rect 2382 471218 37826 471454
rect 38062 471218 38146 471454
rect 38382 471218 61008 471454
rect 61244 471218 195376 471454
rect 195612 471218 221008 471454
rect 221244 471218 355376 471454
rect 355612 471218 361826 471454
rect 362062 471218 362146 471454
rect 362382 471218 397826 471454
rect 398062 471218 398146 471454
rect 398382 471218 433826 471454
rect 434062 471218 434146 471454
rect 434382 471218 469826 471454
rect 470062 471218 470146 471454
rect 470382 471218 505826 471454
rect 506062 471218 506146 471454
rect 506382 471218 541826 471454
rect 542062 471218 542146 471454
rect 542382 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 1826 471134
rect 2062 470898 2146 471134
rect 2382 470898 37826 471134
rect 38062 470898 38146 471134
rect 38382 470898 61008 471134
rect 61244 470898 195376 471134
rect 195612 470898 221008 471134
rect 221244 470898 355376 471134
rect 355612 470898 361826 471134
rect 362062 470898 362146 471134
rect 362382 470898 397826 471134
rect 398062 470898 398146 471134
rect 398382 470898 433826 471134
rect 434062 470898 434146 471134
rect 434382 470898 469826 471134
rect 470062 470898 470146 471134
rect 470382 470898 505826 471134
rect 506062 470898 506146 471134
rect 506382 470898 541826 471134
rect 542062 470898 542146 471134
rect 542382 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 30986 464614
rect 31222 464378 31306 464614
rect 31542 464378 210986 464614
rect 211222 464378 211306 464614
rect 211542 464378 390986 464614
rect 391222 464378 391306 464614
rect 391542 464378 426986 464614
rect 427222 464378 427306 464614
rect 427542 464378 462986 464614
rect 463222 464378 463306 464614
rect 463542 464378 498986 464614
rect 499222 464378 499306 464614
rect 499542 464378 534986 464614
rect 535222 464378 535306 464614
rect 535542 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 30986 464294
rect 31222 464058 31306 464294
rect 31542 464058 210986 464294
rect 211222 464058 211306 464294
rect 211542 464058 390986 464294
rect 391222 464058 391306 464294
rect 391542 464058 426986 464294
rect 427222 464058 427306 464294
rect 427542 464058 462986 464294
rect 463222 464058 463306 464294
rect 463542 464058 498986 464294
rect 499222 464058 499306 464294
rect 499542 464058 534986 464294
rect 535222 464058 535306 464294
rect 535542 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 27266 460894
rect 27502 460658 27586 460894
rect 27822 460658 207266 460894
rect 207502 460658 207586 460894
rect 207822 460658 387266 460894
rect 387502 460658 387586 460894
rect 387822 460658 423266 460894
rect 423502 460658 423586 460894
rect 423822 460658 459266 460894
rect 459502 460658 459586 460894
rect 459822 460658 495266 460894
rect 495502 460658 495586 460894
rect 495822 460658 531266 460894
rect 531502 460658 531586 460894
rect 531822 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 27266 460574
rect 27502 460338 27586 460574
rect 27822 460338 207266 460574
rect 207502 460338 207586 460574
rect 207822 460338 387266 460574
rect 387502 460338 387586 460574
rect 387822 460338 423266 460574
rect 423502 460338 423586 460574
rect 423822 460338 459266 460574
rect 459502 460338 459586 460574
rect 459822 460338 495266 460574
rect 495502 460338 495586 460574
rect 495822 460338 531266 460574
rect 531502 460338 531586 460574
rect 531822 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 23546 457174
rect 23782 456938 23866 457174
rect 24102 456938 203546 457174
rect 203782 456938 203866 457174
rect 204102 456938 383546 457174
rect 383782 456938 383866 457174
rect 384102 456938 419546 457174
rect 419782 456938 419866 457174
rect 420102 456938 455546 457174
rect 455782 456938 455866 457174
rect 456102 456938 491546 457174
rect 491782 456938 491866 457174
rect 492102 456938 527546 457174
rect 527782 456938 527866 457174
rect 528102 456938 563546 457174
rect 563782 456938 563866 457174
rect 564102 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 23546 456854
rect 23782 456618 23866 456854
rect 24102 456618 203546 456854
rect 203782 456618 203866 456854
rect 204102 456618 383546 456854
rect 383782 456618 383866 456854
rect 384102 456618 419546 456854
rect 419782 456618 419866 456854
rect 420102 456618 455546 456854
rect 455782 456618 455866 456854
rect 456102 456618 491546 456854
rect 491782 456618 491866 456854
rect 492102 456618 527546 456854
rect 527782 456618 527866 456854
rect 528102 456618 563546 456854
rect 563782 456618 563866 456854
rect 564102 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 19826 453454
rect 20062 453218 20146 453454
rect 20382 453218 55826 453454
rect 56062 453218 56146 453454
rect 56382 453218 60328 453454
rect 60564 453218 196056 453454
rect 196292 453218 199826 453454
rect 200062 453218 200146 453454
rect 200382 453218 220328 453454
rect 220564 453218 356056 453454
rect 356292 453218 379826 453454
rect 380062 453218 380146 453454
rect 380382 453218 415826 453454
rect 416062 453218 416146 453454
rect 416382 453218 451826 453454
rect 452062 453218 452146 453454
rect 452382 453218 487826 453454
rect 488062 453218 488146 453454
rect 488382 453218 523826 453454
rect 524062 453218 524146 453454
rect 524382 453218 559826 453454
rect 560062 453218 560146 453454
rect 560382 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 19826 453134
rect 20062 452898 20146 453134
rect 20382 452898 55826 453134
rect 56062 452898 56146 453134
rect 56382 452898 60328 453134
rect 60564 452898 196056 453134
rect 196292 452898 199826 453134
rect 200062 452898 200146 453134
rect 200382 452898 220328 453134
rect 220564 452898 356056 453134
rect 356292 452898 379826 453134
rect 380062 452898 380146 453134
rect 380382 452898 415826 453134
rect 416062 452898 416146 453134
rect 416382 452898 451826 453134
rect 452062 452898 452146 453134
rect 452382 452898 487826 453134
rect 488062 452898 488146 453134
rect 488382 452898 523826 453134
rect 524062 452898 524146 453134
rect 524382 452898 559826 453134
rect 560062 452898 560146 453134
rect 560382 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 12986 446614
rect 13222 446378 13306 446614
rect 13542 446378 48986 446614
rect 49222 446378 49306 446614
rect 49542 446378 372986 446614
rect 373222 446378 373306 446614
rect 373542 446378 408986 446614
rect 409222 446378 409306 446614
rect 409542 446378 444986 446614
rect 445222 446378 445306 446614
rect 445542 446378 480986 446614
rect 481222 446378 481306 446614
rect 481542 446378 516986 446614
rect 517222 446378 517306 446614
rect 517542 446378 552986 446614
rect 553222 446378 553306 446614
rect 553542 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 12986 446294
rect 13222 446058 13306 446294
rect 13542 446058 48986 446294
rect 49222 446058 49306 446294
rect 49542 446058 372986 446294
rect 373222 446058 373306 446294
rect 373542 446058 408986 446294
rect 409222 446058 409306 446294
rect 409542 446058 444986 446294
rect 445222 446058 445306 446294
rect 445542 446058 480986 446294
rect 481222 446058 481306 446294
rect 481542 446058 516986 446294
rect 517222 446058 517306 446294
rect 517542 446058 552986 446294
rect 553222 446058 553306 446294
rect 553542 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 9266 442894
rect 9502 442658 9586 442894
rect 9822 442658 45266 442894
rect 45502 442658 45586 442894
rect 45822 442658 369266 442894
rect 369502 442658 369586 442894
rect 369822 442658 405266 442894
rect 405502 442658 405586 442894
rect 405822 442658 441266 442894
rect 441502 442658 441586 442894
rect 441822 442658 477266 442894
rect 477502 442658 477586 442894
rect 477822 442658 513266 442894
rect 513502 442658 513586 442894
rect 513822 442658 549266 442894
rect 549502 442658 549586 442894
rect 549822 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 9266 442574
rect 9502 442338 9586 442574
rect 9822 442338 45266 442574
rect 45502 442338 45586 442574
rect 45822 442338 369266 442574
rect 369502 442338 369586 442574
rect 369822 442338 405266 442574
rect 405502 442338 405586 442574
rect 405822 442338 441266 442574
rect 441502 442338 441586 442574
rect 441822 442338 477266 442574
rect 477502 442338 477586 442574
rect 477822 442338 513266 442574
rect 513502 442338 513586 442574
rect 513822 442338 549266 442574
rect 549502 442338 549586 442574
rect 549822 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 5546 439174
rect 5782 438938 5866 439174
rect 6102 438938 41546 439174
rect 41782 438938 41866 439174
rect 42102 438938 365546 439174
rect 365782 438938 365866 439174
rect 366102 438938 401546 439174
rect 401782 438938 401866 439174
rect 402102 438938 437546 439174
rect 437782 438938 437866 439174
rect 438102 438938 473546 439174
rect 473782 438938 473866 439174
rect 474102 438938 509546 439174
rect 509782 438938 509866 439174
rect 510102 438938 545546 439174
rect 545782 438938 545866 439174
rect 546102 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 5546 438854
rect 5782 438618 5866 438854
rect 6102 438618 41546 438854
rect 41782 438618 41866 438854
rect 42102 438618 365546 438854
rect 365782 438618 365866 438854
rect 366102 438618 401546 438854
rect 401782 438618 401866 438854
rect 402102 438618 437546 438854
rect 437782 438618 437866 438854
rect 438102 438618 473546 438854
rect 473782 438618 473866 438854
rect 474102 438618 509546 438854
rect 509782 438618 509866 438854
rect 510102 438618 545546 438854
rect 545782 438618 545866 438854
rect 546102 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 1826 435454
rect 2062 435218 2146 435454
rect 2382 435218 37826 435454
rect 38062 435218 38146 435454
rect 38382 435218 61008 435454
rect 61244 435218 195376 435454
rect 195612 435218 221008 435454
rect 221244 435218 355376 435454
rect 355612 435218 361826 435454
rect 362062 435218 362146 435454
rect 362382 435218 397826 435454
rect 398062 435218 398146 435454
rect 398382 435218 433826 435454
rect 434062 435218 434146 435454
rect 434382 435218 469826 435454
rect 470062 435218 470146 435454
rect 470382 435218 505826 435454
rect 506062 435218 506146 435454
rect 506382 435218 541826 435454
rect 542062 435218 542146 435454
rect 542382 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 1826 435134
rect 2062 434898 2146 435134
rect 2382 434898 37826 435134
rect 38062 434898 38146 435134
rect 38382 434898 61008 435134
rect 61244 434898 195376 435134
rect 195612 434898 221008 435134
rect 221244 434898 355376 435134
rect 355612 434898 361826 435134
rect 362062 434898 362146 435134
rect 362382 434898 397826 435134
rect 398062 434898 398146 435134
rect 398382 434898 433826 435134
rect 434062 434898 434146 435134
rect 434382 434898 469826 435134
rect 470062 434898 470146 435134
rect 470382 434898 505826 435134
rect 506062 434898 506146 435134
rect 506382 434898 541826 435134
rect 542062 434898 542146 435134
rect 542382 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 30986 428614
rect 31222 428378 31306 428614
rect 31542 428378 210986 428614
rect 211222 428378 211306 428614
rect 211542 428378 390986 428614
rect 391222 428378 391306 428614
rect 391542 428378 426986 428614
rect 427222 428378 427306 428614
rect 427542 428378 462986 428614
rect 463222 428378 463306 428614
rect 463542 428378 498986 428614
rect 499222 428378 499306 428614
rect 499542 428378 534986 428614
rect 535222 428378 535306 428614
rect 535542 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 30986 428294
rect 31222 428058 31306 428294
rect 31542 428058 210986 428294
rect 211222 428058 211306 428294
rect 211542 428058 390986 428294
rect 391222 428058 391306 428294
rect 391542 428058 426986 428294
rect 427222 428058 427306 428294
rect 427542 428058 462986 428294
rect 463222 428058 463306 428294
rect 463542 428058 498986 428294
rect 499222 428058 499306 428294
rect 499542 428058 534986 428294
rect 535222 428058 535306 428294
rect 535542 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 27266 424894
rect 27502 424658 27586 424894
rect 27822 424658 207266 424894
rect 207502 424658 207586 424894
rect 207822 424658 387266 424894
rect 387502 424658 387586 424894
rect 387822 424658 423266 424894
rect 423502 424658 423586 424894
rect 423822 424658 459266 424894
rect 459502 424658 459586 424894
rect 459822 424658 495266 424894
rect 495502 424658 495586 424894
rect 495822 424658 531266 424894
rect 531502 424658 531586 424894
rect 531822 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 27266 424574
rect 27502 424338 27586 424574
rect 27822 424338 207266 424574
rect 207502 424338 207586 424574
rect 207822 424338 387266 424574
rect 387502 424338 387586 424574
rect 387822 424338 423266 424574
rect 423502 424338 423586 424574
rect 423822 424338 459266 424574
rect 459502 424338 459586 424574
rect 459822 424338 495266 424574
rect 495502 424338 495586 424574
rect 495822 424338 531266 424574
rect 531502 424338 531586 424574
rect 531822 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 23546 421174
rect 23782 420938 23866 421174
rect 24102 420938 203546 421174
rect 203782 420938 203866 421174
rect 204102 420938 383546 421174
rect 383782 420938 383866 421174
rect 384102 420938 419546 421174
rect 419782 420938 419866 421174
rect 420102 420938 455546 421174
rect 455782 420938 455866 421174
rect 456102 420938 491546 421174
rect 491782 420938 491866 421174
rect 492102 420938 527546 421174
rect 527782 420938 527866 421174
rect 528102 420938 563546 421174
rect 563782 420938 563866 421174
rect 564102 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 23546 420854
rect 23782 420618 23866 420854
rect 24102 420618 203546 420854
rect 203782 420618 203866 420854
rect 204102 420618 383546 420854
rect 383782 420618 383866 420854
rect 384102 420618 419546 420854
rect 419782 420618 419866 420854
rect 420102 420618 455546 420854
rect 455782 420618 455866 420854
rect 456102 420618 491546 420854
rect 491782 420618 491866 420854
rect 492102 420618 527546 420854
rect 527782 420618 527866 420854
rect 528102 420618 563546 420854
rect 563782 420618 563866 420854
rect 564102 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 19826 417454
rect 20062 417218 20146 417454
rect 20382 417218 55826 417454
rect 56062 417218 56146 417454
rect 56382 417218 60328 417454
rect 60564 417218 196056 417454
rect 196292 417218 199826 417454
rect 200062 417218 200146 417454
rect 200382 417218 220328 417454
rect 220564 417218 356056 417454
rect 356292 417218 379826 417454
rect 380062 417218 380146 417454
rect 380382 417218 415826 417454
rect 416062 417218 416146 417454
rect 416382 417218 451826 417454
rect 452062 417218 452146 417454
rect 452382 417218 487826 417454
rect 488062 417218 488146 417454
rect 488382 417218 523826 417454
rect 524062 417218 524146 417454
rect 524382 417218 559826 417454
rect 560062 417218 560146 417454
rect 560382 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 19826 417134
rect 20062 416898 20146 417134
rect 20382 416898 55826 417134
rect 56062 416898 56146 417134
rect 56382 416898 60328 417134
rect 60564 416898 196056 417134
rect 196292 416898 199826 417134
rect 200062 416898 200146 417134
rect 200382 416898 220328 417134
rect 220564 416898 356056 417134
rect 356292 416898 379826 417134
rect 380062 416898 380146 417134
rect 380382 416898 415826 417134
rect 416062 416898 416146 417134
rect 416382 416898 451826 417134
rect 452062 416898 452146 417134
rect 452382 416898 487826 417134
rect 488062 416898 488146 417134
rect 488382 416898 523826 417134
rect 524062 416898 524146 417134
rect 524382 416898 559826 417134
rect 560062 416898 560146 417134
rect 560382 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 12986 410614
rect 13222 410378 13306 410614
rect 13542 410378 48986 410614
rect 49222 410378 49306 410614
rect 49542 410378 372986 410614
rect 373222 410378 373306 410614
rect 373542 410378 408986 410614
rect 409222 410378 409306 410614
rect 409542 410378 444986 410614
rect 445222 410378 445306 410614
rect 445542 410378 480986 410614
rect 481222 410378 481306 410614
rect 481542 410378 516986 410614
rect 517222 410378 517306 410614
rect 517542 410378 552986 410614
rect 553222 410378 553306 410614
rect 553542 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 12986 410294
rect 13222 410058 13306 410294
rect 13542 410058 48986 410294
rect 49222 410058 49306 410294
rect 49542 410058 372986 410294
rect 373222 410058 373306 410294
rect 373542 410058 408986 410294
rect 409222 410058 409306 410294
rect 409542 410058 444986 410294
rect 445222 410058 445306 410294
rect 445542 410058 480986 410294
rect 481222 410058 481306 410294
rect 481542 410058 516986 410294
rect 517222 410058 517306 410294
rect 517542 410058 552986 410294
rect 553222 410058 553306 410294
rect 553542 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 9266 406894
rect 9502 406658 9586 406894
rect 9822 406658 45266 406894
rect 45502 406658 45586 406894
rect 45822 406658 369266 406894
rect 369502 406658 369586 406894
rect 369822 406658 405266 406894
rect 405502 406658 405586 406894
rect 405822 406658 441266 406894
rect 441502 406658 441586 406894
rect 441822 406658 477266 406894
rect 477502 406658 477586 406894
rect 477822 406658 513266 406894
rect 513502 406658 513586 406894
rect 513822 406658 549266 406894
rect 549502 406658 549586 406894
rect 549822 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 9266 406574
rect 9502 406338 9586 406574
rect 9822 406338 45266 406574
rect 45502 406338 45586 406574
rect 45822 406338 369266 406574
rect 369502 406338 369586 406574
rect 369822 406338 405266 406574
rect 405502 406338 405586 406574
rect 405822 406338 441266 406574
rect 441502 406338 441586 406574
rect 441822 406338 477266 406574
rect 477502 406338 477586 406574
rect 477822 406338 513266 406574
rect 513502 406338 513586 406574
rect 513822 406338 549266 406574
rect 549502 406338 549586 406574
rect 549822 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 5546 403174
rect 5782 402938 5866 403174
rect 6102 402938 41546 403174
rect 41782 402938 41866 403174
rect 42102 402938 365546 403174
rect 365782 402938 365866 403174
rect 366102 402938 401546 403174
rect 401782 402938 401866 403174
rect 402102 402938 437546 403174
rect 437782 402938 437866 403174
rect 438102 402938 473546 403174
rect 473782 402938 473866 403174
rect 474102 402938 509546 403174
rect 509782 402938 509866 403174
rect 510102 402938 545546 403174
rect 545782 402938 545866 403174
rect 546102 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 5546 402854
rect 5782 402618 5866 402854
rect 6102 402618 41546 402854
rect 41782 402618 41866 402854
rect 42102 402618 365546 402854
rect 365782 402618 365866 402854
rect 366102 402618 401546 402854
rect 401782 402618 401866 402854
rect 402102 402618 437546 402854
rect 437782 402618 437866 402854
rect 438102 402618 473546 402854
rect 473782 402618 473866 402854
rect 474102 402618 509546 402854
rect 509782 402618 509866 402854
rect 510102 402618 545546 402854
rect 545782 402618 545866 402854
rect 546102 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 1826 399454
rect 2062 399218 2146 399454
rect 2382 399218 37826 399454
rect 38062 399218 38146 399454
rect 38382 399218 361826 399454
rect 362062 399218 362146 399454
rect 362382 399218 397826 399454
rect 398062 399218 398146 399454
rect 398382 399218 433826 399454
rect 434062 399218 434146 399454
rect 434382 399218 469826 399454
rect 470062 399218 470146 399454
rect 470382 399218 505826 399454
rect 506062 399218 506146 399454
rect 506382 399218 541826 399454
rect 542062 399218 542146 399454
rect 542382 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 1826 399134
rect 2062 398898 2146 399134
rect 2382 398898 37826 399134
rect 38062 398898 38146 399134
rect 38382 398898 361826 399134
rect 362062 398898 362146 399134
rect 362382 398898 397826 399134
rect 398062 398898 398146 399134
rect 398382 398898 433826 399134
rect 434062 398898 434146 399134
rect 434382 398898 469826 399134
rect 470062 398898 470146 399134
rect 470382 398898 505826 399134
rect 506062 398898 506146 399134
rect 506382 398898 541826 399134
rect 542062 398898 542146 399134
rect 542382 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 30986 392614
rect 31222 392378 31306 392614
rect 31542 392378 66986 392614
rect 67222 392378 67306 392614
rect 67542 392378 102986 392614
rect 103222 392378 103306 392614
rect 103542 392378 138986 392614
rect 139222 392378 139306 392614
rect 139542 392378 174986 392614
rect 175222 392378 175306 392614
rect 175542 392378 210986 392614
rect 211222 392378 211306 392614
rect 211542 392378 246986 392614
rect 247222 392378 247306 392614
rect 247542 392378 282986 392614
rect 283222 392378 283306 392614
rect 283542 392378 318986 392614
rect 319222 392378 319306 392614
rect 319542 392378 354986 392614
rect 355222 392378 355306 392614
rect 355542 392378 390986 392614
rect 391222 392378 391306 392614
rect 391542 392378 426986 392614
rect 427222 392378 427306 392614
rect 427542 392378 462986 392614
rect 463222 392378 463306 392614
rect 463542 392378 498986 392614
rect 499222 392378 499306 392614
rect 499542 392378 534986 392614
rect 535222 392378 535306 392614
rect 535542 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 30986 392294
rect 31222 392058 31306 392294
rect 31542 392058 66986 392294
rect 67222 392058 67306 392294
rect 67542 392058 102986 392294
rect 103222 392058 103306 392294
rect 103542 392058 138986 392294
rect 139222 392058 139306 392294
rect 139542 392058 174986 392294
rect 175222 392058 175306 392294
rect 175542 392058 210986 392294
rect 211222 392058 211306 392294
rect 211542 392058 246986 392294
rect 247222 392058 247306 392294
rect 247542 392058 282986 392294
rect 283222 392058 283306 392294
rect 283542 392058 318986 392294
rect 319222 392058 319306 392294
rect 319542 392058 354986 392294
rect 355222 392058 355306 392294
rect 355542 392058 390986 392294
rect 391222 392058 391306 392294
rect 391542 392058 426986 392294
rect 427222 392058 427306 392294
rect 427542 392058 462986 392294
rect 463222 392058 463306 392294
rect 463542 392058 498986 392294
rect 499222 392058 499306 392294
rect 499542 392058 534986 392294
rect 535222 392058 535306 392294
rect 535542 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 27266 388894
rect 27502 388658 27586 388894
rect 27822 388658 63266 388894
rect 63502 388658 63586 388894
rect 63822 388658 99266 388894
rect 99502 388658 99586 388894
rect 99822 388658 135266 388894
rect 135502 388658 135586 388894
rect 135822 388658 171266 388894
rect 171502 388658 171586 388894
rect 171822 388658 207266 388894
rect 207502 388658 207586 388894
rect 207822 388658 243266 388894
rect 243502 388658 243586 388894
rect 243822 388658 279266 388894
rect 279502 388658 279586 388894
rect 279822 388658 315266 388894
rect 315502 388658 315586 388894
rect 315822 388658 351266 388894
rect 351502 388658 351586 388894
rect 351822 388658 387266 388894
rect 387502 388658 387586 388894
rect 387822 388658 423266 388894
rect 423502 388658 423586 388894
rect 423822 388658 459266 388894
rect 459502 388658 459586 388894
rect 459822 388658 495266 388894
rect 495502 388658 495586 388894
rect 495822 388658 531266 388894
rect 531502 388658 531586 388894
rect 531822 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 27266 388574
rect 27502 388338 27586 388574
rect 27822 388338 63266 388574
rect 63502 388338 63586 388574
rect 63822 388338 99266 388574
rect 99502 388338 99586 388574
rect 99822 388338 135266 388574
rect 135502 388338 135586 388574
rect 135822 388338 171266 388574
rect 171502 388338 171586 388574
rect 171822 388338 207266 388574
rect 207502 388338 207586 388574
rect 207822 388338 243266 388574
rect 243502 388338 243586 388574
rect 243822 388338 279266 388574
rect 279502 388338 279586 388574
rect 279822 388338 315266 388574
rect 315502 388338 315586 388574
rect 315822 388338 351266 388574
rect 351502 388338 351586 388574
rect 351822 388338 387266 388574
rect 387502 388338 387586 388574
rect 387822 388338 423266 388574
rect 423502 388338 423586 388574
rect 423822 388338 459266 388574
rect 459502 388338 459586 388574
rect 459822 388338 495266 388574
rect 495502 388338 495586 388574
rect 495822 388338 531266 388574
rect 531502 388338 531586 388574
rect 531822 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 23546 385174
rect 23782 384938 23866 385174
rect 24102 384938 59546 385174
rect 59782 384938 59866 385174
rect 60102 384938 95546 385174
rect 95782 384938 95866 385174
rect 96102 384938 131546 385174
rect 131782 384938 131866 385174
rect 132102 384938 167546 385174
rect 167782 384938 167866 385174
rect 168102 384938 203546 385174
rect 203782 384938 203866 385174
rect 204102 384938 239546 385174
rect 239782 384938 239866 385174
rect 240102 384938 275546 385174
rect 275782 384938 275866 385174
rect 276102 384938 311546 385174
rect 311782 384938 311866 385174
rect 312102 384938 347546 385174
rect 347782 384938 347866 385174
rect 348102 384938 383546 385174
rect 383782 384938 383866 385174
rect 384102 384938 419546 385174
rect 419782 384938 419866 385174
rect 420102 384938 455546 385174
rect 455782 384938 455866 385174
rect 456102 384938 491546 385174
rect 491782 384938 491866 385174
rect 492102 384938 527546 385174
rect 527782 384938 527866 385174
rect 528102 384938 563546 385174
rect 563782 384938 563866 385174
rect 564102 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 23546 384854
rect 23782 384618 23866 384854
rect 24102 384618 59546 384854
rect 59782 384618 59866 384854
rect 60102 384618 95546 384854
rect 95782 384618 95866 384854
rect 96102 384618 131546 384854
rect 131782 384618 131866 384854
rect 132102 384618 167546 384854
rect 167782 384618 167866 384854
rect 168102 384618 203546 384854
rect 203782 384618 203866 384854
rect 204102 384618 239546 384854
rect 239782 384618 239866 384854
rect 240102 384618 275546 384854
rect 275782 384618 275866 384854
rect 276102 384618 311546 384854
rect 311782 384618 311866 384854
rect 312102 384618 347546 384854
rect 347782 384618 347866 384854
rect 348102 384618 383546 384854
rect 383782 384618 383866 384854
rect 384102 384618 419546 384854
rect 419782 384618 419866 384854
rect 420102 384618 455546 384854
rect 455782 384618 455866 384854
rect 456102 384618 491546 384854
rect 491782 384618 491866 384854
rect 492102 384618 527546 384854
rect 527782 384618 527866 384854
rect 528102 384618 563546 384854
rect 563782 384618 563866 384854
rect 564102 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 19826 381454
rect 20062 381218 20146 381454
rect 20382 381218 55826 381454
rect 56062 381218 56146 381454
rect 56382 381218 91826 381454
rect 92062 381218 92146 381454
rect 92382 381218 127826 381454
rect 128062 381218 128146 381454
rect 128382 381218 163826 381454
rect 164062 381218 164146 381454
rect 164382 381218 199826 381454
rect 200062 381218 200146 381454
rect 200382 381218 235826 381454
rect 236062 381218 236146 381454
rect 236382 381218 271826 381454
rect 272062 381218 272146 381454
rect 272382 381218 307826 381454
rect 308062 381218 308146 381454
rect 308382 381218 343826 381454
rect 344062 381218 344146 381454
rect 344382 381218 379826 381454
rect 380062 381218 380146 381454
rect 380382 381218 415826 381454
rect 416062 381218 416146 381454
rect 416382 381218 451826 381454
rect 452062 381218 452146 381454
rect 452382 381218 487826 381454
rect 488062 381218 488146 381454
rect 488382 381218 523826 381454
rect 524062 381218 524146 381454
rect 524382 381218 559826 381454
rect 560062 381218 560146 381454
rect 560382 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 19826 381134
rect 20062 380898 20146 381134
rect 20382 380898 55826 381134
rect 56062 380898 56146 381134
rect 56382 380898 91826 381134
rect 92062 380898 92146 381134
rect 92382 380898 127826 381134
rect 128062 380898 128146 381134
rect 128382 380898 163826 381134
rect 164062 380898 164146 381134
rect 164382 380898 199826 381134
rect 200062 380898 200146 381134
rect 200382 380898 235826 381134
rect 236062 380898 236146 381134
rect 236382 380898 271826 381134
rect 272062 380898 272146 381134
rect 272382 380898 307826 381134
rect 308062 380898 308146 381134
rect 308382 380898 343826 381134
rect 344062 380898 344146 381134
rect 344382 380898 379826 381134
rect 380062 380898 380146 381134
rect 380382 380898 415826 381134
rect 416062 380898 416146 381134
rect 416382 380898 451826 381134
rect 452062 380898 452146 381134
rect 452382 380898 487826 381134
rect 488062 380898 488146 381134
rect 488382 380898 523826 381134
rect 524062 380898 524146 381134
rect 524382 380898 559826 381134
rect 560062 380898 560146 381134
rect 560382 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 12986 374614
rect 13222 374378 13306 374614
rect 13542 374378 48986 374614
rect 49222 374378 49306 374614
rect 49542 374378 84986 374614
rect 85222 374378 85306 374614
rect 85542 374378 120986 374614
rect 121222 374378 121306 374614
rect 121542 374378 156986 374614
rect 157222 374378 157306 374614
rect 157542 374378 192986 374614
rect 193222 374378 193306 374614
rect 193542 374378 228986 374614
rect 229222 374378 229306 374614
rect 229542 374378 264986 374614
rect 265222 374378 265306 374614
rect 265542 374378 300986 374614
rect 301222 374378 301306 374614
rect 301542 374378 336986 374614
rect 337222 374378 337306 374614
rect 337542 374378 372986 374614
rect 373222 374378 373306 374614
rect 373542 374378 408986 374614
rect 409222 374378 409306 374614
rect 409542 374378 444986 374614
rect 445222 374378 445306 374614
rect 445542 374378 480986 374614
rect 481222 374378 481306 374614
rect 481542 374378 516986 374614
rect 517222 374378 517306 374614
rect 517542 374378 552986 374614
rect 553222 374378 553306 374614
rect 553542 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 12986 374294
rect 13222 374058 13306 374294
rect 13542 374058 48986 374294
rect 49222 374058 49306 374294
rect 49542 374058 84986 374294
rect 85222 374058 85306 374294
rect 85542 374058 120986 374294
rect 121222 374058 121306 374294
rect 121542 374058 156986 374294
rect 157222 374058 157306 374294
rect 157542 374058 192986 374294
rect 193222 374058 193306 374294
rect 193542 374058 228986 374294
rect 229222 374058 229306 374294
rect 229542 374058 264986 374294
rect 265222 374058 265306 374294
rect 265542 374058 300986 374294
rect 301222 374058 301306 374294
rect 301542 374058 336986 374294
rect 337222 374058 337306 374294
rect 337542 374058 372986 374294
rect 373222 374058 373306 374294
rect 373542 374058 408986 374294
rect 409222 374058 409306 374294
rect 409542 374058 444986 374294
rect 445222 374058 445306 374294
rect 445542 374058 480986 374294
rect 481222 374058 481306 374294
rect 481542 374058 516986 374294
rect 517222 374058 517306 374294
rect 517542 374058 552986 374294
rect 553222 374058 553306 374294
rect 553542 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 9266 370894
rect 9502 370658 9586 370894
rect 9822 370658 45266 370894
rect 45502 370658 45586 370894
rect 45822 370658 81266 370894
rect 81502 370658 81586 370894
rect 81822 370658 117266 370894
rect 117502 370658 117586 370894
rect 117822 370658 153266 370894
rect 153502 370658 153586 370894
rect 153822 370658 189266 370894
rect 189502 370658 189586 370894
rect 189822 370658 225266 370894
rect 225502 370658 225586 370894
rect 225822 370658 261266 370894
rect 261502 370658 261586 370894
rect 261822 370658 297266 370894
rect 297502 370658 297586 370894
rect 297822 370658 333266 370894
rect 333502 370658 333586 370894
rect 333822 370658 369266 370894
rect 369502 370658 369586 370894
rect 369822 370658 405266 370894
rect 405502 370658 405586 370894
rect 405822 370658 441266 370894
rect 441502 370658 441586 370894
rect 441822 370658 477266 370894
rect 477502 370658 477586 370894
rect 477822 370658 513266 370894
rect 513502 370658 513586 370894
rect 513822 370658 549266 370894
rect 549502 370658 549586 370894
rect 549822 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 9266 370574
rect 9502 370338 9586 370574
rect 9822 370338 45266 370574
rect 45502 370338 45586 370574
rect 45822 370338 81266 370574
rect 81502 370338 81586 370574
rect 81822 370338 117266 370574
rect 117502 370338 117586 370574
rect 117822 370338 153266 370574
rect 153502 370338 153586 370574
rect 153822 370338 189266 370574
rect 189502 370338 189586 370574
rect 189822 370338 225266 370574
rect 225502 370338 225586 370574
rect 225822 370338 261266 370574
rect 261502 370338 261586 370574
rect 261822 370338 297266 370574
rect 297502 370338 297586 370574
rect 297822 370338 333266 370574
rect 333502 370338 333586 370574
rect 333822 370338 369266 370574
rect 369502 370338 369586 370574
rect 369822 370338 405266 370574
rect 405502 370338 405586 370574
rect 405822 370338 441266 370574
rect 441502 370338 441586 370574
rect 441822 370338 477266 370574
rect 477502 370338 477586 370574
rect 477822 370338 513266 370574
rect 513502 370338 513586 370574
rect 513822 370338 549266 370574
rect 549502 370338 549586 370574
rect 549822 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 5546 367174
rect 5782 366938 5866 367174
rect 6102 366938 41546 367174
rect 41782 366938 41866 367174
rect 42102 366938 77546 367174
rect 77782 366938 77866 367174
rect 78102 366938 113546 367174
rect 113782 366938 113866 367174
rect 114102 366938 149546 367174
rect 149782 366938 149866 367174
rect 150102 366938 185546 367174
rect 185782 366938 185866 367174
rect 186102 366938 221546 367174
rect 221782 366938 221866 367174
rect 222102 366938 257546 367174
rect 257782 366938 257866 367174
rect 258102 366938 293546 367174
rect 293782 366938 293866 367174
rect 294102 366938 329546 367174
rect 329782 366938 329866 367174
rect 330102 366938 365546 367174
rect 365782 366938 365866 367174
rect 366102 366938 401546 367174
rect 401782 366938 401866 367174
rect 402102 366938 437546 367174
rect 437782 366938 437866 367174
rect 438102 366938 473546 367174
rect 473782 366938 473866 367174
rect 474102 366938 509546 367174
rect 509782 366938 509866 367174
rect 510102 366938 545546 367174
rect 545782 366938 545866 367174
rect 546102 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 5546 366854
rect 5782 366618 5866 366854
rect 6102 366618 41546 366854
rect 41782 366618 41866 366854
rect 42102 366618 77546 366854
rect 77782 366618 77866 366854
rect 78102 366618 113546 366854
rect 113782 366618 113866 366854
rect 114102 366618 149546 366854
rect 149782 366618 149866 366854
rect 150102 366618 185546 366854
rect 185782 366618 185866 366854
rect 186102 366618 221546 366854
rect 221782 366618 221866 366854
rect 222102 366618 257546 366854
rect 257782 366618 257866 366854
rect 258102 366618 293546 366854
rect 293782 366618 293866 366854
rect 294102 366618 329546 366854
rect 329782 366618 329866 366854
rect 330102 366618 365546 366854
rect 365782 366618 365866 366854
rect 366102 366618 401546 366854
rect 401782 366618 401866 366854
rect 402102 366618 437546 366854
rect 437782 366618 437866 366854
rect 438102 366618 473546 366854
rect 473782 366618 473866 366854
rect 474102 366618 509546 366854
rect 509782 366618 509866 366854
rect 510102 366618 545546 366854
rect 545782 366618 545866 366854
rect 546102 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 1826 363454
rect 2062 363218 2146 363454
rect 2382 363218 37826 363454
rect 38062 363218 38146 363454
rect 38382 363218 73826 363454
rect 74062 363218 74146 363454
rect 74382 363218 109826 363454
rect 110062 363218 110146 363454
rect 110382 363218 145826 363454
rect 146062 363218 146146 363454
rect 146382 363218 181826 363454
rect 182062 363218 182146 363454
rect 182382 363218 217826 363454
rect 218062 363218 218146 363454
rect 218382 363218 253826 363454
rect 254062 363218 254146 363454
rect 254382 363218 289826 363454
rect 290062 363218 290146 363454
rect 290382 363218 325826 363454
rect 326062 363218 326146 363454
rect 326382 363218 361826 363454
rect 362062 363218 362146 363454
rect 362382 363218 397826 363454
rect 398062 363218 398146 363454
rect 398382 363218 433826 363454
rect 434062 363218 434146 363454
rect 434382 363218 469826 363454
rect 470062 363218 470146 363454
rect 470382 363218 505826 363454
rect 506062 363218 506146 363454
rect 506382 363218 541826 363454
rect 542062 363218 542146 363454
rect 542382 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 1826 363134
rect 2062 362898 2146 363134
rect 2382 362898 37826 363134
rect 38062 362898 38146 363134
rect 38382 362898 73826 363134
rect 74062 362898 74146 363134
rect 74382 362898 109826 363134
rect 110062 362898 110146 363134
rect 110382 362898 145826 363134
rect 146062 362898 146146 363134
rect 146382 362898 181826 363134
rect 182062 362898 182146 363134
rect 182382 362898 217826 363134
rect 218062 362898 218146 363134
rect 218382 362898 253826 363134
rect 254062 362898 254146 363134
rect 254382 362898 289826 363134
rect 290062 362898 290146 363134
rect 290382 362898 325826 363134
rect 326062 362898 326146 363134
rect 326382 362898 361826 363134
rect 362062 362898 362146 363134
rect 362382 362898 397826 363134
rect 398062 362898 398146 363134
rect 398382 362898 433826 363134
rect 434062 362898 434146 363134
rect 434382 362898 469826 363134
rect 470062 362898 470146 363134
rect 470382 362898 505826 363134
rect 506062 362898 506146 363134
rect 506382 362898 541826 363134
rect 542062 362898 542146 363134
rect 542382 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 30986 356614
rect 31222 356378 31306 356614
rect 31542 356378 66986 356614
rect 67222 356378 67306 356614
rect 67542 356378 102986 356614
rect 103222 356378 103306 356614
rect 103542 356378 138986 356614
rect 139222 356378 139306 356614
rect 139542 356378 174986 356614
rect 175222 356378 175306 356614
rect 175542 356378 210986 356614
rect 211222 356378 211306 356614
rect 211542 356378 246986 356614
rect 247222 356378 247306 356614
rect 247542 356378 282986 356614
rect 283222 356378 283306 356614
rect 283542 356378 318986 356614
rect 319222 356378 319306 356614
rect 319542 356378 354986 356614
rect 355222 356378 355306 356614
rect 355542 356378 390986 356614
rect 391222 356378 391306 356614
rect 391542 356378 426986 356614
rect 427222 356378 427306 356614
rect 427542 356378 462986 356614
rect 463222 356378 463306 356614
rect 463542 356378 498986 356614
rect 499222 356378 499306 356614
rect 499542 356378 534986 356614
rect 535222 356378 535306 356614
rect 535542 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 30986 356294
rect 31222 356058 31306 356294
rect 31542 356058 66986 356294
rect 67222 356058 67306 356294
rect 67542 356058 102986 356294
rect 103222 356058 103306 356294
rect 103542 356058 138986 356294
rect 139222 356058 139306 356294
rect 139542 356058 174986 356294
rect 175222 356058 175306 356294
rect 175542 356058 210986 356294
rect 211222 356058 211306 356294
rect 211542 356058 246986 356294
rect 247222 356058 247306 356294
rect 247542 356058 282986 356294
rect 283222 356058 283306 356294
rect 283542 356058 318986 356294
rect 319222 356058 319306 356294
rect 319542 356058 354986 356294
rect 355222 356058 355306 356294
rect 355542 356058 390986 356294
rect 391222 356058 391306 356294
rect 391542 356058 426986 356294
rect 427222 356058 427306 356294
rect 427542 356058 462986 356294
rect 463222 356058 463306 356294
rect 463542 356058 498986 356294
rect 499222 356058 499306 356294
rect 499542 356058 534986 356294
rect 535222 356058 535306 356294
rect 535542 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 27266 352894
rect 27502 352658 27586 352894
rect 27822 352658 63266 352894
rect 63502 352658 63586 352894
rect 63822 352658 99266 352894
rect 99502 352658 99586 352894
rect 99822 352658 135266 352894
rect 135502 352658 135586 352894
rect 135822 352658 171266 352894
rect 171502 352658 171586 352894
rect 171822 352658 207266 352894
rect 207502 352658 207586 352894
rect 207822 352658 243266 352894
rect 243502 352658 243586 352894
rect 243822 352658 279266 352894
rect 279502 352658 279586 352894
rect 279822 352658 315266 352894
rect 315502 352658 315586 352894
rect 315822 352658 351266 352894
rect 351502 352658 351586 352894
rect 351822 352658 387266 352894
rect 387502 352658 387586 352894
rect 387822 352658 423266 352894
rect 423502 352658 423586 352894
rect 423822 352658 459266 352894
rect 459502 352658 459586 352894
rect 459822 352658 495266 352894
rect 495502 352658 495586 352894
rect 495822 352658 531266 352894
rect 531502 352658 531586 352894
rect 531822 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 27266 352574
rect 27502 352338 27586 352574
rect 27822 352338 63266 352574
rect 63502 352338 63586 352574
rect 63822 352338 99266 352574
rect 99502 352338 99586 352574
rect 99822 352338 135266 352574
rect 135502 352338 135586 352574
rect 135822 352338 171266 352574
rect 171502 352338 171586 352574
rect 171822 352338 207266 352574
rect 207502 352338 207586 352574
rect 207822 352338 243266 352574
rect 243502 352338 243586 352574
rect 243822 352338 279266 352574
rect 279502 352338 279586 352574
rect 279822 352338 315266 352574
rect 315502 352338 315586 352574
rect 315822 352338 351266 352574
rect 351502 352338 351586 352574
rect 351822 352338 387266 352574
rect 387502 352338 387586 352574
rect 387822 352338 423266 352574
rect 423502 352338 423586 352574
rect 423822 352338 459266 352574
rect 459502 352338 459586 352574
rect 459822 352338 495266 352574
rect 495502 352338 495586 352574
rect 495822 352338 531266 352574
rect 531502 352338 531586 352574
rect 531822 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 23546 349174
rect 23782 348938 23866 349174
rect 24102 348938 59546 349174
rect 59782 348938 59866 349174
rect 60102 348938 95546 349174
rect 95782 348938 95866 349174
rect 96102 348938 131546 349174
rect 131782 348938 131866 349174
rect 132102 348938 167546 349174
rect 167782 348938 167866 349174
rect 168102 348938 203546 349174
rect 203782 348938 203866 349174
rect 204102 348938 239546 349174
rect 239782 348938 239866 349174
rect 240102 348938 275546 349174
rect 275782 348938 275866 349174
rect 276102 348938 311546 349174
rect 311782 348938 311866 349174
rect 312102 348938 347546 349174
rect 347782 348938 347866 349174
rect 348102 348938 383546 349174
rect 383782 348938 383866 349174
rect 384102 348938 419546 349174
rect 419782 348938 419866 349174
rect 420102 348938 455546 349174
rect 455782 348938 455866 349174
rect 456102 348938 491546 349174
rect 491782 348938 491866 349174
rect 492102 348938 527546 349174
rect 527782 348938 527866 349174
rect 528102 348938 563546 349174
rect 563782 348938 563866 349174
rect 564102 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 23546 348854
rect 23782 348618 23866 348854
rect 24102 348618 59546 348854
rect 59782 348618 59866 348854
rect 60102 348618 95546 348854
rect 95782 348618 95866 348854
rect 96102 348618 131546 348854
rect 131782 348618 131866 348854
rect 132102 348618 167546 348854
rect 167782 348618 167866 348854
rect 168102 348618 203546 348854
rect 203782 348618 203866 348854
rect 204102 348618 239546 348854
rect 239782 348618 239866 348854
rect 240102 348618 275546 348854
rect 275782 348618 275866 348854
rect 276102 348618 311546 348854
rect 311782 348618 311866 348854
rect 312102 348618 347546 348854
rect 347782 348618 347866 348854
rect 348102 348618 383546 348854
rect 383782 348618 383866 348854
rect 384102 348618 419546 348854
rect 419782 348618 419866 348854
rect 420102 348618 455546 348854
rect 455782 348618 455866 348854
rect 456102 348618 491546 348854
rect 491782 348618 491866 348854
rect 492102 348618 527546 348854
rect 527782 348618 527866 348854
rect 528102 348618 563546 348854
rect 563782 348618 563866 348854
rect 564102 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 19826 345454
rect 20062 345218 20146 345454
rect 20382 345218 55826 345454
rect 56062 345218 56146 345454
rect 56382 345218 91826 345454
rect 92062 345218 92146 345454
rect 92382 345218 127826 345454
rect 128062 345218 128146 345454
rect 128382 345218 163826 345454
rect 164062 345218 164146 345454
rect 164382 345218 199826 345454
rect 200062 345218 200146 345454
rect 200382 345218 235826 345454
rect 236062 345218 236146 345454
rect 236382 345218 271826 345454
rect 272062 345218 272146 345454
rect 272382 345218 307826 345454
rect 308062 345218 308146 345454
rect 308382 345218 343826 345454
rect 344062 345218 344146 345454
rect 344382 345218 379826 345454
rect 380062 345218 380146 345454
rect 380382 345218 415826 345454
rect 416062 345218 416146 345454
rect 416382 345218 451826 345454
rect 452062 345218 452146 345454
rect 452382 345218 487826 345454
rect 488062 345218 488146 345454
rect 488382 345218 523826 345454
rect 524062 345218 524146 345454
rect 524382 345218 559826 345454
rect 560062 345218 560146 345454
rect 560382 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 19826 345134
rect 20062 344898 20146 345134
rect 20382 344898 55826 345134
rect 56062 344898 56146 345134
rect 56382 344898 91826 345134
rect 92062 344898 92146 345134
rect 92382 344898 127826 345134
rect 128062 344898 128146 345134
rect 128382 344898 163826 345134
rect 164062 344898 164146 345134
rect 164382 344898 199826 345134
rect 200062 344898 200146 345134
rect 200382 344898 235826 345134
rect 236062 344898 236146 345134
rect 236382 344898 271826 345134
rect 272062 344898 272146 345134
rect 272382 344898 307826 345134
rect 308062 344898 308146 345134
rect 308382 344898 343826 345134
rect 344062 344898 344146 345134
rect 344382 344898 379826 345134
rect 380062 344898 380146 345134
rect 380382 344898 415826 345134
rect 416062 344898 416146 345134
rect 416382 344898 451826 345134
rect 452062 344898 452146 345134
rect 452382 344898 487826 345134
rect 488062 344898 488146 345134
rect 488382 344898 523826 345134
rect 524062 344898 524146 345134
rect 524382 344898 559826 345134
rect 560062 344898 560146 345134
rect 560382 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 12986 338614
rect 13222 338378 13306 338614
rect 13542 338378 48986 338614
rect 49222 338378 49306 338614
rect 49542 338378 84986 338614
rect 85222 338378 85306 338614
rect 85542 338378 120986 338614
rect 121222 338378 121306 338614
rect 121542 338378 156986 338614
rect 157222 338378 157306 338614
rect 157542 338378 192986 338614
rect 193222 338378 193306 338614
rect 193542 338378 228986 338614
rect 229222 338378 229306 338614
rect 229542 338378 264986 338614
rect 265222 338378 265306 338614
rect 265542 338378 300986 338614
rect 301222 338378 301306 338614
rect 301542 338378 336986 338614
rect 337222 338378 337306 338614
rect 337542 338378 372986 338614
rect 373222 338378 373306 338614
rect 373542 338378 408986 338614
rect 409222 338378 409306 338614
rect 409542 338378 444986 338614
rect 445222 338378 445306 338614
rect 445542 338378 480986 338614
rect 481222 338378 481306 338614
rect 481542 338378 516986 338614
rect 517222 338378 517306 338614
rect 517542 338378 552986 338614
rect 553222 338378 553306 338614
rect 553542 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 12986 338294
rect 13222 338058 13306 338294
rect 13542 338058 48986 338294
rect 49222 338058 49306 338294
rect 49542 338058 84986 338294
rect 85222 338058 85306 338294
rect 85542 338058 120986 338294
rect 121222 338058 121306 338294
rect 121542 338058 156986 338294
rect 157222 338058 157306 338294
rect 157542 338058 192986 338294
rect 193222 338058 193306 338294
rect 193542 338058 228986 338294
rect 229222 338058 229306 338294
rect 229542 338058 264986 338294
rect 265222 338058 265306 338294
rect 265542 338058 300986 338294
rect 301222 338058 301306 338294
rect 301542 338058 336986 338294
rect 337222 338058 337306 338294
rect 337542 338058 372986 338294
rect 373222 338058 373306 338294
rect 373542 338058 408986 338294
rect 409222 338058 409306 338294
rect 409542 338058 444986 338294
rect 445222 338058 445306 338294
rect 445542 338058 480986 338294
rect 481222 338058 481306 338294
rect 481542 338058 516986 338294
rect 517222 338058 517306 338294
rect 517542 338058 552986 338294
rect 553222 338058 553306 338294
rect 553542 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 9266 334894
rect 9502 334658 9586 334894
rect 9822 334658 45266 334894
rect 45502 334658 45586 334894
rect 45822 334658 81266 334894
rect 81502 334658 81586 334894
rect 81822 334658 117266 334894
rect 117502 334658 117586 334894
rect 117822 334658 153266 334894
rect 153502 334658 153586 334894
rect 153822 334658 189266 334894
rect 189502 334658 189586 334894
rect 189822 334658 225266 334894
rect 225502 334658 225586 334894
rect 225822 334658 261266 334894
rect 261502 334658 261586 334894
rect 261822 334658 297266 334894
rect 297502 334658 297586 334894
rect 297822 334658 333266 334894
rect 333502 334658 333586 334894
rect 333822 334658 369266 334894
rect 369502 334658 369586 334894
rect 369822 334658 405266 334894
rect 405502 334658 405586 334894
rect 405822 334658 441266 334894
rect 441502 334658 441586 334894
rect 441822 334658 477266 334894
rect 477502 334658 477586 334894
rect 477822 334658 513266 334894
rect 513502 334658 513586 334894
rect 513822 334658 549266 334894
rect 549502 334658 549586 334894
rect 549822 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 9266 334574
rect 9502 334338 9586 334574
rect 9822 334338 45266 334574
rect 45502 334338 45586 334574
rect 45822 334338 81266 334574
rect 81502 334338 81586 334574
rect 81822 334338 117266 334574
rect 117502 334338 117586 334574
rect 117822 334338 153266 334574
rect 153502 334338 153586 334574
rect 153822 334338 189266 334574
rect 189502 334338 189586 334574
rect 189822 334338 225266 334574
rect 225502 334338 225586 334574
rect 225822 334338 261266 334574
rect 261502 334338 261586 334574
rect 261822 334338 297266 334574
rect 297502 334338 297586 334574
rect 297822 334338 333266 334574
rect 333502 334338 333586 334574
rect 333822 334338 369266 334574
rect 369502 334338 369586 334574
rect 369822 334338 405266 334574
rect 405502 334338 405586 334574
rect 405822 334338 441266 334574
rect 441502 334338 441586 334574
rect 441822 334338 477266 334574
rect 477502 334338 477586 334574
rect 477822 334338 513266 334574
rect 513502 334338 513586 334574
rect 513822 334338 549266 334574
rect 549502 334338 549586 334574
rect 549822 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 5546 331174
rect 5782 330938 5866 331174
rect 6102 330938 41546 331174
rect 41782 330938 41866 331174
rect 42102 330938 77546 331174
rect 77782 330938 77866 331174
rect 78102 330938 113546 331174
rect 113782 330938 113866 331174
rect 114102 330938 149546 331174
rect 149782 330938 149866 331174
rect 150102 330938 185546 331174
rect 185782 330938 185866 331174
rect 186102 330938 221546 331174
rect 221782 330938 221866 331174
rect 222102 330938 257546 331174
rect 257782 330938 257866 331174
rect 258102 330938 293546 331174
rect 293782 330938 293866 331174
rect 294102 330938 329546 331174
rect 329782 330938 329866 331174
rect 330102 330938 365546 331174
rect 365782 330938 365866 331174
rect 366102 330938 401546 331174
rect 401782 330938 401866 331174
rect 402102 330938 437546 331174
rect 437782 330938 437866 331174
rect 438102 330938 473546 331174
rect 473782 330938 473866 331174
rect 474102 330938 509546 331174
rect 509782 330938 509866 331174
rect 510102 330938 545546 331174
rect 545782 330938 545866 331174
rect 546102 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 5546 330854
rect 5782 330618 5866 330854
rect 6102 330618 41546 330854
rect 41782 330618 41866 330854
rect 42102 330618 77546 330854
rect 77782 330618 77866 330854
rect 78102 330618 113546 330854
rect 113782 330618 113866 330854
rect 114102 330618 149546 330854
rect 149782 330618 149866 330854
rect 150102 330618 185546 330854
rect 185782 330618 185866 330854
rect 186102 330618 221546 330854
rect 221782 330618 221866 330854
rect 222102 330618 257546 330854
rect 257782 330618 257866 330854
rect 258102 330618 293546 330854
rect 293782 330618 293866 330854
rect 294102 330618 329546 330854
rect 329782 330618 329866 330854
rect 330102 330618 365546 330854
rect 365782 330618 365866 330854
rect 366102 330618 401546 330854
rect 401782 330618 401866 330854
rect 402102 330618 437546 330854
rect 437782 330618 437866 330854
rect 438102 330618 473546 330854
rect 473782 330618 473866 330854
rect 474102 330618 509546 330854
rect 509782 330618 509866 330854
rect 510102 330618 545546 330854
rect 545782 330618 545866 330854
rect 546102 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 1826 327454
rect 2062 327218 2146 327454
rect 2382 327218 37826 327454
rect 38062 327218 38146 327454
rect 38382 327218 73826 327454
rect 74062 327218 74146 327454
rect 74382 327218 109826 327454
rect 110062 327218 110146 327454
rect 110382 327218 145826 327454
rect 146062 327218 146146 327454
rect 146382 327218 181826 327454
rect 182062 327218 182146 327454
rect 182382 327218 217826 327454
rect 218062 327218 218146 327454
rect 218382 327218 253826 327454
rect 254062 327218 254146 327454
rect 254382 327218 289826 327454
rect 290062 327218 290146 327454
rect 290382 327218 325826 327454
rect 326062 327218 326146 327454
rect 326382 327218 361826 327454
rect 362062 327218 362146 327454
rect 362382 327218 397826 327454
rect 398062 327218 398146 327454
rect 398382 327218 433826 327454
rect 434062 327218 434146 327454
rect 434382 327218 469826 327454
rect 470062 327218 470146 327454
rect 470382 327218 505826 327454
rect 506062 327218 506146 327454
rect 506382 327218 541826 327454
rect 542062 327218 542146 327454
rect 542382 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 1826 327134
rect 2062 326898 2146 327134
rect 2382 326898 37826 327134
rect 38062 326898 38146 327134
rect 38382 326898 73826 327134
rect 74062 326898 74146 327134
rect 74382 326898 109826 327134
rect 110062 326898 110146 327134
rect 110382 326898 145826 327134
rect 146062 326898 146146 327134
rect 146382 326898 181826 327134
rect 182062 326898 182146 327134
rect 182382 326898 217826 327134
rect 218062 326898 218146 327134
rect 218382 326898 253826 327134
rect 254062 326898 254146 327134
rect 254382 326898 289826 327134
rect 290062 326898 290146 327134
rect 290382 326898 325826 327134
rect 326062 326898 326146 327134
rect 326382 326898 361826 327134
rect 362062 326898 362146 327134
rect 362382 326898 397826 327134
rect 398062 326898 398146 327134
rect 398382 326898 433826 327134
rect 434062 326898 434146 327134
rect 434382 326898 469826 327134
rect 470062 326898 470146 327134
rect 470382 326898 505826 327134
rect 506062 326898 506146 327134
rect 506382 326898 541826 327134
rect 542062 326898 542146 327134
rect 542382 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 30986 320614
rect 31222 320378 31306 320614
rect 31542 320378 66986 320614
rect 67222 320378 67306 320614
rect 67542 320378 102986 320614
rect 103222 320378 103306 320614
rect 103542 320378 138986 320614
rect 139222 320378 139306 320614
rect 139542 320378 174986 320614
rect 175222 320378 175306 320614
rect 175542 320378 210986 320614
rect 211222 320378 211306 320614
rect 211542 320378 246986 320614
rect 247222 320378 247306 320614
rect 247542 320378 282986 320614
rect 283222 320378 283306 320614
rect 283542 320378 318986 320614
rect 319222 320378 319306 320614
rect 319542 320378 354986 320614
rect 355222 320378 355306 320614
rect 355542 320378 390986 320614
rect 391222 320378 391306 320614
rect 391542 320378 426986 320614
rect 427222 320378 427306 320614
rect 427542 320378 462986 320614
rect 463222 320378 463306 320614
rect 463542 320378 498986 320614
rect 499222 320378 499306 320614
rect 499542 320378 534986 320614
rect 535222 320378 535306 320614
rect 535542 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 30986 320294
rect 31222 320058 31306 320294
rect 31542 320058 66986 320294
rect 67222 320058 67306 320294
rect 67542 320058 102986 320294
rect 103222 320058 103306 320294
rect 103542 320058 138986 320294
rect 139222 320058 139306 320294
rect 139542 320058 174986 320294
rect 175222 320058 175306 320294
rect 175542 320058 210986 320294
rect 211222 320058 211306 320294
rect 211542 320058 246986 320294
rect 247222 320058 247306 320294
rect 247542 320058 282986 320294
rect 283222 320058 283306 320294
rect 283542 320058 318986 320294
rect 319222 320058 319306 320294
rect 319542 320058 354986 320294
rect 355222 320058 355306 320294
rect 355542 320058 390986 320294
rect 391222 320058 391306 320294
rect 391542 320058 426986 320294
rect 427222 320058 427306 320294
rect 427542 320058 462986 320294
rect 463222 320058 463306 320294
rect 463542 320058 498986 320294
rect 499222 320058 499306 320294
rect 499542 320058 534986 320294
rect 535222 320058 535306 320294
rect 535542 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 27266 316894
rect 27502 316658 27586 316894
rect 27822 316658 63266 316894
rect 63502 316658 63586 316894
rect 63822 316658 99266 316894
rect 99502 316658 99586 316894
rect 99822 316658 135266 316894
rect 135502 316658 135586 316894
rect 135822 316658 171266 316894
rect 171502 316658 171586 316894
rect 171822 316658 207266 316894
rect 207502 316658 207586 316894
rect 207822 316658 243266 316894
rect 243502 316658 243586 316894
rect 243822 316658 279266 316894
rect 279502 316658 279586 316894
rect 279822 316658 315266 316894
rect 315502 316658 315586 316894
rect 315822 316658 351266 316894
rect 351502 316658 351586 316894
rect 351822 316658 387266 316894
rect 387502 316658 387586 316894
rect 387822 316658 423266 316894
rect 423502 316658 423586 316894
rect 423822 316658 459266 316894
rect 459502 316658 459586 316894
rect 459822 316658 495266 316894
rect 495502 316658 495586 316894
rect 495822 316658 531266 316894
rect 531502 316658 531586 316894
rect 531822 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 27266 316574
rect 27502 316338 27586 316574
rect 27822 316338 63266 316574
rect 63502 316338 63586 316574
rect 63822 316338 99266 316574
rect 99502 316338 99586 316574
rect 99822 316338 135266 316574
rect 135502 316338 135586 316574
rect 135822 316338 171266 316574
rect 171502 316338 171586 316574
rect 171822 316338 207266 316574
rect 207502 316338 207586 316574
rect 207822 316338 243266 316574
rect 243502 316338 243586 316574
rect 243822 316338 279266 316574
rect 279502 316338 279586 316574
rect 279822 316338 315266 316574
rect 315502 316338 315586 316574
rect 315822 316338 351266 316574
rect 351502 316338 351586 316574
rect 351822 316338 387266 316574
rect 387502 316338 387586 316574
rect 387822 316338 423266 316574
rect 423502 316338 423586 316574
rect 423822 316338 459266 316574
rect 459502 316338 459586 316574
rect 459822 316338 495266 316574
rect 495502 316338 495586 316574
rect 495822 316338 531266 316574
rect 531502 316338 531586 316574
rect 531822 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 23546 313174
rect 23782 312938 23866 313174
rect 24102 312938 59546 313174
rect 59782 312938 59866 313174
rect 60102 312938 95546 313174
rect 95782 312938 95866 313174
rect 96102 312938 131546 313174
rect 131782 312938 131866 313174
rect 132102 312938 167546 313174
rect 167782 312938 167866 313174
rect 168102 312938 203546 313174
rect 203782 312938 203866 313174
rect 204102 312938 239546 313174
rect 239782 312938 239866 313174
rect 240102 312938 275546 313174
rect 275782 312938 275866 313174
rect 276102 312938 311546 313174
rect 311782 312938 311866 313174
rect 312102 312938 347546 313174
rect 347782 312938 347866 313174
rect 348102 312938 383546 313174
rect 383782 312938 383866 313174
rect 384102 312938 419546 313174
rect 419782 312938 419866 313174
rect 420102 312938 455546 313174
rect 455782 312938 455866 313174
rect 456102 312938 491546 313174
rect 491782 312938 491866 313174
rect 492102 312938 527546 313174
rect 527782 312938 527866 313174
rect 528102 312938 563546 313174
rect 563782 312938 563866 313174
rect 564102 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 23546 312854
rect 23782 312618 23866 312854
rect 24102 312618 59546 312854
rect 59782 312618 59866 312854
rect 60102 312618 95546 312854
rect 95782 312618 95866 312854
rect 96102 312618 131546 312854
rect 131782 312618 131866 312854
rect 132102 312618 167546 312854
rect 167782 312618 167866 312854
rect 168102 312618 203546 312854
rect 203782 312618 203866 312854
rect 204102 312618 239546 312854
rect 239782 312618 239866 312854
rect 240102 312618 275546 312854
rect 275782 312618 275866 312854
rect 276102 312618 311546 312854
rect 311782 312618 311866 312854
rect 312102 312618 347546 312854
rect 347782 312618 347866 312854
rect 348102 312618 383546 312854
rect 383782 312618 383866 312854
rect 384102 312618 419546 312854
rect 419782 312618 419866 312854
rect 420102 312618 455546 312854
rect 455782 312618 455866 312854
rect 456102 312618 491546 312854
rect 491782 312618 491866 312854
rect 492102 312618 527546 312854
rect 527782 312618 527866 312854
rect 528102 312618 563546 312854
rect 563782 312618 563866 312854
rect 564102 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 19826 309454
rect 20062 309218 20146 309454
rect 20382 309218 55826 309454
rect 56062 309218 56146 309454
rect 56382 309218 91826 309454
rect 92062 309218 92146 309454
rect 92382 309218 127826 309454
rect 128062 309218 128146 309454
rect 128382 309218 163826 309454
rect 164062 309218 164146 309454
rect 164382 309218 199826 309454
rect 200062 309218 200146 309454
rect 200382 309218 235826 309454
rect 236062 309218 236146 309454
rect 236382 309218 271826 309454
rect 272062 309218 272146 309454
rect 272382 309218 307826 309454
rect 308062 309218 308146 309454
rect 308382 309218 343826 309454
rect 344062 309218 344146 309454
rect 344382 309218 379826 309454
rect 380062 309218 380146 309454
rect 380382 309218 415826 309454
rect 416062 309218 416146 309454
rect 416382 309218 451826 309454
rect 452062 309218 452146 309454
rect 452382 309218 487826 309454
rect 488062 309218 488146 309454
rect 488382 309218 523826 309454
rect 524062 309218 524146 309454
rect 524382 309218 559826 309454
rect 560062 309218 560146 309454
rect 560382 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 19826 309134
rect 20062 308898 20146 309134
rect 20382 308898 55826 309134
rect 56062 308898 56146 309134
rect 56382 308898 91826 309134
rect 92062 308898 92146 309134
rect 92382 308898 127826 309134
rect 128062 308898 128146 309134
rect 128382 308898 163826 309134
rect 164062 308898 164146 309134
rect 164382 308898 199826 309134
rect 200062 308898 200146 309134
rect 200382 308898 235826 309134
rect 236062 308898 236146 309134
rect 236382 308898 271826 309134
rect 272062 308898 272146 309134
rect 272382 308898 307826 309134
rect 308062 308898 308146 309134
rect 308382 308898 343826 309134
rect 344062 308898 344146 309134
rect 344382 308898 379826 309134
rect 380062 308898 380146 309134
rect 380382 308898 415826 309134
rect 416062 308898 416146 309134
rect 416382 308898 451826 309134
rect 452062 308898 452146 309134
rect 452382 308898 487826 309134
rect 488062 308898 488146 309134
rect 488382 308898 523826 309134
rect 524062 308898 524146 309134
rect 524382 308898 559826 309134
rect 560062 308898 560146 309134
rect 560382 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 12986 302614
rect 13222 302378 13306 302614
rect 13542 302378 48986 302614
rect 49222 302378 49306 302614
rect 49542 302378 84986 302614
rect 85222 302378 85306 302614
rect 85542 302378 120986 302614
rect 121222 302378 121306 302614
rect 121542 302378 156986 302614
rect 157222 302378 157306 302614
rect 157542 302378 192986 302614
rect 193222 302378 193306 302614
rect 193542 302378 228986 302614
rect 229222 302378 229306 302614
rect 229542 302378 264986 302614
rect 265222 302378 265306 302614
rect 265542 302378 300986 302614
rect 301222 302378 301306 302614
rect 301542 302378 336986 302614
rect 337222 302378 337306 302614
rect 337542 302378 372986 302614
rect 373222 302378 373306 302614
rect 373542 302378 408986 302614
rect 409222 302378 409306 302614
rect 409542 302378 444986 302614
rect 445222 302378 445306 302614
rect 445542 302378 480986 302614
rect 481222 302378 481306 302614
rect 481542 302378 516986 302614
rect 517222 302378 517306 302614
rect 517542 302378 552986 302614
rect 553222 302378 553306 302614
rect 553542 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 12986 302294
rect 13222 302058 13306 302294
rect 13542 302058 48986 302294
rect 49222 302058 49306 302294
rect 49542 302058 84986 302294
rect 85222 302058 85306 302294
rect 85542 302058 120986 302294
rect 121222 302058 121306 302294
rect 121542 302058 156986 302294
rect 157222 302058 157306 302294
rect 157542 302058 192986 302294
rect 193222 302058 193306 302294
rect 193542 302058 228986 302294
rect 229222 302058 229306 302294
rect 229542 302058 264986 302294
rect 265222 302058 265306 302294
rect 265542 302058 300986 302294
rect 301222 302058 301306 302294
rect 301542 302058 336986 302294
rect 337222 302058 337306 302294
rect 337542 302058 372986 302294
rect 373222 302058 373306 302294
rect 373542 302058 408986 302294
rect 409222 302058 409306 302294
rect 409542 302058 444986 302294
rect 445222 302058 445306 302294
rect 445542 302058 480986 302294
rect 481222 302058 481306 302294
rect 481542 302058 516986 302294
rect 517222 302058 517306 302294
rect 517542 302058 552986 302294
rect 553222 302058 553306 302294
rect 553542 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 9266 298894
rect 9502 298658 9586 298894
rect 9822 298658 45266 298894
rect 45502 298658 45586 298894
rect 45822 298658 81266 298894
rect 81502 298658 81586 298894
rect 81822 298658 117266 298894
rect 117502 298658 117586 298894
rect 117822 298658 153266 298894
rect 153502 298658 153586 298894
rect 153822 298658 189266 298894
rect 189502 298658 189586 298894
rect 189822 298658 225266 298894
rect 225502 298658 225586 298894
rect 225822 298658 261266 298894
rect 261502 298658 261586 298894
rect 261822 298658 297266 298894
rect 297502 298658 297586 298894
rect 297822 298658 333266 298894
rect 333502 298658 333586 298894
rect 333822 298658 369266 298894
rect 369502 298658 369586 298894
rect 369822 298658 405266 298894
rect 405502 298658 405586 298894
rect 405822 298658 441266 298894
rect 441502 298658 441586 298894
rect 441822 298658 477266 298894
rect 477502 298658 477586 298894
rect 477822 298658 513266 298894
rect 513502 298658 513586 298894
rect 513822 298658 549266 298894
rect 549502 298658 549586 298894
rect 549822 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 9266 298574
rect 9502 298338 9586 298574
rect 9822 298338 45266 298574
rect 45502 298338 45586 298574
rect 45822 298338 81266 298574
rect 81502 298338 81586 298574
rect 81822 298338 117266 298574
rect 117502 298338 117586 298574
rect 117822 298338 153266 298574
rect 153502 298338 153586 298574
rect 153822 298338 189266 298574
rect 189502 298338 189586 298574
rect 189822 298338 225266 298574
rect 225502 298338 225586 298574
rect 225822 298338 261266 298574
rect 261502 298338 261586 298574
rect 261822 298338 297266 298574
rect 297502 298338 297586 298574
rect 297822 298338 333266 298574
rect 333502 298338 333586 298574
rect 333822 298338 369266 298574
rect 369502 298338 369586 298574
rect 369822 298338 405266 298574
rect 405502 298338 405586 298574
rect 405822 298338 441266 298574
rect 441502 298338 441586 298574
rect 441822 298338 477266 298574
rect 477502 298338 477586 298574
rect 477822 298338 513266 298574
rect 513502 298338 513586 298574
rect 513822 298338 549266 298574
rect 549502 298338 549586 298574
rect 549822 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 5546 295174
rect 5782 294938 5866 295174
rect 6102 294938 41546 295174
rect 41782 294938 41866 295174
rect 42102 294938 77546 295174
rect 77782 294938 77866 295174
rect 78102 294938 113546 295174
rect 113782 294938 113866 295174
rect 114102 294938 149546 295174
rect 149782 294938 149866 295174
rect 150102 294938 185546 295174
rect 185782 294938 185866 295174
rect 186102 294938 221546 295174
rect 221782 294938 221866 295174
rect 222102 294938 257546 295174
rect 257782 294938 257866 295174
rect 258102 294938 293546 295174
rect 293782 294938 293866 295174
rect 294102 294938 329546 295174
rect 329782 294938 329866 295174
rect 330102 294938 365546 295174
rect 365782 294938 365866 295174
rect 366102 294938 401546 295174
rect 401782 294938 401866 295174
rect 402102 294938 437546 295174
rect 437782 294938 437866 295174
rect 438102 294938 473546 295174
rect 473782 294938 473866 295174
rect 474102 294938 509546 295174
rect 509782 294938 509866 295174
rect 510102 294938 545546 295174
rect 545782 294938 545866 295174
rect 546102 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 5546 294854
rect 5782 294618 5866 294854
rect 6102 294618 41546 294854
rect 41782 294618 41866 294854
rect 42102 294618 77546 294854
rect 77782 294618 77866 294854
rect 78102 294618 113546 294854
rect 113782 294618 113866 294854
rect 114102 294618 149546 294854
rect 149782 294618 149866 294854
rect 150102 294618 185546 294854
rect 185782 294618 185866 294854
rect 186102 294618 221546 294854
rect 221782 294618 221866 294854
rect 222102 294618 257546 294854
rect 257782 294618 257866 294854
rect 258102 294618 293546 294854
rect 293782 294618 293866 294854
rect 294102 294618 329546 294854
rect 329782 294618 329866 294854
rect 330102 294618 365546 294854
rect 365782 294618 365866 294854
rect 366102 294618 401546 294854
rect 401782 294618 401866 294854
rect 402102 294618 437546 294854
rect 437782 294618 437866 294854
rect 438102 294618 473546 294854
rect 473782 294618 473866 294854
rect 474102 294618 509546 294854
rect 509782 294618 509866 294854
rect 510102 294618 545546 294854
rect 545782 294618 545866 294854
rect 546102 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 1826 291454
rect 2062 291218 2146 291454
rect 2382 291218 37826 291454
rect 38062 291218 38146 291454
rect 38382 291218 73826 291454
rect 74062 291218 74146 291454
rect 74382 291218 109826 291454
rect 110062 291218 110146 291454
rect 110382 291218 145826 291454
rect 146062 291218 146146 291454
rect 146382 291218 181826 291454
rect 182062 291218 182146 291454
rect 182382 291218 217826 291454
rect 218062 291218 218146 291454
rect 218382 291218 253826 291454
rect 254062 291218 254146 291454
rect 254382 291218 289826 291454
rect 290062 291218 290146 291454
rect 290382 291218 325826 291454
rect 326062 291218 326146 291454
rect 326382 291218 361826 291454
rect 362062 291218 362146 291454
rect 362382 291218 397826 291454
rect 398062 291218 398146 291454
rect 398382 291218 433826 291454
rect 434062 291218 434146 291454
rect 434382 291218 469826 291454
rect 470062 291218 470146 291454
rect 470382 291218 505826 291454
rect 506062 291218 506146 291454
rect 506382 291218 541826 291454
rect 542062 291218 542146 291454
rect 542382 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 1826 291134
rect 2062 290898 2146 291134
rect 2382 290898 37826 291134
rect 38062 290898 38146 291134
rect 38382 290898 73826 291134
rect 74062 290898 74146 291134
rect 74382 290898 109826 291134
rect 110062 290898 110146 291134
rect 110382 290898 145826 291134
rect 146062 290898 146146 291134
rect 146382 290898 181826 291134
rect 182062 290898 182146 291134
rect 182382 290898 217826 291134
rect 218062 290898 218146 291134
rect 218382 290898 253826 291134
rect 254062 290898 254146 291134
rect 254382 290898 289826 291134
rect 290062 290898 290146 291134
rect 290382 290898 325826 291134
rect 326062 290898 326146 291134
rect 326382 290898 361826 291134
rect 362062 290898 362146 291134
rect 362382 290898 397826 291134
rect 398062 290898 398146 291134
rect 398382 290898 433826 291134
rect 434062 290898 434146 291134
rect 434382 290898 469826 291134
rect 470062 290898 470146 291134
rect 470382 290898 505826 291134
rect 506062 290898 506146 291134
rect 506382 290898 541826 291134
rect 542062 290898 542146 291134
rect 542382 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 30986 284614
rect 31222 284378 31306 284614
rect 31542 284378 66986 284614
rect 67222 284378 67306 284614
rect 67542 284378 102986 284614
rect 103222 284378 103306 284614
rect 103542 284378 138986 284614
rect 139222 284378 139306 284614
rect 139542 284378 174986 284614
rect 175222 284378 175306 284614
rect 175542 284378 210986 284614
rect 211222 284378 211306 284614
rect 211542 284378 246986 284614
rect 247222 284378 247306 284614
rect 247542 284378 282986 284614
rect 283222 284378 283306 284614
rect 283542 284378 318986 284614
rect 319222 284378 319306 284614
rect 319542 284378 354986 284614
rect 355222 284378 355306 284614
rect 355542 284378 390986 284614
rect 391222 284378 391306 284614
rect 391542 284378 426986 284614
rect 427222 284378 427306 284614
rect 427542 284378 462986 284614
rect 463222 284378 463306 284614
rect 463542 284378 498986 284614
rect 499222 284378 499306 284614
rect 499542 284378 534986 284614
rect 535222 284378 535306 284614
rect 535542 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 30986 284294
rect 31222 284058 31306 284294
rect 31542 284058 66986 284294
rect 67222 284058 67306 284294
rect 67542 284058 102986 284294
rect 103222 284058 103306 284294
rect 103542 284058 138986 284294
rect 139222 284058 139306 284294
rect 139542 284058 174986 284294
rect 175222 284058 175306 284294
rect 175542 284058 210986 284294
rect 211222 284058 211306 284294
rect 211542 284058 246986 284294
rect 247222 284058 247306 284294
rect 247542 284058 282986 284294
rect 283222 284058 283306 284294
rect 283542 284058 318986 284294
rect 319222 284058 319306 284294
rect 319542 284058 354986 284294
rect 355222 284058 355306 284294
rect 355542 284058 390986 284294
rect 391222 284058 391306 284294
rect 391542 284058 426986 284294
rect 427222 284058 427306 284294
rect 427542 284058 462986 284294
rect 463222 284058 463306 284294
rect 463542 284058 498986 284294
rect 499222 284058 499306 284294
rect 499542 284058 534986 284294
rect 535222 284058 535306 284294
rect 535542 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 27266 280894
rect 27502 280658 27586 280894
rect 27822 280658 63266 280894
rect 63502 280658 63586 280894
rect 63822 280658 99266 280894
rect 99502 280658 99586 280894
rect 99822 280658 135266 280894
rect 135502 280658 135586 280894
rect 135822 280658 171266 280894
rect 171502 280658 171586 280894
rect 171822 280658 207266 280894
rect 207502 280658 207586 280894
rect 207822 280658 243266 280894
rect 243502 280658 243586 280894
rect 243822 280658 279266 280894
rect 279502 280658 279586 280894
rect 279822 280658 315266 280894
rect 315502 280658 315586 280894
rect 315822 280658 351266 280894
rect 351502 280658 351586 280894
rect 351822 280658 387266 280894
rect 387502 280658 387586 280894
rect 387822 280658 423266 280894
rect 423502 280658 423586 280894
rect 423822 280658 459266 280894
rect 459502 280658 459586 280894
rect 459822 280658 495266 280894
rect 495502 280658 495586 280894
rect 495822 280658 531266 280894
rect 531502 280658 531586 280894
rect 531822 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 27266 280574
rect 27502 280338 27586 280574
rect 27822 280338 63266 280574
rect 63502 280338 63586 280574
rect 63822 280338 99266 280574
rect 99502 280338 99586 280574
rect 99822 280338 135266 280574
rect 135502 280338 135586 280574
rect 135822 280338 171266 280574
rect 171502 280338 171586 280574
rect 171822 280338 207266 280574
rect 207502 280338 207586 280574
rect 207822 280338 243266 280574
rect 243502 280338 243586 280574
rect 243822 280338 279266 280574
rect 279502 280338 279586 280574
rect 279822 280338 315266 280574
rect 315502 280338 315586 280574
rect 315822 280338 351266 280574
rect 351502 280338 351586 280574
rect 351822 280338 387266 280574
rect 387502 280338 387586 280574
rect 387822 280338 423266 280574
rect 423502 280338 423586 280574
rect 423822 280338 459266 280574
rect 459502 280338 459586 280574
rect 459822 280338 495266 280574
rect 495502 280338 495586 280574
rect 495822 280338 531266 280574
rect 531502 280338 531586 280574
rect 531822 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 23546 277174
rect 23782 276938 23866 277174
rect 24102 276938 59546 277174
rect 59782 276938 59866 277174
rect 60102 276938 95546 277174
rect 95782 276938 95866 277174
rect 96102 276938 131546 277174
rect 131782 276938 131866 277174
rect 132102 276938 167546 277174
rect 167782 276938 167866 277174
rect 168102 276938 203546 277174
rect 203782 276938 203866 277174
rect 204102 276938 239546 277174
rect 239782 276938 239866 277174
rect 240102 276938 275546 277174
rect 275782 276938 275866 277174
rect 276102 276938 311546 277174
rect 311782 276938 311866 277174
rect 312102 276938 347546 277174
rect 347782 276938 347866 277174
rect 348102 276938 383546 277174
rect 383782 276938 383866 277174
rect 384102 276938 419546 277174
rect 419782 276938 419866 277174
rect 420102 276938 455546 277174
rect 455782 276938 455866 277174
rect 456102 276938 491546 277174
rect 491782 276938 491866 277174
rect 492102 276938 527546 277174
rect 527782 276938 527866 277174
rect 528102 276938 563546 277174
rect 563782 276938 563866 277174
rect 564102 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 23546 276854
rect 23782 276618 23866 276854
rect 24102 276618 59546 276854
rect 59782 276618 59866 276854
rect 60102 276618 95546 276854
rect 95782 276618 95866 276854
rect 96102 276618 131546 276854
rect 131782 276618 131866 276854
rect 132102 276618 167546 276854
rect 167782 276618 167866 276854
rect 168102 276618 203546 276854
rect 203782 276618 203866 276854
rect 204102 276618 239546 276854
rect 239782 276618 239866 276854
rect 240102 276618 275546 276854
rect 275782 276618 275866 276854
rect 276102 276618 311546 276854
rect 311782 276618 311866 276854
rect 312102 276618 347546 276854
rect 347782 276618 347866 276854
rect 348102 276618 383546 276854
rect 383782 276618 383866 276854
rect 384102 276618 419546 276854
rect 419782 276618 419866 276854
rect 420102 276618 455546 276854
rect 455782 276618 455866 276854
rect 456102 276618 491546 276854
rect 491782 276618 491866 276854
rect 492102 276618 527546 276854
rect 527782 276618 527866 276854
rect 528102 276618 563546 276854
rect 563782 276618 563866 276854
rect 564102 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 19826 273454
rect 20062 273218 20146 273454
rect 20382 273218 55826 273454
rect 56062 273218 56146 273454
rect 56382 273218 91826 273454
rect 92062 273218 92146 273454
rect 92382 273218 127826 273454
rect 128062 273218 128146 273454
rect 128382 273218 163826 273454
rect 164062 273218 164146 273454
rect 164382 273218 199826 273454
rect 200062 273218 200146 273454
rect 200382 273218 235826 273454
rect 236062 273218 236146 273454
rect 236382 273218 271826 273454
rect 272062 273218 272146 273454
rect 272382 273218 307826 273454
rect 308062 273218 308146 273454
rect 308382 273218 343826 273454
rect 344062 273218 344146 273454
rect 344382 273218 379826 273454
rect 380062 273218 380146 273454
rect 380382 273218 415826 273454
rect 416062 273218 416146 273454
rect 416382 273218 451826 273454
rect 452062 273218 452146 273454
rect 452382 273218 487826 273454
rect 488062 273218 488146 273454
rect 488382 273218 523826 273454
rect 524062 273218 524146 273454
rect 524382 273218 559826 273454
rect 560062 273218 560146 273454
rect 560382 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 19826 273134
rect 20062 272898 20146 273134
rect 20382 272898 55826 273134
rect 56062 272898 56146 273134
rect 56382 272898 91826 273134
rect 92062 272898 92146 273134
rect 92382 272898 127826 273134
rect 128062 272898 128146 273134
rect 128382 272898 163826 273134
rect 164062 272898 164146 273134
rect 164382 272898 199826 273134
rect 200062 272898 200146 273134
rect 200382 272898 235826 273134
rect 236062 272898 236146 273134
rect 236382 272898 271826 273134
rect 272062 272898 272146 273134
rect 272382 272898 307826 273134
rect 308062 272898 308146 273134
rect 308382 272898 343826 273134
rect 344062 272898 344146 273134
rect 344382 272898 379826 273134
rect 380062 272898 380146 273134
rect 380382 272898 415826 273134
rect 416062 272898 416146 273134
rect 416382 272898 451826 273134
rect 452062 272898 452146 273134
rect 452382 272898 487826 273134
rect 488062 272898 488146 273134
rect 488382 272898 523826 273134
rect 524062 272898 524146 273134
rect 524382 272898 559826 273134
rect 560062 272898 560146 273134
rect 560382 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 12986 266614
rect 13222 266378 13306 266614
rect 13542 266378 48986 266614
rect 49222 266378 49306 266614
rect 49542 266378 84986 266614
rect 85222 266378 85306 266614
rect 85542 266378 120986 266614
rect 121222 266378 121306 266614
rect 121542 266378 156986 266614
rect 157222 266378 157306 266614
rect 157542 266378 192986 266614
rect 193222 266378 193306 266614
rect 193542 266378 228986 266614
rect 229222 266378 229306 266614
rect 229542 266378 264986 266614
rect 265222 266378 265306 266614
rect 265542 266378 300986 266614
rect 301222 266378 301306 266614
rect 301542 266378 336986 266614
rect 337222 266378 337306 266614
rect 337542 266378 372986 266614
rect 373222 266378 373306 266614
rect 373542 266378 408986 266614
rect 409222 266378 409306 266614
rect 409542 266378 444986 266614
rect 445222 266378 445306 266614
rect 445542 266378 480986 266614
rect 481222 266378 481306 266614
rect 481542 266378 516986 266614
rect 517222 266378 517306 266614
rect 517542 266378 552986 266614
rect 553222 266378 553306 266614
rect 553542 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 12986 266294
rect 13222 266058 13306 266294
rect 13542 266058 48986 266294
rect 49222 266058 49306 266294
rect 49542 266058 84986 266294
rect 85222 266058 85306 266294
rect 85542 266058 120986 266294
rect 121222 266058 121306 266294
rect 121542 266058 156986 266294
rect 157222 266058 157306 266294
rect 157542 266058 192986 266294
rect 193222 266058 193306 266294
rect 193542 266058 228986 266294
rect 229222 266058 229306 266294
rect 229542 266058 264986 266294
rect 265222 266058 265306 266294
rect 265542 266058 300986 266294
rect 301222 266058 301306 266294
rect 301542 266058 336986 266294
rect 337222 266058 337306 266294
rect 337542 266058 372986 266294
rect 373222 266058 373306 266294
rect 373542 266058 408986 266294
rect 409222 266058 409306 266294
rect 409542 266058 444986 266294
rect 445222 266058 445306 266294
rect 445542 266058 480986 266294
rect 481222 266058 481306 266294
rect 481542 266058 516986 266294
rect 517222 266058 517306 266294
rect 517542 266058 552986 266294
rect 553222 266058 553306 266294
rect 553542 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 9266 262894
rect 9502 262658 9586 262894
rect 9822 262658 45266 262894
rect 45502 262658 45586 262894
rect 45822 262658 81266 262894
rect 81502 262658 81586 262894
rect 81822 262658 117266 262894
rect 117502 262658 117586 262894
rect 117822 262658 153266 262894
rect 153502 262658 153586 262894
rect 153822 262658 189266 262894
rect 189502 262658 189586 262894
rect 189822 262658 225266 262894
rect 225502 262658 225586 262894
rect 225822 262658 261266 262894
rect 261502 262658 261586 262894
rect 261822 262658 297266 262894
rect 297502 262658 297586 262894
rect 297822 262658 333266 262894
rect 333502 262658 333586 262894
rect 333822 262658 369266 262894
rect 369502 262658 369586 262894
rect 369822 262658 405266 262894
rect 405502 262658 405586 262894
rect 405822 262658 441266 262894
rect 441502 262658 441586 262894
rect 441822 262658 477266 262894
rect 477502 262658 477586 262894
rect 477822 262658 513266 262894
rect 513502 262658 513586 262894
rect 513822 262658 549266 262894
rect 549502 262658 549586 262894
rect 549822 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 9266 262574
rect 9502 262338 9586 262574
rect 9822 262338 45266 262574
rect 45502 262338 45586 262574
rect 45822 262338 81266 262574
rect 81502 262338 81586 262574
rect 81822 262338 117266 262574
rect 117502 262338 117586 262574
rect 117822 262338 153266 262574
rect 153502 262338 153586 262574
rect 153822 262338 189266 262574
rect 189502 262338 189586 262574
rect 189822 262338 225266 262574
rect 225502 262338 225586 262574
rect 225822 262338 261266 262574
rect 261502 262338 261586 262574
rect 261822 262338 297266 262574
rect 297502 262338 297586 262574
rect 297822 262338 333266 262574
rect 333502 262338 333586 262574
rect 333822 262338 369266 262574
rect 369502 262338 369586 262574
rect 369822 262338 405266 262574
rect 405502 262338 405586 262574
rect 405822 262338 441266 262574
rect 441502 262338 441586 262574
rect 441822 262338 477266 262574
rect 477502 262338 477586 262574
rect 477822 262338 513266 262574
rect 513502 262338 513586 262574
rect 513822 262338 549266 262574
rect 549502 262338 549586 262574
rect 549822 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 5546 259174
rect 5782 258938 5866 259174
rect 6102 258938 41546 259174
rect 41782 258938 41866 259174
rect 42102 258938 77546 259174
rect 77782 258938 77866 259174
rect 78102 258938 113546 259174
rect 113782 258938 113866 259174
rect 114102 258938 149546 259174
rect 149782 258938 149866 259174
rect 150102 258938 185546 259174
rect 185782 258938 185866 259174
rect 186102 258938 221546 259174
rect 221782 258938 221866 259174
rect 222102 258938 257546 259174
rect 257782 258938 257866 259174
rect 258102 258938 293546 259174
rect 293782 258938 293866 259174
rect 294102 258938 329546 259174
rect 329782 258938 329866 259174
rect 330102 258938 365546 259174
rect 365782 258938 365866 259174
rect 366102 258938 401546 259174
rect 401782 258938 401866 259174
rect 402102 258938 437546 259174
rect 437782 258938 437866 259174
rect 438102 258938 473546 259174
rect 473782 258938 473866 259174
rect 474102 258938 509546 259174
rect 509782 258938 509866 259174
rect 510102 258938 545546 259174
rect 545782 258938 545866 259174
rect 546102 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 5546 258854
rect 5782 258618 5866 258854
rect 6102 258618 41546 258854
rect 41782 258618 41866 258854
rect 42102 258618 77546 258854
rect 77782 258618 77866 258854
rect 78102 258618 113546 258854
rect 113782 258618 113866 258854
rect 114102 258618 149546 258854
rect 149782 258618 149866 258854
rect 150102 258618 185546 258854
rect 185782 258618 185866 258854
rect 186102 258618 221546 258854
rect 221782 258618 221866 258854
rect 222102 258618 257546 258854
rect 257782 258618 257866 258854
rect 258102 258618 293546 258854
rect 293782 258618 293866 258854
rect 294102 258618 329546 258854
rect 329782 258618 329866 258854
rect 330102 258618 365546 258854
rect 365782 258618 365866 258854
rect 366102 258618 401546 258854
rect 401782 258618 401866 258854
rect 402102 258618 437546 258854
rect 437782 258618 437866 258854
rect 438102 258618 473546 258854
rect 473782 258618 473866 258854
rect 474102 258618 509546 258854
rect 509782 258618 509866 258854
rect 510102 258618 545546 258854
rect 545782 258618 545866 258854
rect 546102 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 1826 255454
rect 2062 255218 2146 255454
rect 2382 255218 37826 255454
rect 38062 255218 38146 255454
rect 38382 255218 73826 255454
rect 74062 255218 74146 255454
rect 74382 255218 109826 255454
rect 110062 255218 110146 255454
rect 110382 255218 145826 255454
rect 146062 255218 146146 255454
rect 146382 255218 181826 255454
rect 182062 255218 182146 255454
rect 182382 255218 217826 255454
rect 218062 255218 218146 255454
rect 218382 255218 253826 255454
rect 254062 255218 254146 255454
rect 254382 255218 289826 255454
rect 290062 255218 290146 255454
rect 290382 255218 325826 255454
rect 326062 255218 326146 255454
rect 326382 255218 361826 255454
rect 362062 255218 362146 255454
rect 362382 255218 397826 255454
rect 398062 255218 398146 255454
rect 398382 255218 433826 255454
rect 434062 255218 434146 255454
rect 434382 255218 469826 255454
rect 470062 255218 470146 255454
rect 470382 255218 505826 255454
rect 506062 255218 506146 255454
rect 506382 255218 541826 255454
rect 542062 255218 542146 255454
rect 542382 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 1826 255134
rect 2062 254898 2146 255134
rect 2382 254898 37826 255134
rect 38062 254898 38146 255134
rect 38382 254898 73826 255134
rect 74062 254898 74146 255134
rect 74382 254898 109826 255134
rect 110062 254898 110146 255134
rect 110382 254898 145826 255134
rect 146062 254898 146146 255134
rect 146382 254898 181826 255134
rect 182062 254898 182146 255134
rect 182382 254898 217826 255134
rect 218062 254898 218146 255134
rect 218382 254898 253826 255134
rect 254062 254898 254146 255134
rect 254382 254898 289826 255134
rect 290062 254898 290146 255134
rect 290382 254898 325826 255134
rect 326062 254898 326146 255134
rect 326382 254898 361826 255134
rect 362062 254898 362146 255134
rect 362382 254898 397826 255134
rect 398062 254898 398146 255134
rect 398382 254898 433826 255134
rect 434062 254898 434146 255134
rect 434382 254898 469826 255134
rect 470062 254898 470146 255134
rect 470382 254898 505826 255134
rect 506062 254898 506146 255134
rect 506382 254898 541826 255134
rect 542062 254898 542146 255134
rect 542382 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 30986 248614
rect 31222 248378 31306 248614
rect 31542 248378 66986 248614
rect 67222 248378 67306 248614
rect 67542 248378 102986 248614
rect 103222 248378 103306 248614
rect 103542 248378 138986 248614
rect 139222 248378 139306 248614
rect 139542 248378 174986 248614
rect 175222 248378 175306 248614
rect 175542 248378 210986 248614
rect 211222 248378 211306 248614
rect 211542 248378 246986 248614
rect 247222 248378 247306 248614
rect 247542 248378 282986 248614
rect 283222 248378 283306 248614
rect 283542 248378 318986 248614
rect 319222 248378 319306 248614
rect 319542 248378 354986 248614
rect 355222 248378 355306 248614
rect 355542 248378 390986 248614
rect 391222 248378 391306 248614
rect 391542 248378 426986 248614
rect 427222 248378 427306 248614
rect 427542 248378 462986 248614
rect 463222 248378 463306 248614
rect 463542 248378 498986 248614
rect 499222 248378 499306 248614
rect 499542 248378 534986 248614
rect 535222 248378 535306 248614
rect 535542 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 30986 248294
rect 31222 248058 31306 248294
rect 31542 248058 66986 248294
rect 67222 248058 67306 248294
rect 67542 248058 102986 248294
rect 103222 248058 103306 248294
rect 103542 248058 138986 248294
rect 139222 248058 139306 248294
rect 139542 248058 174986 248294
rect 175222 248058 175306 248294
rect 175542 248058 210986 248294
rect 211222 248058 211306 248294
rect 211542 248058 246986 248294
rect 247222 248058 247306 248294
rect 247542 248058 282986 248294
rect 283222 248058 283306 248294
rect 283542 248058 318986 248294
rect 319222 248058 319306 248294
rect 319542 248058 354986 248294
rect 355222 248058 355306 248294
rect 355542 248058 390986 248294
rect 391222 248058 391306 248294
rect 391542 248058 426986 248294
rect 427222 248058 427306 248294
rect 427542 248058 462986 248294
rect 463222 248058 463306 248294
rect 463542 248058 498986 248294
rect 499222 248058 499306 248294
rect 499542 248058 534986 248294
rect 535222 248058 535306 248294
rect 535542 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 27266 244894
rect 27502 244658 27586 244894
rect 27822 244658 63266 244894
rect 63502 244658 63586 244894
rect 63822 244658 99266 244894
rect 99502 244658 99586 244894
rect 99822 244658 135266 244894
rect 135502 244658 135586 244894
rect 135822 244658 171266 244894
rect 171502 244658 171586 244894
rect 171822 244658 207266 244894
rect 207502 244658 207586 244894
rect 207822 244658 243266 244894
rect 243502 244658 243586 244894
rect 243822 244658 279266 244894
rect 279502 244658 279586 244894
rect 279822 244658 315266 244894
rect 315502 244658 315586 244894
rect 315822 244658 351266 244894
rect 351502 244658 351586 244894
rect 351822 244658 387266 244894
rect 387502 244658 387586 244894
rect 387822 244658 423266 244894
rect 423502 244658 423586 244894
rect 423822 244658 459266 244894
rect 459502 244658 459586 244894
rect 459822 244658 495266 244894
rect 495502 244658 495586 244894
rect 495822 244658 531266 244894
rect 531502 244658 531586 244894
rect 531822 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 27266 244574
rect 27502 244338 27586 244574
rect 27822 244338 63266 244574
rect 63502 244338 63586 244574
rect 63822 244338 99266 244574
rect 99502 244338 99586 244574
rect 99822 244338 135266 244574
rect 135502 244338 135586 244574
rect 135822 244338 171266 244574
rect 171502 244338 171586 244574
rect 171822 244338 207266 244574
rect 207502 244338 207586 244574
rect 207822 244338 243266 244574
rect 243502 244338 243586 244574
rect 243822 244338 279266 244574
rect 279502 244338 279586 244574
rect 279822 244338 315266 244574
rect 315502 244338 315586 244574
rect 315822 244338 351266 244574
rect 351502 244338 351586 244574
rect 351822 244338 387266 244574
rect 387502 244338 387586 244574
rect 387822 244338 423266 244574
rect 423502 244338 423586 244574
rect 423822 244338 459266 244574
rect 459502 244338 459586 244574
rect 459822 244338 495266 244574
rect 495502 244338 495586 244574
rect 495822 244338 531266 244574
rect 531502 244338 531586 244574
rect 531822 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 23546 241174
rect 23782 240938 23866 241174
rect 24102 240938 59546 241174
rect 59782 240938 59866 241174
rect 60102 240938 95546 241174
rect 95782 240938 95866 241174
rect 96102 240938 131546 241174
rect 131782 240938 131866 241174
rect 132102 240938 167546 241174
rect 167782 240938 167866 241174
rect 168102 240938 203546 241174
rect 203782 240938 203866 241174
rect 204102 240938 239546 241174
rect 239782 240938 239866 241174
rect 240102 240938 275546 241174
rect 275782 240938 275866 241174
rect 276102 240938 311546 241174
rect 311782 240938 311866 241174
rect 312102 240938 347546 241174
rect 347782 240938 347866 241174
rect 348102 240938 383546 241174
rect 383782 240938 383866 241174
rect 384102 240938 419546 241174
rect 419782 240938 419866 241174
rect 420102 240938 455546 241174
rect 455782 240938 455866 241174
rect 456102 240938 491546 241174
rect 491782 240938 491866 241174
rect 492102 240938 527546 241174
rect 527782 240938 527866 241174
rect 528102 240938 563546 241174
rect 563782 240938 563866 241174
rect 564102 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 23546 240854
rect 23782 240618 23866 240854
rect 24102 240618 59546 240854
rect 59782 240618 59866 240854
rect 60102 240618 95546 240854
rect 95782 240618 95866 240854
rect 96102 240618 131546 240854
rect 131782 240618 131866 240854
rect 132102 240618 167546 240854
rect 167782 240618 167866 240854
rect 168102 240618 203546 240854
rect 203782 240618 203866 240854
rect 204102 240618 239546 240854
rect 239782 240618 239866 240854
rect 240102 240618 275546 240854
rect 275782 240618 275866 240854
rect 276102 240618 311546 240854
rect 311782 240618 311866 240854
rect 312102 240618 347546 240854
rect 347782 240618 347866 240854
rect 348102 240618 383546 240854
rect 383782 240618 383866 240854
rect 384102 240618 419546 240854
rect 419782 240618 419866 240854
rect 420102 240618 455546 240854
rect 455782 240618 455866 240854
rect 456102 240618 491546 240854
rect 491782 240618 491866 240854
rect 492102 240618 527546 240854
rect 527782 240618 527866 240854
rect 528102 240618 563546 240854
rect 563782 240618 563866 240854
rect 564102 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 19826 237454
rect 20062 237218 20146 237454
rect 20382 237218 55826 237454
rect 56062 237218 56146 237454
rect 56382 237218 91826 237454
rect 92062 237218 92146 237454
rect 92382 237218 127826 237454
rect 128062 237218 128146 237454
rect 128382 237218 163826 237454
rect 164062 237218 164146 237454
rect 164382 237218 199826 237454
rect 200062 237218 200146 237454
rect 200382 237218 235826 237454
rect 236062 237218 236146 237454
rect 236382 237218 271826 237454
rect 272062 237218 272146 237454
rect 272382 237218 307826 237454
rect 308062 237218 308146 237454
rect 308382 237218 343826 237454
rect 344062 237218 344146 237454
rect 344382 237218 379826 237454
rect 380062 237218 380146 237454
rect 380382 237218 415826 237454
rect 416062 237218 416146 237454
rect 416382 237218 451826 237454
rect 452062 237218 452146 237454
rect 452382 237218 487826 237454
rect 488062 237218 488146 237454
rect 488382 237218 523826 237454
rect 524062 237218 524146 237454
rect 524382 237218 559826 237454
rect 560062 237218 560146 237454
rect 560382 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 19826 237134
rect 20062 236898 20146 237134
rect 20382 236898 55826 237134
rect 56062 236898 56146 237134
rect 56382 236898 91826 237134
rect 92062 236898 92146 237134
rect 92382 236898 127826 237134
rect 128062 236898 128146 237134
rect 128382 236898 163826 237134
rect 164062 236898 164146 237134
rect 164382 236898 199826 237134
rect 200062 236898 200146 237134
rect 200382 236898 235826 237134
rect 236062 236898 236146 237134
rect 236382 236898 271826 237134
rect 272062 236898 272146 237134
rect 272382 236898 307826 237134
rect 308062 236898 308146 237134
rect 308382 236898 343826 237134
rect 344062 236898 344146 237134
rect 344382 236898 379826 237134
rect 380062 236898 380146 237134
rect 380382 236898 415826 237134
rect 416062 236898 416146 237134
rect 416382 236898 451826 237134
rect 452062 236898 452146 237134
rect 452382 236898 487826 237134
rect 488062 236898 488146 237134
rect 488382 236898 523826 237134
rect 524062 236898 524146 237134
rect 524382 236898 559826 237134
rect 560062 236898 560146 237134
rect 560382 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 12986 230614
rect 13222 230378 13306 230614
rect 13542 230378 48986 230614
rect 49222 230378 49306 230614
rect 49542 230378 84986 230614
rect 85222 230378 85306 230614
rect 85542 230378 120986 230614
rect 121222 230378 121306 230614
rect 121542 230378 156986 230614
rect 157222 230378 157306 230614
rect 157542 230378 192986 230614
rect 193222 230378 193306 230614
rect 193542 230378 228986 230614
rect 229222 230378 229306 230614
rect 229542 230378 264986 230614
rect 265222 230378 265306 230614
rect 265542 230378 300986 230614
rect 301222 230378 301306 230614
rect 301542 230378 336986 230614
rect 337222 230378 337306 230614
rect 337542 230378 372986 230614
rect 373222 230378 373306 230614
rect 373542 230378 408986 230614
rect 409222 230378 409306 230614
rect 409542 230378 444986 230614
rect 445222 230378 445306 230614
rect 445542 230378 480986 230614
rect 481222 230378 481306 230614
rect 481542 230378 516986 230614
rect 517222 230378 517306 230614
rect 517542 230378 552986 230614
rect 553222 230378 553306 230614
rect 553542 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 12986 230294
rect 13222 230058 13306 230294
rect 13542 230058 48986 230294
rect 49222 230058 49306 230294
rect 49542 230058 84986 230294
rect 85222 230058 85306 230294
rect 85542 230058 120986 230294
rect 121222 230058 121306 230294
rect 121542 230058 156986 230294
rect 157222 230058 157306 230294
rect 157542 230058 192986 230294
rect 193222 230058 193306 230294
rect 193542 230058 228986 230294
rect 229222 230058 229306 230294
rect 229542 230058 264986 230294
rect 265222 230058 265306 230294
rect 265542 230058 300986 230294
rect 301222 230058 301306 230294
rect 301542 230058 336986 230294
rect 337222 230058 337306 230294
rect 337542 230058 372986 230294
rect 373222 230058 373306 230294
rect 373542 230058 408986 230294
rect 409222 230058 409306 230294
rect 409542 230058 444986 230294
rect 445222 230058 445306 230294
rect 445542 230058 480986 230294
rect 481222 230058 481306 230294
rect 481542 230058 516986 230294
rect 517222 230058 517306 230294
rect 517542 230058 552986 230294
rect 553222 230058 553306 230294
rect 553542 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 9266 226894
rect 9502 226658 9586 226894
rect 9822 226658 45266 226894
rect 45502 226658 45586 226894
rect 45822 226658 261266 226894
rect 261502 226658 261586 226894
rect 261822 226658 297266 226894
rect 297502 226658 297586 226894
rect 297822 226658 333266 226894
rect 333502 226658 333586 226894
rect 333822 226658 369266 226894
rect 369502 226658 369586 226894
rect 369822 226658 405266 226894
rect 405502 226658 405586 226894
rect 405822 226658 441266 226894
rect 441502 226658 441586 226894
rect 441822 226658 477266 226894
rect 477502 226658 477586 226894
rect 477822 226658 513266 226894
rect 513502 226658 513586 226894
rect 513822 226658 549266 226894
rect 549502 226658 549586 226894
rect 549822 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 9266 226574
rect 9502 226338 9586 226574
rect 9822 226338 45266 226574
rect 45502 226338 45586 226574
rect 45822 226338 261266 226574
rect 261502 226338 261586 226574
rect 261822 226338 297266 226574
rect 297502 226338 297586 226574
rect 297822 226338 333266 226574
rect 333502 226338 333586 226574
rect 333822 226338 369266 226574
rect 369502 226338 369586 226574
rect 369822 226338 405266 226574
rect 405502 226338 405586 226574
rect 405822 226338 441266 226574
rect 441502 226338 441586 226574
rect 441822 226338 477266 226574
rect 477502 226338 477586 226574
rect 477822 226338 513266 226574
rect 513502 226338 513586 226574
rect 513822 226338 549266 226574
rect 549502 226338 549586 226574
rect 549822 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 5546 223174
rect 5782 222938 5866 223174
rect 6102 222938 41546 223174
rect 41782 222938 41866 223174
rect 42102 222938 257546 223174
rect 257782 222938 257866 223174
rect 258102 222938 293546 223174
rect 293782 222938 293866 223174
rect 294102 222938 329546 223174
rect 329782 222938 329866 223174
rect 330102 222938 365546 223174
rect 365782 222938 365866 223174
rect 366102 222938 401546 223174
rect 401782 222938 401866 223174
rect 402102 222938 437546 223174
rect 437782 222938 437866 223174
rect 438102 222938 473546 223174
rect 473782 222938 473866 223174
rect 474102 222938 509546 223174
rect 509782 222938 509866 223174
rect 510102 222938 545546 223174
rect 545782 222938 545866 223174
rect 546102 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 5546 222854
rect 5782 222618 5866 222854
rect 6102 222618 41546 222854
rect 41782 222618 41866 222854
rect 42102 222618 257546 222854
rect 257782 222618 257866 222854
rect 258102 222618 293546 222854
rect 293782 222618 293866 222854
rect 294102 222618 329546 222854
rect 329782 222618 329866 222854
rect 330102 222618 365546 222854
rect 365782 222618 365866 222854
rect 366102 222618 401546 222854
rect 401782 222618 401866 222854
rect 402102 222618 437546 222854
rect 437782 222618 437866 222854
rect 438102 222618 473546 222854
rect 473782 222618 473866 222854
rect 474102 222618 509546 222854
rect 509782 222618 509866 222854
rect 510102 222618 545546 222854
rect 545782 222618 545866 222854
rect 546102 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 1826 219454
rect 2062 219218 2146 219454
rect 2382 219218 37826 219454
rect 38062 219218 38146 219454
rect 38382 219218 64250 219454
rect 64486 219218 94970 219454
rect 95206 219218 125690 219454
rect 125926 219218 156410 219454
rect 156646 219218 187130 219454
rect 187366 219218 217850 219454
rect 218086 219218 253826 219454
rect 254062 219218 254146 219454
rect 254382 219218 289826 219454
rect 290062 219218 290146 219454
rect 290382 219218 325826 219454
rect 326062 219218 326146 219454
rect 326382 219218 361826 219454
rect 362062 219218 362146 219454
rect 362382 219218 397826 219454
rect 398062 219218 398146 219454
rect 398382 219218 433826 219454
rect 434062 219218 434146 219454
rect 434382 219218 469826 219454
rect 470062 219218 470146 219454
rect 470382 219218 505826 219454
rect 506062 219218 506146 219454
rect 506382 219218 541826 219454
rect 542062 219218 542146 219454
rect 542382 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 1826 219134
rect 2062 218898 2146 219134
rect 2382 218898 37826 219134
rect 38062 218898 38146 219134
rect 38382 218898 64250 219134
rect 64486 218898 94970 219134
rect 95206 218898 125690 219134
rect 125926 218898 156410 219134
rect 156646 218898 187130 219134
rect 187366 218898 217850 219134
rect 218086 218898 253826 219134
rect 254062 218898 254146 219134
rect 254382 218898 289826 219134
rect 290062 218898 290146 219134
rect 290382 218898 325826 219134
rect 326062 218898 326146 219134
rect 326382 218898 361826 219134
rect 362062 218898 362146 219134
rect 362382 218898 397826 219134
rect 398062 218898 398146 219134
rect 398382 218898 433826 219134
rect 434062 218898 434146 219134
rect 434382 218898 469826 219134
rect 470062 218898 470146 219134
rect 470382 218898 505826 219134
rect 506062 218898 506146 219134
rect 506382 218898 541826 219134
rect 542062 218898 542146 219134
rect 542382 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 30986 212614
rect 31222 212378 31306 212614
rect 31542 212378 246986 212614
rect 247222 212378 247306 212614
rect 247542 212378 282986 212614
rect 283222 212378 283306 212614
rect 283542 212378 318986 212614
rect 319222 212378 319306 212614
rect 319542 212378 354986 212614
rect 355222 212378 355306 212614
rect 355542 212378 390986 212614
rect 391222 212378 391306 212614
rect 391542 212378 426986 212614
rect 427222 212378 427306 212614
rect 427542 212378 462986 212614
rect 463222 212378 463306 212614
rect 463542 212378 498986 212614
rect 499222 212378 499306 212614
rect 499542 212378 534986 212614
rect 535222 212378 535306 212614
rect 535542 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 30986 212294
rect 31222 212058 31306 212294
rect 31542 212058 246986 212294
rect 247222 212058 247306 212294
rect 247542 212058 282986 212294
rect 283222 212058 283306 212294
rect 283542 212058 318986 212294
rect 319222 212058 319306 212294
rect 319542 212058 354986 212294
rect 355222 212058 355306 212294
rect 355542 212058 390986 212294
rect 391222 212058 391306 212294
rect 391542 212058 426986 212294
rect 427222 212058 427306 212294
rect 427542 212058 462986 212294
rect 463222 212058 463306 212294
rect 463542 212058 498986 212294
rect 499222 212058 499306 212294
rect 499542 212058 534986 212294
rect 535222 212058 535306 212294
rect 535542 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 27266 208894
rect 27502 208658 27586 208894
rect 27822 208658 243266 208894
rect 243502 208658 243586 208894
rect 243822 208658 279266 208894
rect 279502 208658 279586 208894
rect 279822 208658 315266 208894
rect 315502 208658 315586 208894
rect 315822 208658 351266 208894
rect 351502 208658 351586 208894
rect 351822 208658 387266 208894
rect 387502 208658 387586 208894
rect 387822 208658 423266 208894
rect 423502 208658 423586 208894
rect 423822 208658 459266 208894
rect 459502 208658 459586 208894
rect 459822 208658 495266 208894
rect 495502 208658 495586 208894
rect 495822 208658 531266 208894
rect 531502 208658 531586 208894
rect 531822 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 27266 208574
rect 27502 208338 27586 208574
rect 27822 208338 243266 208574
rect 243502 208338 243586 208574
rect 243822 208338 279266 208574
rect 279502 208338 279586 208574
rect 279822 208338 315266 208574
rect 315502 208338 315586 208574
rect 315822 208338 351266 208574
rect 351502 208338 351586 208574
rect 351822 208338 387266 208574
rect 387502 208338 387586 208574
rect 387822 208338 423266 208574
rect 423502 208338 423586 208574
rect 423822 208338 459266 208574
rect 459502 208338 459586 208574
rect 459822 208338 495266 208574
rect 495502 208338 495586 208574
rect 495822 208338 531266 208574
rect 531502 208338 531586 208574
rect 531822 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 23546 205174
rect 23782 204938 23866 205174
rect 24102 204938 239546 205174
rect 239782 204938 239866 205174
rect 240102 204938 275546 205174
rect 275782 204938 275866 205174
rect 276102 204938 311546 205174
rect 311782 204938 311866 205174
rect 312102 204938 347546 205174
rect 347782 204938 347866 205174
rect 348102 204938 383546 205174
rect 383782 204938 383866 205174
rect 384102 204938 419546 205174
rect 419782 204938 419866 205174
rect 420102 204938 455546 205174
rect 455782 204938 455866 205174
rect 456102 204938 491546 205174
rect 491782 204938 491866 205174
rect 492102 204938 527546 205174
rect 527782 204938 527866 205174
rect 528102 204938 563546 205174
rect 563782 204938 563866 205174
rect 564102 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 23546 204854
rect 23782 204618 23866 204854
rect 24102 204618 239546 204854
rect 239782 204618 239866 204854
rect 240102 204618 275546 204854
rect 275782 204618 275866 204854
rect 276102 204618 311546 204854
rect 311782 204618 311866 204854
rect 312102 204618 347546 204854
rect 347782 204618 347866 204854
rect 348102 204618 383546 204854
rect 383782 204618 383866 204854
rect 384102 204618 419546 204854
rect 419782 204618 419866 204854
rect 420102 204618 455546 204854
rect 455782 204618 455866 204854
rect 456102 204618 491546 204854
rect 491782 204618 491866 204854
rect 492102 204618 527546 204854
rect 527782 204618 527866 204854
rect 528102 204618 563546 204854
rect 563782 204618 563866 204854
rect 564102 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 19826 201454
rect 20062 201218 20146 201454
rect 20382 201218 55826 201454
rect 56062 201218 56146 201454
rect 56382 201218 79610 201454
rect 79846 201218 110330 201454
rect 110566 201218 141050 201454
rect 141286 201218 171770 201454
rect 172006 201218 202490 201454
rect 202726 201218 235826 201454
rect 236062 201218 236146 201454
rect 236382 201218 271826 201454
rect 272062 201218 272146 201454
rect 272382 201218 307826 201454
rect 308062 201218 308146 201454
rect 308382 201218 343826 201454
rect 344062 201218 344146 201454
rect 344382 201218 379826 201454
rect 380062 201218 380146 201454
rect 380382 201218 415826 201454
rect 416062 201218 416146 201454
rect 416382 201218 451826 201454
rect 452062 201218 452146 201454
rect 452382 201218 487826 201454
rect 488062 201218 488146 201454
rect 488382 201218 523826 201454
rect 524062 201218 524146 201454
rect 524382 201218 559826 201454
rect 560062 201218 560146 201454
rect 560382 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 19826 201134
rect 20062 200898 20146 201134
rect 20382 200898 55826 201134
rect 56062 200898 56146 201134
rect 56382 200898 79610 201134
rect 79846 200898 110330 201134
rect 110566 200898 141050 201134
rect 141286 200898 171770 201134
rect 172006 200898 202490 201134
rect 202726 200898 235826 201134
rect 236062 200898 236146 201134
rect 236382 200898 271826 201134
rect 272062 200898 272146 201134
rect 272382 200898 307826 201134
rect 308062 200898 308146 201134
rect 308382 200898 343826 201134
rect 344062 200898 344146 201134
rect 344382 200898 379826 201134
rect 380062 200898 380146 201134
rect 380382 200898 415826 201134
rect 416062 200898 416146 201134
rect 416382 200898 451826 201134
rect 452062 200898 452146 201134
rect 452382 200898 487826 201134
rect 488062 200898 488146 201134
rect 488382 200898 523826 201134
rect 524062 200898 524146 201134
rect 524382 200898 559826 201134
rect 560062 200898 560146 201134
rect 560382 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 12986 194614
rect 13222 194378 13306 194614
rect 13542 194378 48986 194614
rect 49222 194378 49306 194614
rect 49542 194378 228986 194614
rect 229222 194378 229306 194614
rect 229542 194378 264986 194614
rect 265222 194378 265306 194614
rect 265542 194378 300986 194614
rect 301222 194378 301306 194614
rect 301542 194378 336986 194614
rect 337222 194378 337306 194614
rect 337542 194378 372986 194614
rect 373222 194378 373306 194614
rect 373542 194378 408986 194614
rect 409222 194378 409306 194614
rect 409542 194378 444986 194614
rect 445222 194378 445306 194614
rect 445542 194378 480986 194614
rect 481222 194378 481306 194614
rect 481542 194378 516986 194614
rect 517222 194378 517306 194614
rect 517542 194378 552986 194614
rect 553222 194378 553306 194614
rect 553542 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 12986 194294
rect 13222 194058 13306 194294
rect 13542 194058 48986 194294
rect 49222 194058 49306 194294
rect 49542 194058 228986 194294
rect 229222 194058 229306 194294
rect 229542 194058 264986 194294
rect 265222 194058 265306 194294
rect 265542 194058 300986 194294
rect 301222 194058 301306 194294
rect 301542 194058 336986 194294
rect 337222 194058 337306 194294
rect 337542 194058 372986 194294
rect 373222 194058 373306 194294
rect 373542 194058 408986 194294
rect 409222 194058 409306 194294
rect 409542 194058 444986 194294
rect 445222 194058 445306 194294
rect 445542 194058 480986 194294
rect 481222 194058 481306 194294
rect 481542 194058 516986 194294
rect 517222 194058 517306 194294
rect 517542 194058 552986 194294
rect 553222 194058 553306 194294
rect 553542 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 9266 190894
rect 9502 190658 9586 190894
rect 9822 190658 45266 190894
rect 45502 190658 45586 190894
rect 45822 190658 261266 190894
rect 261502 190658 261586 190894
rect 261822 190658 297266 190894
rect 297502 190658 297586 190894
rect 297822 190658 333266 190894
rect 333502 190658 333586 190894
rect 333822 190658 369266 190894
rect 369502 190658 369586 190894
rect 369822 190658 405266 190894
rect 405502 190658 405586 190894
rect 405822 190658 441266 190894
rect 441502 190658 441586 190894
rect 441822 190658 477266 190894
rect 477502 190658 477586 190894
rect 477822 190658 513266 190894
rect 513502 190658 513586 190894
rect 513822 190658 549266 190894
rect 549502 190658 549586 190894
rect 549822 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 9266 190574
rect 9502 190338 9586 190574
rect 9822 190338 45266 190574
rect 45502 190338 45586 190574
rect 45822 190338 261266 190574
rect 261502 190338 261586 190574
rect 261822 190338 297266 190574
rect 297502 190338 297586 190574
rect 297822 190338 333266 190574
rect 333502 190338 333586 190574
rect 333822 190338 369266 190574
rect 369502 190338 369586 190574
rect 369822 190338 405266 190574
rect 405502 190338 405586 190574
rect 405822 190338 441266 190574
rect 441502 190338 441586 190574
rect 441822 190338 477266 190574
rect 477502 190338 477586 190574
rect 477822 190338 513266 190574
rect 513502 190338 513586 190574
rect 513822 190338 549266 190574
rect 549502 190338 549586 190574
rect 549822 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 5546 187174
rect 5782 186938 5866 187174
rect 6102 186938 41546 187174
rect 41782 186938 41866 187174
rect 42102 186938 257546 187174
rect 257782 186938 257866 187174
rect 258102 186938 293546 187174
rect 293782 186938 293866 187174
rect 294102 186938 329546 187174
rect 329782 186938 329866 187174
rect 330102 186938 365546 187174
rect 365782 186938 365866 187174
rect 366102 186938 401546 187174
rect 401782 186938 401866 187174
rect 402102 186938 437546 187174
rect 437782 186938 437866 187174
rect 438102 186938 473546 187174
rect 473782 186938 473866 187174
rect 474102 186938 509546 187174
rect 509782 186938 509866 187174
rect 510102 186938 545546 187174
rect 545782 186938 545866 187174
rect 546102 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 5546 186854
rect 5782 186618 5866 186854
rect 6102 186618 41546 186854
rect 41782 186618 41866 186854
rect 42102 186618 257546 186854
rect 257782 186618 257866 186854
rect 258102 186618 293546 186854
rect 293782 186618 293866 186854
rect 294102 186618 329546 186854
rect 329782 186618 329866 186854
rect 330102 186618 365546 186854
rect 365782 186618 365866 186854
rect 366102 186618 401546 186854
rect 401782 186618 401866 186854
rect 402102 186618 437546 186854
rect 437782 186618 437866 186854
rect 438102 186618 473546 186854
rect 473782 186618 473866 186854
rect 474102 186618 509546 186854
rect 509782 186618 509866 186854
rect 510102 186618 545546 186854
rect 545782 186618 545866 186854
rect 546102 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 1826 183454
rect 2062 183218 2146 183454
rect 2382 183218 37826 183454
rect 38062 183218 38146 183454
rect 38382 183218 64250 183454
rect 64486 183218 94970 183454
rect 95206 183218 125690 183454
rect 125926 183218 156410 183454
rect 156646 183218 187130 183454
rect 187366 183218 217850 183454
rect 218086 183218 253826 183454
rect 254062 183218 254146 183454
rect 254382 183218 289826 183454
rect 290062 183218 290146 183454
rect 290382 183218 325826 183454
rect 326062 183218 326146 183454
rect 326382 183218 361826 183454
rect 362062 183218 362146 183454
rect 362382 183218 397826 183454
rect 398062 183218 398146 183454
rect 398382 183218 433826 183454
rect 434062 183218 434146 183454
rect 434382 183218 469826 183454
rect 470062 183218 470146 183454
rect 470382 183218 505826 183454
rect 506062 183218 506146 183454
rect 506382 183218 541826 183454
rect 542062 183218 542146 183454
rect 542382 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 1826 183134
rect 2062 182898 2146 183134
rect 2382 182898 37826 183134
rect 38062 182898 38146 183134
rect 38382 182898 64250 183134
rect 64486 182898 94970 183134
rect 95206 182898 125690 183134
rect 125926 182898 156410 183134
rect 156646 182898 187130 183134
rect 187366 182898 217850 183134
rect 218086 182898 253826 183134
rect 254062 182898 254146 183134
rect 254382 182898 289826 183134
rect 290062 182898 290146 183134
rect 290382 182898 325826 183134
rect 326062 182898 326146 183134
rect 326382 182898 361826 183134
rect 362062 182898 362146 183134
rect 362382 182898 397826 183134
rect 398062 182898 398146 183134
rect 398382 182898 433826 183134
rect 434062 182898 434146 183134
rect 434382 182898 469826 183134
rect 470062 182898 470146 183134
rect 470382 182898 505826 183134
rect 506062 182898 506146 183134
rect 506382 182898 541826 183134
rect 542062 182898 542146 183134
rect 542382 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 30986 176614
rect 31222 176378 31306 176614
rect 31542 176378 246986 176614
rect 247222 176378 247306 176614
rect 247542 176378 282986 176614
rect 283222 176378 283306 176614
rect 283542 176378 318986 176614
rect 319222 176378 319306 176614
rect 319542 176378 354986 176614
rect 355222 176378 355306 176614
rect 355542 176378 390986 176614
rect 391222 176378 391306 176614
rect 391542 176378 426986 176614
rect 427222 176378 427306 176614
rect 427542 176378 462986 176614
rect 463222 176378 463306 176614
rect 463542 176378 498986 176614
rect 499222 176378 499306 176614
rect 499542 176378 534986 176614
rect 535222 176378 535306 176614
rect 535542 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 30986 176294
rect 31222 176058 31306 176294
rect 31542 176058 246986 176294
rect 247222 176058 247306 176294
rect 247542 176058 282986 176294
rect 283222 176058 283306 176294
rect 283542 176058 318986 176294
rect 319222 176058 319306 176294
rect 319542 176058 354986 176294
rect 355222 176058 355306 176294
rect 355542 176058 390986 176294
rect 391222 176058 391306 176294
rect 391542 176058 426986 176294
rect 427222 176058 427306 176294
rect 427542 176058 462986 176294
rect 463222 176058 463306 176294
rect 463542 176058 498986 176294
rect 499222 176058 499306 176294
rect 499542 176058 534986 176294
rect 535222 176058 535306 176294
rect 535542 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 27266 172894
rect 27502 172658 27586 172894
rect 27822 172658 243266 172894
rect 243502 172658 243586 172894
rect 243822 172658 279266 172894
rect 279502 172658 279586 172894
rect 279822 172658 315266 172894
rect 315502 172658 315586 172894
rect 315822 172658 351266 172894
rect 351502 172658 351586 172894
rect 351822 172658 387266 172894
rect 387502 172658 387586 172894
rect 387822 172658 423266 172894
rect 423502 172658 423586 172894
rect 423822 172658 459266 172894
rect 459502 172658 459586 172894
rect 459822 172658 495266 172894
rect 495502 172658 495586 172894
rect 495822 172658 531266 172894
rect 531502 172658 531586 172894
rect 531822 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 27266 172574
rect 27502 172338 27586 172574
rect 27822 172338 243266 172574
rect 243502 172338 243586 172574
rect 243822 172338 279266 172574
rect 279502 172338 279586 172574
rect 279822 172338 315266 172574
rect 315502 172338 315586 172574
rect 315822 172338 351266 172574
rect 351502 172338 351586 172574
rect 351822 172338 387266 172574
rect 387502 172338 387586 172574
rect 387822 172338 423266 172574
rect 423502 172338 423586 172574
rect 423822 172338 459266 172574
rect 459502 172338 459586 172574
rect 459822 172338 495266 172574
rect 495502 172338 495586 172574
rect 495822 172338 531266 172574
rect 531502 172338 531586 172574
rect 531822 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 23546 169174
rect 23782 168938 23866 169174
rect 24102 168938 239546 169174
rect 239782 168938 239866 169174
rect 240102 168938 275546 169174
rect 275782 168938 275866 169174
rect 276102 168938 311546 169174
rect 311782 168938 311866 169174
rect 312102 168938 347546 169174
rect 347782 168938 347866 169174
rect 348102 168938 383546 169174
rect 383782 168938 383866 169174
rect 384102 168938 419546 169174
rect 419782 168938 419866 169174
rect 420102 168938 455546 169174
rect 455782 168938 455866 169174
rect 456102 168938 491546 169174
rect 491782 168938 491866 169174
rect 492102 168938 527546 169174
rect 527782 168938 527866 169174
rect 528102 168938 563546 169174
rect 563782 168938 563866 169174
rect 564102 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 23546 168854
rect 23782 168618 23866 168854
rect 24102 168618 239546 168854
rect 239782 168618 239866 168854
rect 240102 168618 275546 168854
rect 275782 168618 275866 168854
rect 276102 168618 311546 168854
rect 311782 168618 311866 168854
rect 312102 168618 347546 168854
rect 347782 168618 347866 168854
rect 348102 168618 383546 168854
rect 383782 168618 383866 168854
rect 384102 168618 419546 168854
rect 419782 168618 419866 168854
rect 420102 168618 455546 168854
rect 455782 168618 455866 168854
rect 456102 168618 491546 168854
rect 491782 168618 491866 168854
rect 492102 168618 527546 168854
rect 527782 168618 527866 168854
rect 528102 168618 563546 168854
rect 563782 168618 563866 168854
rect 564102 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 19826 165454
rect 20062 165218 20146 165454
rect 20382 165218 55826 165454
rect 56062 165218 56146 165454
rect 56382 165218 79610 165454
rect 79846 165218 110330 165454
rect 110566 165218 141050 165454
rect 141286 165218 171770 165454
rect 172006 165218 202490 165454
rect 202726 165218 235826 165454
rect 236062 165218 236146 165454
rect 236382 165218 271826 165454
rect 272062 165218 272146 165454
rect 272382 165218 307826 165454
rect 308062 165218 308146 165454
rect 308382 165218 343826 165454
rect 344062 165218 344146 165454
rect 344382 165218 379826 165454
rect 380062 165218 380146 165454
rect 380382 165218 415826 165454
rect 416062 165218 416146 165454
rect 416382 165218 451826 165454
rect 452062 165218 452146 165454
rect 452382 165218 487826 165454
rect 488062 165218 488146 165454
rect 488382 165218 523826 165454
rect 524062 165218 524146 165454
rect 524382 165218 559826 165454
rect 560062 165218 560146 165454
rect 560382 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 19826 165134
rect 20062 164898 20146 165134
rect 20382 164898 55826 165134
rect 56062 164898 56146 165134
rect 56382 164898 79610 165134
rect 79846 164898 110330 165134
rect 110566 164898 141050 165134
rect 141286 164898 171770 165134
rect 172006 164898 202490 165134
rect 202726 164898 235826 165134
rect 236062 164898 236146 165134
rect 236382 164898 271826 165134
rect 272062 164898 272146 165134
rect 272382 164898 307826 165134
rect 308062 164898 308146 165134
rect 308382 164898 343826 165134
rect 344062 164898 344146 165134
rect 344382 164898 379826 165134
rect 380062 164898 380146 165134
rect 380382 164898 415826 165134
rect 416062 164898 416146 165134
rect 416382 164898 451826 165134
rect 452062 164898 452146 165134
rect 452382 164898 487826 165134
rect 488062 164898 488146 165134
rect 488382 164898 523826 165134
rect 524062 164898 524146 165134
rect 524382 164898 559826 165134
rect 560062 164898 560146 165134
rect 560382 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 12986 158614
rect 13222 158378 13306 158614
rect 13542 158378 48986 158614
rect 49222 158378 49306 158614
rect 49542 158378 228986 158614
rect 229222 158378 229306 158614
rect 229542 158378 264986 158614
rect 265222 158378 265306 158614
rect 265542 158378 300986 158614
rect 301222 158378 301306 158614
rect 301542 158378 336986 158614
rect 337222 158378 337306 158614
rect 337542 158378 372986 158614
rect 373222 158378 373306 158614
rect 373542 158378 408986 158614
rect 409222 158378 409306 158614
rect 409542 158378 444986 158614
rect 445222 158378 445306 158614
rect 445542 158378 480986 158614
rect 481222 158378 481306 158614
rect 481542 158378 516986 158614
rect 517222 158378 517306 158614
rect 517542 158378 552986 158614
rect 553222 158378 553306 158614
rect 553542 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 12986 158294
rect 13222 158058 13306 158294
rect 13542 158058 48986 158294
rect 49222 158058 49306 158294
rect 49542 158058 228986 158294
rect 229222 158058 229306 158294
rect 229542 158058 264986 158294
rect 265222 158058 265306 158294
rect 265542 158058 300986 158294
rect 301222 158058 301306 158294
rect 301542 158058 336986 158294
rect 337222 158058 337306 158294
rect 337542 158058 372986 158294
rect 373222 158058 373306 158294
rect 373542 158058 408986 158294
rect 409222 158058 409306 158294
rect 409542 158058 444986 158294
rect 445222 158058 445306 158294
rect 445542 158058 480986 158294
rect 481222 158058 481306 158294
rect 481542 158058 516986 158294
rect 517222 158058 517306 158294
rect 517542 158058 552986 158294
rect 553222 158058 553306 158294
rect 553542 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 9266 154894
rect 9502 154658 9586 154894
rect 9822 154658 45266 154894
rect 45502 154658 45586 154894
rect 45822 154658 261266 154894
rect 261502 154658 261586 154894
rect 261822 154658 297266 154894
rect 297502 154658 297586 154894
rect 297822 154658 333266 154894
rect 333502 154658 333586 154894
rect 333822 154658 369266 154894
rect 369502 154658 369586 154894
rect 369822 154658 405266 154894
rect 405502 154658 405586 154894
rect 405822 154658 441266 154894
rect 441502 154658 441586 154894
rect 441822 154658 477266 154894
rect 477502 154658 477586 154894
rect 477822 154658 513266 154894
rect 513502 154658 513586 154894
rect 513822 154658 549266 154894
rect 549502 154658 549586 154894
rect 549822 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 9266 154574
rect 9502 154338 9586 154574
rect 9822 154338 45266 154574
rect 45502 154338 45586 154574
rect 45822 154338 261266 154574
rect 261502 154338 261586 154574
rect 261822 154338 297266 154574
rect 297502 154338 297586 154574
rect 297822 154338 333266 154574
rect 333502 154338 333586 154574
rect 333822 154338 369266 154574
rect 369502 154338 369586 154574
rect 369822 154338 405266 154574
rect 405502 154338 405586 154574
rect 405822 154338 441266 154574
rect 441502 154338 441586 154574
rect 441822 154338 477266 154574
rect 477502 154338 477586 154574
rect 477822 154338 513266 154574
rect 513502 154338 513586 154574
rect 513822 154338 549266 154574
rect 549502 154338 549586 154574
rect 549822 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 5546 151174
rect 5782 150938 5866 151174
rect 6102 150938 41546 151174
rect 41782 150938 41866 151174
rect 42102 150938 257546 151174
rect 257782 150938 257866 151174
rect 258102 150938 293546 151174
rect 293782 150938 293866 151174
rect 294102 150938 329546 151174
rect 329782 150938 329866 151174
rect 330102 150938 365546 151174
rect 365782 150938 365866 151174
rect 366102 150938 401546 151174
rect 401782 150938 401866 151174
rect 402102 150938 437546 151174
rect 437782 150938 437866 151174
rect 438102 150938 473546 151174
rect 473782 150938 473866 151174
rect 474102 150938 509546 151174
rect 509782 150938 509866 151174
rect 510102 150938 545546 151174
rect 545782 150938 545866 151174
rect 546102 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 5546 150854
rect 5782 150618 5866 150854
rect 6102 150618 41546 150854
rect 41782 150618 41866 150854
rect 42102 150618 257546 150854
rect 257782 150618 257866 150854
rect 258102 150618 293546 150854
rect 293782 150618 293866 150854
rect 294102 150618 329546 150854
rect 329782 150618 329866 150854
rect 330102 150618 365546 150854
rect 365782 150618 365866 150854
rect 366102 150618 401546 150854
rect 401782 150618 401866 150854
rect 402102 150618 437546 150854
rect 437782 150618 437866 150854
rect 438102 150618 473546 150854
rect 473782 150618 473866 150854
rect 474102 150618 509546 150854
rect 509782 150618 509866 150854
rect 510102 150618 545546 150854
rect 545782 150618 545866 150854
rect 546102 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 1826 147454
rect 2062 147218 2146 147454
rect 2382 147218 37826 147454
rect 38062 147218 38146 147454
rect 38382 147218 64250 147454
rect 64486 147218 94970 147454
rect 95206 147218 125690 147454
rect 125926 147218 156410 147454
rect 156646 147218 187130 147454
rect 187366 147218 217850 147454
rect 218086 147218 253826 147454
rect 254062 147218 254146 147454
rect 254382 147218 289826 147454
rect 290062 147218 290146 147454
rect 290382 147218 325826 147454
rect 326062 147218 326146 147454
rect 326382 147218 361826 147454
rect 362062 147218 362146 147454
rect 362382 147218 397826 147454
rect 398062 147218 398146 147454
rect 398382 147218 433826 147454
rect 434062 147218 434146 147454
rect 434382 147218 469826 147454
rect 470062 147218 470146 147454
rect 470382 147218 505826 147454
rect 506062 147218 506146 147454
rect 506382 147218 541826 147454
rect 542062 147218 542146 147454
rect 542382 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 1826 147134
rect 2062 146898 2146 147134
rect 2382 146898 37826 147134
rect 38062 146898 38146 147134
rect 38382 146898 64250 147134
rect 64486 146898 94970 147134
rect 95206 146898 125690 147134
rect 125926 146898 156410 147134
rect 156646 146898 187130 147134
rect 187366 146898 217850 147134
rect 218086 146898 253826 147134
rect 254062 146898 254146 147134
rect 254382 146898 289826 147134
rect 290062 146898 290146 147134
rect 290382 146898 325826 147134
rect 326062 146898 326146 147134
rect 326382 146898 361826 147134
rect 362062 146898 362146 147134
rect 362382 146898 397826 147134
rect 398062 146898 398146 147134
rect 398382 146898 433826 147134
rect 434062 146898 434146 147134
rect 434382 146898 469826 147134
rect 470062 146898 470146 147134
rect 470382 146898 505826 147134
rect 506062 146898 506146 147134
rect 506382 146898 541826 147134
rect 542062 146898 542146 147134
rect 542382 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 30986 140614
rect 31222 140378 31306 140614
rect 31542 140378 246986 140614
rect 247222 140378 247306 140614
rect 247542 140378 282986 140614
rect 283222 140378 283306 140614
rect 283542 140378 318986 140614
rect 319222 140378 319306 140614
rect 319542 140378 354986 140614
rect 355222 140378 355306 140614
rect 355542 140378 390986 140614
rect 391222 140378 391306 140614
rect 391542 140378 426986 140614
rect 427222 140378 427306 140614
rect 427542 140378 462986 140614
rect 463222 140378 463306 140614
rect 463542 140378 498986 140614
rect 499222 140378 499306 140614
rect 499542 140378 534986 140614
rect 535222 140378 535306 140614
rect 535542 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 30986 140294
rect 31222 140058 31306 140294
rect 31542 140058 246986 140294
rect 247222 140058 247306 140294
rect 247542 140058 282986 140294
rect 283222 140058 283306 140294
rect 283542 140058 318986 140294
rect 319222 140058 319306 140294
rect 319542 140058 354986 140294
rect 355222 140058 355306 140294
rect 355542 140058 390986 140294
rect 391222 140058 391306 140294
rect 391542 140058 426986 140294
rect 427222 140058 427306 140294
rect 427542 140058 462986 140294
rect 463222 140058 463306 140294
rect 463542 140058 498986 140294
rect 499222 140058 499306 140294
rect 499542 140058 534986 140294
rect 535222 140058 535306 140294
rect 535542 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 27266 136894
rect 27502 136658 27586 136894
rect 27822 136658 243266 136894
rect 243502 136658 243586 136894
rect 243822 136658 279266 136894
rect 279502 136658 279586 136894
rect 279822 136658 315266 136894
rect 315502 136658 315586 136894
rect 315822 136658 351266 136894
rect 351502 136658 351586 136894
rect 351822 136658 387266 136894
rect 387502 136658 387586 136894
rect 387822 136658 423266 136894
rect 423502 136658 423586 136894
rect 423822 136658 459266 136894
rect 459502 136658 459586 136894
rect 459822 136658 495266 136894
rect 495502 136658 495586 136894
rect 495822 136658 531266 136894
rect 531502 136658 531586 136894
rect 531822 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 27266 136574
rect 27502 136338 27586 136574
rect 27822 136338 243266 136574
rect 243502 136338 243586 136574
rect 243822 136338 279266 136574
rect 279502 136338 279586 136574
rect 279822 136338 315266 136574
rect 315502 136338 315586 136574
rect 315822 136338 351266 136574
rect 351502 136338 351586 136574
rect 351822 136338 387266 136574
rect 387502 136338 387586 136574
rect 387822 136338 423266 136574
rect 423502 136338 423586 136574
rect 423822 136338 459266 136574
rect 459502 136338 459586 136574
rect 459822 136338 495266 136574
rect 495502 136338 495586 136574
rect 495822 136338 531266 136574
rect 531502 136338 531586 136574
rect 531822 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 23546 133174
rect 23782 132938 23866 133174
rect 24102 132938 239546 133174
rect 239782 132938 239866 133174
rect 240102 132938 275546 133174
rect 275782 132938 275866 133174
rect 276102 132938 311546 133174
rect 311782 132938 311866 133174
rect 312102 132938 347546 133174
rect 347782 132938 347866 133174
rect 348102 132938 383546 133174
rect 383782 132938 383866 133174
rect 384102 132938 419546 133174
rect 419782 132938 419866 133174
rect 420102 132938 455546 133174
rect 455782 132938 455866 133174
rect 456102 132938 491546 133174
rect 491782 132938 491866 133174
rect 492102 132938 527546 133174
rect 527782 132938 527866 133174
rect 528102 132938 563546 133174
rect 563782 132938 563866 133174
rect 564102 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 23546 132854
rect 23782 132618 23866 132854
rect 24102 132618 239546 132854
rect 239782 132618 239866 132854
rect 240102 132618 275546 132854
rect 275782 132618 275866 132854
rect 276102 132618 311546 132854
rect 311782 132618 311866 132854
rect 312102 132618 347546 132854
rect 347782 132618 347866 132854
rect 348102 132618 383546 132854
rect 383782 132618 383866 132854
rect 384102 132618 419546 132854
rect 419782 132618 419866 132854
rect 420102 132618 455546 132854
rect 455782 132618 455866 132854
rect 456102 132618 491546 132854
rect 491782 132618 491866 132854
rect 492102 132618 527546 132854
rect 527782 132618 527866 132854
rect 528102 132618 563546 132854
rect 563782 132618 563866 132854
rect 564102 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 19826 129454
rect 20062 129218 20146 129454
rect 20382 129218 55826 129454
rect 56062 129218 56146 129454
rect 56382 129218 79610 129454
rect 79846 129218 110330 129454
rect 110566 129218 141050 129454
rect 141286 129218 171770 129454
rect 172006 129218 202490 129454
rect 202726 129218 235826 129454
rect 236062 129218 236146 129454
rect 236382 129218 271826 129454
rect 272062 129218 272146 129454
rect 272382 129218 307826 129454
rect 308062 129218 308146 129454
rect 308382 129218 343826 129454
rect 344062 129218 344146 129454
rect 344382 129218 379826 129454
rect 380062 129218 380146 129454
rect 380382 129218 415826 129454
rect 416062 129218 416146 129454
rect 416382 129218 451826 129454
rect 452062 129218 452146 129454
rect 452382 129218 487826 129454
rect 488062 129218 488146 129454
rect 488382 129218 523826 129454
rect 524062 129218 524146 129454
rect 524382 129218 559826 129454
rect 560062 129218 560146 129454
rect 560382 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 19826 129134
rect 20062 128898 20146 129134
rect 20382 128898 55826 129134
rect 56062 128898 56146 129134
rect 56382 128898 79610 129134
rect 79846 128898 110330 129134
rect 110566 128898 141050 129134
rect 141286 128898 171770 129134
rect 172006 128898 202490 129134
rect 202726 128898 235826 129134
rect 236062 128898 236146 129134
rect 236382 128898 271826 129134
rect 272062 128898 272146 129134
rect 272382 128898 307826 129134
rect 308062 128898 308146 129134
rect 308382 128898 343826 129134
rect 344062 128898 344146 129134
rect 344382 128898 379826 129134
rect 380062 128898 380146 129134
rect 380382 128898 415826 129134
rect 416062 128898 416146 129134
rect 416382 128898 451826 129134
rect 452062 128898 452146 129134
rect 452382 128898 487826 129134
rect 488062 128898 488146 129134
rect 488382 128898 523826 129134
rect 524062 128898 524146 129134
rect 524382 128898 559826 129134
rect 560062 128898 560146 129134
rect 560382 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 12986 122614
rect 13222 122378 13306 122614
rect 13542 122378 48986 122614
rect 49222 122378 49306 122614
rect 49542 122378 228986 122614
rect 229222 122378 229306 122614
rect 229542 122378 264986 122614
rect 265222 122378 265306 122614
rect 265542 122378 300986 122614
rect 301222 122378 301306 122614
rect 301542 122378 336986 122614
rect 337222 122378 337306 122614
rect 337542 122378 372986 122614
rect 373222 122378 373306 122614
rect 373542 122378 408986 122614
rect 409222 122378 409306 122614
rect 409542 122378 444986 122614
rect 445222 122378 445306 122614
rect 445542 122378 480986 122614
rect 481222 122378 481306 122614
rect 481542 122378 516986 122614
rect 517222 122378 517306 122614
rect 517542 122378 552986 122614
rect 553222 122378 553306 122614
rect 553542 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 12986 122294
rect 13222 122058 13306 122294
rect 13542 122058 48986 122294
rect 49222 122058 49306 122294
rect 49542 122058 228986 122294
rect 229222 122058 229306 122294
rect 229542 122058 264986 122294
rect 265222 122058 265306 122294
rect 265542 122058 300986 122294
rect 301222 122058 301306 122294
rect 301542 122058 336986 122294
rect 337222 122058 337306 122294
rect 337542 122058 372986 122294
rect 373222 122058 373306 122294
rect 373542 122058 408986 122294
rect 409222 122058 409306 122294
rect 409542 122058 444986 122294
rect 445222 122058 445306 122294
rect 445542 122058 480986 122294
rect 481222 122058 481306 122294
rect 481542 122058 516986 122294
rect 517222 122058 517306 122294
rect 517542 122058 552986 122294
rect 553222 122058 553306 122294
rect 553542 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 9266 118894
rect 9502 118658 9586 118894
rect 9822 118658 45266 118894
rect 45502 118658 45586 118894
rect 45822 118658 261266 118894
rect 261502 118658 261586 118894
rect 261822 118658 297266 118894
rect 297502 118658 297586 118894
rect 297822 118658 333266 118894
rect 333502 118658 333586 118894
rect 333822 118658 369266 118894
rect 369502 118658 369586 118894
rect 369822 118658 405266 118894
rect 405502 118658 405586 118894
rect 405822 118658 441266 118894
rect 441502 118658 441586 118894
rect 441822 118658 477266 118894
rect 477502 118658 477586 118894
rect 477822 118658 513266 118894
rect 513502 118658 513586 118894
rect 513822 118658 549266 118894
rect 549502 118658 549586 118894
rect 549822 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 9266 118574
rect 9502 118338 9586 118574
rect 9822 118338 45266 118574
rect 45502 118338 45586 118574
rect 45822 118338 261266 118574
rect 261502 118338 261586 118574
rect 261822 118338 297266 118574
rect 297502 118338 297586 118574
rect 297822 118338 333266 118574
rect 333502 118338 333586 118574
rect 333822 118338 369266 118574
rect 369502 118338 369586 118574
rect 369822 118338 405266 118574
rect 405502 118338 405586 118574
rect 405822 118338 441266 118574
rect 441502 118338 441586 118574
rect 441822 118338 477266 118574
rect 477502 118338 477586 118574
rect 477822 118338 513266 118574
rect 513502 118338 513586 118574
rect 513822 118338 549266 118574
rect 549502 118338 549586 118574
rect 549822 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 5546 115174
rect 5782 114938 5866 115174
rect 6102 114938 41546 115174
rect 41782 114938 41866 115174
rect 42102 114938 257546 115174
rect 257782 114938 257866 115174
rect 258102 114938 293546 115174
rect 293782 114938 293866 115174
rect 294102 114938 329546 115174
rect 329782 114938 329866 115174
rect 330102 114938 365546 115174
rect 365782 114938 365866 115174
rect 366102 114938 401546 115174
rect 401782 114938 401866 115174
rect 402102 114938 437546 115174
rect 437782 114938 437866 115174
rect 438102 114938 473546 115174
rect 473782 114938 473866 115174
rect 474102 114938 509546 115174
rect 509782 114938 509866 115174
rect 510102 114938 545546 115174
rect 545782 114938 545866 115174
rect 546102 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 5546 114854
rect 5782 114618 5866 114854
rect 6102 114618 41546 114854
rect 41782 114618 41866 114854
rect 42102 114618 257546 114854
rect 257782 114618 257866 114854
rect 258102 114618 293546 114854
rect 293782 114618 293866 114854
rect 294102 114618 329546 114854
rect 329782 114618 329866 114854
rect 330102 114618 365546 114854
rect 365782 114618 365866 114854
rect 366102 114618 401546 114854
rect 401782 114618 401866 114854
rect 402102 114618 437546 114854
rect 437782 114618 437866 114854
rect 438102 114618 473546 114854
rect 473782 114618 473866 114854
rect 474102 114618 509546 114854
rect 509782 114618 509866 114854
rect 510102 114618 545546 114854
rect 545782 114618 545866 114854
rect 546102 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 1826 111454
rect 2062 111218 2146 111454
rect 2382 111218 37826 111454
rect 38062 111218 38146 111454
rect 38382 111218 64250 111454
rect 64486 111218 94970 111454
rect 95206 111218 125690 111454
rect 125926 111218 156410 111454
rect 156646 111218 187130 111454
rect 187366 111218 217850 111454
rect 218086 111218 253826 111454
rect 254062 111218 254146 111454
rect 254382 111218 289826 111454
rect 290062 111218 290146 111454
rect 290382 111218 325826 111454
rect 326062 111218 326146 111454
rect 326382 111218 361826 111454
rect 362062 111218 362146 111454
rect 362382 111218 397826 111454
rect 398062 111218 398146 111454
rect 398382 111218 433826 111454
rect 434062 111218 434146 111454
rect 434382 111218 469826 111454
rect 470062 111218 470146 111454
rect 470382 111218 505826 111454
rect 506062 111218 506146 111454
rect 506382 111218 541826 111454
rect 542062 111218 542146 111454
rect 542382 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 1826 111134
rect 2062 110898 2146 111134
rect 2382 110898 37826 111134
rect 38062 110898 38146 111134
rect 38382 110898 64250 111134
rect 64486 110898 94970 111134
rect 95206 110898 125690 111134
rect 125926 110898 156410 111134
rect 156646 110898 187130 111134
rect 187366 110898 217850 111134
rect 218086 110898 253826 111134
rect 254062 110898 254146 111134
rect 254382 110898 289826 111134
rect 290062 110898 290146 111134
rect 290382 110898 325826 111134
rect 326062 110898 326146 111134
rect 326382 110898 361826 111134
rect 362062 110898 362146 111134
rect 362382 110898 397826 111134
rect 398062 110898 398146 111134
rect 398382 110898 433826 111134
rect 434062 110898 434146 111134
rect 434382 110898 469826 111134
rect 470062 110898 470146 111134
rect 470382 110898 505826 111134
rect 506062 110898 506146 111134
rect 506382 110898 541826 111134
rect 542062 110898 542146 111134
rect 542382 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 30986 104614
rect 31222 104378 31306 104614
rect 31542 104378 246986 104614
rect 247222 104378 247306 104614
rect 247542 104378 282986 104614
rect 283222 104378 283306 104614
rect 283542 104378 318986 104614
rect 319222 104378 319306 104614
rect 319542 104378 354986 104614
rect 355222 104378 355306 104614
rect 355542 104378 390986 104614
rect 391222 104378 391306 104614
rect 391542 104378 426986 104614
rect 427222 104378 427306 104614
rect 427542 104378 462986 104614
rect 463222 104378 463306 104614
rect 463542 104378 498986 104614
rect 499222 104378 499306 104614
rect 499542 104378 534986 104614
rect 535222 104378 535306 104614
rect 535542 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 30986 104294
rect 31222 104058 31306 104294
rect 31542 104058 246986 104294
rect 247222 104058 247306 104294
rect 247542 104058 282986 104294
rect 283222 104058 283306 104294
rect 283542 104058 318986 104294
rect 319222 104058 319306 104294
rect 319542 104058 354986 104294
rect 355222 104058 355306 104294
rect 355542 104058 390986 104294
rect 391222 104058 391306 104294
rect 391542 104058 426986 104294
rect 427222 104058 427306 104294
rect 427542 104058 462986 104294
rect 463222 104058 463306 104294
rect 463542 104058 498986 104294
rect 499222 104058 499306 104294
rect 499542 104058 534986 104294
rect 535222 104058 535306 104294
rect 535542 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 27266 100894
rect 27502 100658 27586 100894
rect 27822 100658 243266 100894
rect 243502 100658 243586 100894
rect 243822 100658 279266 100894
rect 279502 100658 279586 100894
rect 279822 100658 315266 100894
rect 315502 100658 315586 100894
rect 315822 100658 351266 100894
rect 351502 100658 351586 100894
rect 351822 100658 387266 100894
rect 387502 100658 387586 100894
rect 387822 100658 423266 100894
rect 423502 100658 423586 100894
rect 423822 100658 459266 100894
rect 459502 100658 459586 100894
rect 459822 100658 495266 100894
rect 495502 100658 495586 100894
rect 495822 100658 531266 100894
rect 531502 100658 531586 100894
rect 531822 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 27266 100574
rect 27502 100338 27586 100574
rect 27822 100338 243266 100574
rect 243502 100338 243586 100574
rect 243822 100338 279266 100574
rect 279502 100338 279586 100574
rect 279822 100338 315266 100574
rect 315502 100338 315586 100574
rect 315822 100338 351266 100574
rect 351502 100338 351586 100574
rect 351822 100338 387266 100574
rect 387502 100338 387586 100574
rect 387822 100338 423266 100574
rect 423502 100338 423586 100574
rect 423822 100338 459266 100574
rect 459502 100338 459586 100574
rect 459822 100338 495266 100574
rect 495502 100338 495586 100574
rect 495822 100338 531266 100574
rect 531502 100338 531586 100574
rect 531822 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 23546 97174
rect 23782 96938 23866 97174
rect 24102 96938 239546 97174
rect 239782 96938 239866 97174
rect 240102 96938 275546 97174
rect 275782 96938 275866 97174
rect 276102 96938 311546 97174
rect 311782 96938 311866 97174
rect 312102 96938 347546 97174
rect 347782 96938 347866 97174
rect 348102 96938 383546 97174
rect 383782 96938 383866 97174
rect 384102 96938 419546 97174
rect 419782 96938 419866 97174
rect 420102 96938 455546 97174
rect 455782 96938 455866 97174
rect 456102 96938 491546 97174
rect 491782 96938 491866 97174
rect 492102 96938 527546 97174
rect 527782 96938 527866 97174
rect 528102 96938 563546 97174
rect 563782 96938 563866 97174
rect 564102 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 23546 96854
rect 23782 96618 23866 96854
rect 24102 96618 239546 96854
rect 239782 96618 239866 96854
rect 240102 96618 275546 96854
rect 275782 96618 275866 96854
rect 276102 96618 311546 96854
rect 311782 96618 311866 96854
rect 312102 96618 347546 96854
rect 347782 96618 347866 96854
rect 348102 96618 383546 96854
rect 383782 96618 383866 96854
rect 384102 96618 419546 96854
rect 419782 96618 419866 96854
rect 420102 96618 455546 96854
rect 455782 96618 455866 96854
rect 456102 96618 491546 96854
rect 491782 96618 491866 96854
rect 492102 96618 527546 96854
rect 527782 96618 527866 96854
rect 528102 96618 563546 96854
rect 563782 96618 563866 96854
rect 564102 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 19826 93454
rect 20062 93218 20146 93454
rect 20382 93218 55826 93454
rect 56062 93218 56146 93454
rect 56382 93218 79610 93454
rect 79846 93218 110330 93454
rect 110566 93218 141050 93454
rect 141286 93218 171770 93454
rect 172006 93218 202490 93454
rect 202726 93218 235826 93454
rect 236062 93218 236146 93454
rect 236382 93218 271826 93454
rect 272062 93218 272146 93454
rect 272382 93218 307826 93454
rect 308062 93218 308146 93454
rect 308382 93218 343826 93454
rect 344062 93218 344146 93454
rect 344382 93218 379826 93454
rect 380062 93218 380146 93454
rect 380382 93218 415826 93454
rect 416062 93218 416146 93454
rect 416382 93218 451826 93454
rect 452062 93218 452146 93454
rect 452382 93218 487826 93454
rect 488062 93218 488146 93454
rect 488382 93218 523826 93454
rect 524062 93218 524146 93454
rect 524382 93218 559826 93454
rect 560062 93218 560146 93454
rect 560382 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 19826 93134
rect 20062 92898 20146 93134
rect 20382 92898 55826 93134
rect 56062 92898 56146 93134
rect 56382 92898 79610 93134
rect 79846 92898 110330 93134
rect 110566 92898 141050 93134
rect 141286 92898 171770 93134
rect 172006 92898 202490 93134
rect 202726 92898 235826 93134
rect 236062 92898 236146 93134
rect 236382 92898 271826 93134
rect 272062 92898 272146 93134
rect 272382 92898 307826 93134
rect 308062 92898 308146 93134
rect 308382 92898 343826 93134
rect 344062 92898 344146 93134
rect 344382 92898 379826 93134
rect 380062 92898 380146 93134
rect 380382 92898 415826 93134
rect 416062 92898 416146 93134
rect 416382 92898 451826 93134
rect 452062 92898 452146 93134
rect 452382 92898 487826 93134
rect 488062 92898 488146 93134
rect 488382 92898 523826 93134
rect 524062 92898 524146 93134
rect 524382 92898 559826 93134
rect 560062 92898 560146 93134
rect 560382 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 12986 86614
rect 13222 86378 13306 86614
rect 13542 86378 48986 86614
rect 49222 86378 49306 86614
rect 49542 86378 228986 86614
rect 229222 86378 229306 86614
rect 229542 86378 264986 86614
rect 265222 86378 265306 86614
rect 265542 86378 300986 86614
rect 301222 86378 301306 86614
rect 301542 86378 336986 86614
rect 337222 86378 337306 86614
rect 337542 86378 372986 86614
rect 373222 86378 373306 86614
rect 373542 86378 408986 86614
rect 409222 86378 409306 86614
rect 409542 86378 444986 86614
rect 445222 86378 445306 86614
rect 445542 86378 480986 86614
rect 481222 86378 481306 86614
rect 481542 86378 516986 86614
rect 517222 86378 517306 86614
rect 517542 86378 552986 86614
rect 553222 86378 553306 86614
rect 553542 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 12986 86294
rect 13222 86058 13306 86294
rect 13542 86058 48986 86294
rect 49222 86058 49306 86294
rect 49542 86058 228986 86294
rect 229222 86058 229306 86294
rect 229542 86058 264986 86294
rect 265222 86058 265306 86294
rect 265542 86058 300986 86294
rect 301222 86058 301306 86294
rect 301542 86058 336986 86294
rect 337222 86058 337306 86294
rect 337542 86058 372986 86294
rect 373222 86058 373306 86294
rect 373542 86058 408986 86294
rect 409222 86058 409306 86294
rect 409542 86058 444986 86294
rect 445222 86058 445306 86294
rect 445542 86058 480986 86294
rect 481222 86058 481306 86294
rect 481542 86058 516986 86294
rect 517222 86058 517306 86294
rect 517542 86058 552986 86294
rect 553222 86058 553306 86294
rect 553542 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 9266 82894
rect 9502 82658 9586 82894
rect 9822 82658 45266 82894
rect 45502 82658 45586 82894
rect 45822 82658 261266 82894
rect 261502 82658 261586 82894
rect 261822 82658 297266 82894
rect 297502 82658 297586 82894
rect 297822 82658 333266 82894
rect 333502 82658 333586 82894
rect 333822 82658 369266 82894
rect 369502 82658 369586 82894
rect 369822 82658 405266 82894
rect 405502 82658 405586 82894
rect 405822 82658 441266 82894
rect 441502 82658 441586 82894
rect 441822 82658 477266 82894
rect 477502 82658 477586 82894
rect 477822 82658 513266 82894
rect 513502 82658 513586 82894
rect 513822 82658 549266 82894
rect 549502 82658 549586 82894
rect 549822 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 9266 82574
rect 9502 82338 9586 82574
rect 9822 82338 45266 82574
rect 45502 82338 45586 82574
rect 45822 82338 261266 82574
rect 261502 82338 261586 82574
rect 261822 82338 297266 82574
rect 297502 82338 297586 82574
rect 297822 82338 333266 82574
rect 333502 82338 333586 82574
rect 333822 82338 369266 82574
rect 369502 82338 369586 82574
rect 369822 82338 405266 82574
rect 405502 82338 405586 82574
rect 405822 82338 441266 82574
rect 441502 82338 441586 82574
rect 441822 82338 477266 82574
rect 477502 82338 477586 82574
rect 477822 82338 513266 82574
rect 513502 82338 513586 82574
rect 513822 82338 549266 82574
rect 549502 82338 549586 82574
rect 549822 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 5546 79174
rect 5782 78938 5866 79174
rect 6102 78938 41546 79174
rect 41782 78938 41866 79174
rect 42102 78938 257546 79174
rect 257782 78938 257866 79174
rect 258102 78938 293546 79174
rect 293782 78938 293866 79174
rect 294102 78938 329546 79174
rect 329782 78938 329866 79174
rect 330102 78938 365546 79174
rect 365782 78938 365866 79174
rect 366102 78938 401546 79174
rect 401782 78938 401866 79174
rect 402102 78938 437546 79174
rect 437782 78938 437866 79174
rect 438102 78938 473546 79174
rect 473782 78938 473866 79174
rect 474102 78938 509546 79174
rect 509782 78938 509866 79174
rect 510102 78938 545546 79174
rect 545782 78938 545866 79174
rect 546102 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 5546 78854
rect 5782 78618 5866 78854
rect 6102 78618 41546 78854
rect 41782 78618 41866 78854
rect 42102 78618 257546 78854
rect 257782 78618 257866 78854
rect 258102 78618 293546 78854
rect 293782 78618 293866 78854
rect 294102 78618 329546 78854
rect 329782 78618 329866 78854
rect 330102 78618 365546 78854
rect 365782 78618 365866 78854
rect 366102 78618 401546 78854
rect 401782 78618 401866 78854
rect 402102 78618 437546 78854
rect 437782 78618 437866 78854
rect 438102 78618 473546 78854
rect 473782 78618 473866 78854
rect 474102 78618 509546 78854
rect 509782 78618 509866 78854
rect 510102 78618 545546 78854
rect 545782 78618 545866 78854
rect 546102 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 1826 75454
rect 2062 75218 2146 75454
rect 2382 75218 37826 75454
rect 38062 75218 38146 75454
rect 38382 75218 64250 75454
rect 64486 75218 94970 75454
rect 95206 75218 125690 75454
rect 125926 75218 156410 75454
rect 156646 75218 187130 75454
rect 187366 75218 217850 75454
rect 218086 75218 253826 75454
rect 254062 75218 254146 75454
rect 254382 75218 289826 75454
rect 290062 75218 290146 75454
rect 290382 75218 325826 75454
rect 326062 75218 326146 75454
rect 326382 75218 361826 75454
rect 362062 75218 362146 75454
rect 362382 75218 397826 75454
rect 398062 75218 398146 75454
rect 398382 75218 433826 75454
rect 434062 75218 434146 75454
rect 434382 75218 469826 75454
rect 470062 75218 470146 75454
rect 470382 75218 505826 75454
rect 506062 75218 506146 75454
rect 506382 75218 541826 75454
rect 542062 75218 542146 75454
rect 542382 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 1826 75134
rect 2062 74898 2146 75134
rect 2382 74898 37826 75134
rect 38062 74898 38146 75134
rect 38382 74898 64250 75134
rect 64486 74898 94970 75134
rect 95206 74898 125690 75134
rect 125926 74898 156410 75134
rect 156646 74898 187130 75134
rect 187366 74898 217850 75134
rect 218086 74898 253826 75134
rect 254062 74898 254146 75134
rect 254382 74898 289826 75134
rect 290062 74898 290146 75134
rect 290382 74898 325826 75134
rect 326062 74898 326146 75134
rect 326382 74898 361826 75134
rect 362062 74898 362146 75134
rect 362382 74898 397826 75134
rect 398062 74898 398146 75134
rect 398382 74898 433826 75134
rect 434062 74898 434146 75134
rect 434382 74898 469826 75134
rect 470062 74898 470146 75134
rect 470382 74898 505826 75134
rect 506062 74898 506146 75134
rect 506382 74898 541826 75134
rect 542062 74898 542146 75134
rect 542382 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 30986 68614
rect 31222 68378 31306 68614
rect 31542 68378 246986 68614
rect 247222 68378 247306 68614
rect 247542 68378 282986 68614
rect 283222 68378 283306 68614
rect 283542 68378 318986 68614
rect 319222 68378 319306 68614
rect 319542 68378 354986 68614
rect 355222 68378 355306 68614
rect 355542 68378 390986 68614
rect 391222 68378 391306 68614
rect 391542 68378 426986 68614
rect 427222 68378 427306 68614
rect 427542 68378 462986 68614
rect 463222 68378 463306 68614
rect 463542 68378 498986 68614
rect 499222 68378 499306 68614
rect 499542 68378 534986 68614
rect 535222 68378 535306 68614
rect 535542 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 30986 68294
rect 31222 68058 31306 68294
rect 31542 68058 246986 68294
rect 247222 68058 247306 68294
rect 247542 68058 282986 68294
rect 283222 68058 283306 68294
rect 283542 68058 318986 68294
rect 319222 68058 319306 68294
rect 319542 68058 354986 68294
rect 355222 68058 355306 68294
rect 355542 68058 390986 68294
rect 391222 68058 391306 68294
rect 391542 68058 426986 68294
rect 427222 68058 427306 68294
rect 427542 68058 462986 68294
rect 463222 68058 463306 68294
rect 463542 68058 498986 68294
rect 499222 68058 499306 68294
rect 499542 68058 534986 68294
rect 535222 68058 535306 68294
rect 535542 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 27266 64894
rect 27502 64658 27586 64894
rect 27822 64658 243266 64894
rect 243502 64658 243586 64894
rect 243822 64658 279266 64894
rect 279502 64658 279586 64894
rect 279822 64658 315266 64894
rect 315502 64658 315586 64894
rect 315822 64658 351266 64894
rect 351502 64658 351586 64894
rect 351822 64658 387266 64894
rect 387502 64658 387586 64894
rect 387822 64658 423266 64894
rect 423502 64658 423586 64894
rect 423822 64658 459266 64894
rect 459502 64658 459586 64894
rect 459822 64658 495266 64894
rect 495502 64658 495586 64894
rect 495822 64658 531266 64894
rect 531502 64658 531586 64894
rect 531822 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 27266 64574
rect 27502 64338 27586 64574
rect 27822 64338 243266 64574
rect 243502 64338 243586 64574
rect 243822 64338 279266 64574
rect 279502 64338 279586 64574
rect 279822 64338 315266 64574
rect 315502 64338 315586 64574
rect 315822 64338 351266 64574
rect 351502 64338 351586 64574
rect 351822 64338 387266 64574
rect 387502 64338 387586 64574
rect 387822 64338 423266 64574
rect 423502 64338 423586 64574
rect 423822 64338 459266 64574
rect 459502 64338 459586 64574
rect 459822 64338 495266 64574
rect 495502 64338 495586 64574
rect 495822 64338 531266 64574
rect 531502 64338 531586 64574
rect 531822 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 23546 61174
rect 23782 60938 23866 61174
rect 24102 60938 239546 61174
rect 239782 60938 239866 61174
rect 240102 60938 275546 61174
rect 275782 60938 275866 61174
rect 276102 60938 311546 61174
rect 311782 60938 311866 61174
rect 312102 60938 347546 61174
rect 347782 60938 347866 61174
rect 348102 60938 383546 61174
rect 383782 60938 383866 61174
rect 384102 60938 419546 61174
rect 419782 60938 419866 61174
rect 420102 60938 455546 61174
rect 455782 60938 455866 61174
rect 456102 60938 491546 61174
rect 491782 60938 491866 61174
rect 492102 60938 527546 61174
rect 527782 60938 527866 61174
rect 528102 60938 563546 61174
rect 563782 60938 563866 61174
rect 564102 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 23546 60854
rect 23782 60618 23866 60854
rect 24102 60618 239546 60854
rect 239782 60618 239866 60854
rect 240102 60618 275546 60854
rect 275782 60618 275866 60854
rect 276102 60618 311546 60854
rect 311782 60618 311866 60854
rect 312102 60618 347546 60854
rect 347782 60618 347866 60854
rect 348102 60618 383546 60854
rect 383782 60618 383866 60854
rect 384102 60618 419546 60854
rect 419782 60618 419866 60854
rect 420102 60618 455546 60854
rect 455782 60618 455866 60854
rect 456102 60618 491546 60854
rect 491782 60618 491866 60854
rect 492102 60618 527546 60854
rect 527782 60618 527866 60854
rect 528102 60618 563546 60854
rect 563782 60618 563866 60854
rect 564102 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 19826 57454
rect 20062 57218 20146 57454
rect 20382 57218 55826 57454
rect 56062 57218 56146 57454
rect 56382 57218 91826 57454
rect 92062 57218 92146 57454
rect 92382 57218 127826 57454
rect 128062 57218 128146 57454
rect 128382 57218 163826 57454
rect 164062 57218 164146 57454
rect 164382 57218 199826 57454
rect 200062 57218 200146 57454
rect 200382 57218 235826 57454
rect 236062 57218 236146 57454
rect 236382 57218 271826 57454
rect 272062 57218 272146 57454
rect 272382 57218 307826 57454
rect 308062 57218 308146 57454
rect 308382 57218 343826 57454
rect 344062 57218 344146 57454
rect 344382 57218 379826 57454
rect 380062 57218 380146 57454
rect 380382 57218 415826 57454
rect 416062 57218 416146 57454
rect 416382 57218 451826 57454
rect 452062 57218 452146 57454
rect 452382 57218 487826 57454
rect 488062 57218 488146 57454
rect 488382 57218 523826 57454
rect 524062 57218 524146 57454
rect 524382 57218 559826 57454
rect 560062 57218 560146 57454
rect 560382 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 19826 57134
rect 20062 56898 20146 57134
rect 20382 56898 55826 57134
rect 56062 56898 56146 57134
rect 56382 56898 91826 57134
rect 92062 56898 92146 57134
rect 92382 56898 127826 57134
rect 128062 56898 128146 57134
rect 128382 56898 163826 57134
rect 164062 56898 164146 57134
rect 164382 56898 199826 57134
rect 200062 56898 200146 57134
rect 200382 56898 235826 57134
rect 236062 56898 236146 57134
rect 236382 56898 271826 57134
rect 272062 56898 272146 57134
rect 272382 56898 307826 57134
rect 308062 56898 308146 57134
rect 308382 56898 343826 57134
rect 344062 56898 344146 57134
rect 344382 56898 379826 57134
rect 380062 56898 380146 57134
rect 380382 56898 415826 57134
rect 416062 56898 416146 57134
rect 416382 56898 451826 57134
rect 452062 56898 452146 57134
rect 452382 56898 487826 57134
rect 488062 56898 488146 57134
rect 488382 56898 523826 57134
rect 524062 56898 524146 57134
rect 524382 56898 559826 57134
rect 560062 56898 560146 57134
rect 560382 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 12986 50614
rect 13222 50378 13306 50614
rect 13542 50378 48986 50614
rect 49222 50378 49306 50614
rect 49542 50378 84986 50614
rect 85222 50378 85306 50614
rect 85542 50378 120986 50614
rect 121222 50378 121306 50614
rect 121542 50378 156986 50614
rect 157222 50378 157306 50614
rect 157542 50378 192986 50614
rect 193222 50378 193306 50614
rect 193542 50378 228986 50614
rect 229222 50378 229306 50614
rect 229542 50378 264986 50614
rect 265222 50378 265306 50614
rect 265542 50378 300986 50614
rect 301222 50378 301306 50614
rect 301542 50378 336986 50614
rect 337222 50378 337306 50614
rect 337542 50378 372986 50614
rect 373222 50378 373306 50614
rect 373542 50378 408986 50614
rect 409222 50378 409306 50614
rect 409542 50378 444986 50614
rect 445222 50378 445306 50614
rect 445542 50378 480986 50614
rect 481222 50378 481306 50614
rect 481542 50378 516986 50614
rect 517222 50378 517306 50614
rect 517542 50378 552986 50614
rect 553222 50378 553306 50614
rect 553542 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 12986 50294
rect 13222 50058 13306 50294
rect 13542 50058 48986 50294
rect 49222 50058 49306 50294
rect 49542 50058 84986 50294
rect 85222 50058 85306 50294
rect 85542 50058 120986 50294
rect 121222 50058 121306 50294
rect 121542 50058 156986 50294
rect 157222 50058 157306 50294
rect 157542 50058 192986 50294
rect 193222 50058 193306 50294
rect 193542 50058 228986 50294
rect 229222 50058 229306 50294
rect 229542 50058 264986 50294
rect 265222 50058 265306 50294
rect 265542 50058 300986 50294
rect 301222 50058 301306 50294
rect 301542 50058 336986 50294
rect 337222 50058 337306 50294
rect 337542 50058 372986 50294
rect 373222 50058 373306 50294
rect 373542 50058 408986 50294
rect 409222 50058 409306 50294
rect 409542 50058 444986 50294
rect 445222 50058 445306 50294
rect 445542 50058 480986 50294
rect 481222 50058 481306 50294
rect 481542 50058 516986 50294
rect 517222 50058 517306 50294
rect 517542 50058 552986 50294
rect 553222 50058 553306 50294
rect 553542 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 9266 46894
rect 9502 46658 9586 46894
rect 9822 46658 45266 46894
rect 45502 46658 45586 46894
rect 45822 46658 81266 46894
rect 81502 46658 81586 46894
rect 81822 46658 117266 46894
rect 117502 46658 117586 46894
rect 117822 46658 153266 46894
rect 153502 46658 153586 46894
rect 153822 46658 189266 46894
rect 189502 46658 189586 46894
rect 189822 46658 225266 46894
rect 225502 46658 225586 46894
rect 225822 46658 261266 46894
rect 261502 46658 261586 46894
rect 261822 46658 297266 46894
rect 297502 46658 297586 46894
rect 297822 46658 333266 46894
rect 333502 46658 333586 46894
rect 333822 46658 369266 46894
rect 369502 46658 369586 46894
rect 369822 46658 405266 46894
rect 405502 46658 405586 46894
rect 405822 46658 441266 46894
rect 441502 46658 441586 46894
rect 441822 46658 477266 46894
rect 477502 46658 477586 46894
rect 477822 46658 513266 46894
rect 513502 46658 513586 46894
rect 513822 46658 549266 46894
rect 549502 46658 549586 46894
rect 549822 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 9266 46574
rect 9502 46338 9586 46574
rect 9822 46338 45266 46574
rect 45502 46338 45586 46574
rect 45822 46338 81266 46574
rect 81502 46338 81586 46574
rect 81822 46338 117266 46574
rect 117502 46338 117586 46574
rect 117822 46338 153266 46574
rect 153502 46338 153586 46574
rect 153822 46338 189266 46574
rect 189502 46338 189586 46574
rect 189822 46338 225266 46574
rect 225502 46338 225586 46574
rect 225822 46338 261266 46574
rect 261502 46338 261586 46574
rect 261822 46338 297266 46574
rect 297502 46338 297586 46574
rect 297822 46338 333266 46574
rect 333502 46338 333586 46574
rect 333822 46338 369266 46574
rect 369502 46338 369586 46574
rect 369822 46338 405266 46574
rect 405502 46338 405586 46574
rect 405822 46338 441266 46574
rect 441502 46338 441586 46574
rect 441822 46338 477266 46574
rect 477502 46338 477586 46574
rect 477822 46338 513266 46574
rect 513502 46338 513586 46574
rect 513822 46338 549266 46574
rect 549502 46338 549586 46574
rect 549822 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 5546 43174
rect 5782 42938 5866 43174
rect 6102 42938 41546 43174
rect 41782 42938 41866 43174
rect 42102 42938 77546 43174
rect 77782 42938 77866 43174
rect 78102 42938 113546 43174
rect 113782 42938 113866 43174
rect 114102 42938 149546 43174
rect 149782 42938 149866 43174
rect 150102 42938 185546 43174
rect 185782 42938 185866 43174
rect 186102 42938 221546 43174
rect 221782 42938 221866 43174
rect 222102 42938 257546 43174
rect 257782 42938 257866 43174
rect 258102 42938 293546 43174
rect 293782 42938 293866 43174
rect 294102 42938 329546 43174
rect 329782 42938 329866 43174
rect 330102 42938 365546 43174
rect 365782 42938 365866 43174
rect 366102 42938 401546 43174
rect 401782 42938 401866 43174
rect 402102 42938 437546 43174
rect 437782 42938 437866 43174
rect 438102 42938 473546 43174
rect 473782 42938 473866 43174
rect 474102 42938 509546 43174
rect 509782 42938 509866 43174
rect 510102 42938 545546 43174
rect 545782 42938 545866 43174
rect 546102 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 5546 42854
rect 5782 42618 5866 42854
rect 6102 42618 41546 42854
rect 41782 42618 41866 42854
rect 42102 42618 77546 42854
rect 77782 42618 77866 42854
rect 78102 42618 113546 42854
rect 113782 42618 113866 42854
rect 114102 42618 149546 42854
rect 149782 42618 149866 42854
rect 150102 42618 185546 42854
rect 185782 42618 185866 42854
rect 186102 42618 221546 42854
rect 221782 42618 221866 42854
rect 222102 42618 257546 42854
rect 257782 42618 257866 42854
rect 258102 42618 293546 42854
rect 293782 42618 293866 42854
rect 294102 42618 329546 42854
rect 329782 42618 329866 42854
rect 330102 42618 365546 42854
rect 365782 42618 365866 42854
rect 366102 42618 401546 42854
rect 401782 42618 401866 42854
rect 402102 42618 437546 42854
rect 437782 42618 437866 42854
rect 438102 42618 473546 42854
rect 473782 42618 473866 42854
rect 474102 42618 509546 42854
rect 509782 42618 509866 42854
rect 510102 42618 545546 42854
rect 545782 42618 545866 42854
rect 546102 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 1826 39454
rect 2062 39218 2146 39454
rect 2382 39218 37826 39454
rect 38062 39218 38146 39454
rect 38382 39218 73826 39454
rect 74062 39218 74146 39454
rect 74382 39218 109826 39454
rect 110062 39218 110146 39454
rect 110382 39218 145826 39454
rect 146062 39218 146146 39454
rect 146382 39218 181826 39454
rect 182062 39218 182146 39454
rect 182382 39218 217826 39454
rect 218062 39218 218146 39454
rect 218382 39218 253826 39454
rect 254062 39218 254146 39454
rect 254382 39218 289826 39454
rect 290062 39218 290146 39454
rect 290382 39218 325826 39454
rect 326062 39218 326146 39454
rect 326382 39218 361826 39454
rect 362062 39218 362146 39454
rect 362382 39218 397826 39454
rect 398062 39218 398146 39454
rect 398382 39218 433826 39454
rect 434062 39218 434146 39454
rect 434382 39218 469826 39454
rect 470062 39218 470146 39454
rect 470382 39218 505826 39454
rect 506062 39218 506146 39454
rect 506382 39218 541826 39454
rect 542062 39218 542146 39454
rect 542382 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 1826 39134
rect 2062 38898 2146 39134
rect 2382 38898 37826 39134
rect 38062 38898 38146 39134
rect 38382 38898 73826 39134
rect 74062 38898 74146 39134
rect 74382 38898 109826 39134
rect 110062 38898 110146 39134
rect 110382 38898 145826 39134
rect 146062 38898 146146 39134
rect 146382 38898 181826 39134
rect 182062 38898 182146 39134
rect 182382 38898 217826 39134
rect 218062 38898 218146 39134
rect 218382 38898 253826 39134
rect 254062 38898 254146 39134
rect 254382 38898 289826 39134
rect 290062 38898 290146 39134
rect 290382 38898 325826 39134
rect 326062 38898 326146 39134
rect 326382 38898 361826 39134
rect 362062 38898 362146 39134
rect 362382 38898 397826 39134
rect 398062 38898 398146 39134
rect 398382 38898 433826 39134
rect 434062 38898 434146 39134
rect 434382 38898 469826 39134
rect 470062 38898 470146 39134
rect 470382 38898 505826 39134
rect 506062 38898 506146 39134
rect 506382 38898 541826 39134
rect 542062 38898 542146 39134
rect 542382 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 30986 32614
rect 31222 32378 31306 32614
rect 31542 32378 66986 32614
rect 67222 32378 67306 32614
rect 67542 32378 102986 32614
rect 103222 32378 103306 32614
rect 103542 32378 138986 32614
rect 139222 32378 139306 32614
rect 139542 32378 174986 32614
rect 175222 32378 175306 32614
rect 175542 32378 210986 32614
rect 211222 32378 211306 32614
rect 211542 32378 246986 32614
rect 247222 32378 247306 32614
rect 247542 32378 282986 32614
rect 283222 32378 283306 32614
rect 283542 32378 318986 32614
rect 319222 32378 319306 32614
rect 319542 32378 354986 32614
rect 355222 32378 355306 32614
rect 355542 32378 390986 32614
rect 391222 32378 391306 32614
rect 391542 32378 426986 32614
rect 427222 32378 427306 32614
rect 427542 32378 462986 32614
rect 463222 32378 463306 32614
rect 463542 32378 498986 32614
rect 499222 32378 499306 32614
rect 499542 32378 534986 32614
rect 535222 32378 535306 32614
rect 535542 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 30986 32294
rect 31222 32058 31306 32294
rect 31542 32058 66986 32294
rect 67222 32058 67306 32294
rect 67542 32058 102986 32294
rect 103222 32058 103306 32294
rect 103542 32058 138986 32294
rect 139222 32058 139306 32294
rect 139542 32058 174986 32294
rect 175222 32058 175306 32294
rect 175542 32058 210986 32294
rect 211222 32058 211306 32294
rect 211542 32058 246986 32294
rect 247222 32058 247306 32294
rect 247542 32058 282986 32294
rect 283222 32058 283306 32294
rect 283542 32058 318986 32294
rect 319222 32058 319306 32294
rect 319542 32058 354986 32294
rect 355222 32058 355306 32294
rect 355542 32058 390986 32294
rect 391222 32058 391306 32294
rect 391542 32058 426986 32294
rect 427222 32058 427306 32294
rect 427542 32058 462986 32294
rect 463222 32058 463306 32294
rect 463542 32058 498986 32294
rect 499222 32058 499306 32294
rect 499542 32058 534986 32294
rect 535222 32058 535306 32294
rect 535542 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 27266 28894
rect 27502 28658 27586 28894
rect 27822 28658 63266 28894
rect 63502 28658 63586 28894
rect 63822 28658 99266 28894
rect 99502 28658 99586 28894
rect 99822 28658 135266 28894
rect 135502 28658 135586 28894
rect 135822 28658 171266 28894
rect 171502 28658 171586 28894
rect 171822 28658 207266 28894
rect 207502 28658 207586 28894
rect 207822 28658 243266 28894
rect 243502 28658 243586 28894
rect 243822 28658 279266 28894
rect 279502 28658 279586 28894
rect 279822 28658 315266 28894
rect 315502 28658 315586 28894
rect 315822 28658 351266 28894
rect 351502 28658 351586 28894
rect 351822 28658 387266 28894
rect 387502 28658 387586 28894
rect 387822 28658 423266 28894
rect 423502 28658 423586 28894
rect 423822 28658 459266 28894
rect 459502 28658 459586 28894
rect 459822 28658 495266 28894
rect 495502 28658 495586 28894
rect 495822 28658 531266 28894
rect 531502 28658 531586 28894
rect 531822 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 27266 28574
rect 27502 28338 27586 28574
rect 27822 28338 63266 28574
rect 63502 28338 63586 28574
rect 63822 28338 99266 28574
rect 99502 28338 99586 28574
rect 99822 28338 135266 28574
rect 135502 28338 135586 28574
rect 135822 28338 171266 28574
rect 171502 28338 171586 28574
rect 171822 28338 207266 28574
rect 207502 28338 207586 28574
rect 207822 28338 243266 28574
rect 243502 28338 243586 28574
rect 243822 28338 279266 28574
rect 279502 28338 279586 28574
rect 279822 28338 315266 28574
rect 315502 28338 315586 28574
rect 315822 28338 351266 28574
rect 351502 28338 351586 28574
rect 351822 28338 387266 28574
rect 387502 28338 387586 28574
rect 387822 28338 423266 28574
rect 423502 28338 423586 28574
rect 423822 28338 459266 28574
rect 459502 28338 459586 28574
rect 459822 28338 495266 28574
rect 495502 28338 495586 28574
rect 495822 28338 531266 28574
rect 531502 28338 531586 28574
rect 531822 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 23546 25174
rect 23782 24938 23866 25174
rect 24102 24938 59546 25174
rect 59782 24938 59866 25174
rect 60102 24938 95546 25174
rect 95782 24938 95866 25174
rect 96102 24938 131546 25174
rect 131782 24938 131866 25174
rect 132102 24938 167546 25174
rect 167782 24938 167866 25174
rect 168102 24938 203546 25174
rect 203782 24938 203866 25174
rect 204102 24938 239546 25174
rect 239782 24938 239866 25174
rect 240102 24938 275546 25174
rect 275782 24938 275866 25174
rect 276102 24938 311546 25174
rect 311782 24938 311866 25174
rect 312102 24938 347546 25174
rect 347782 24938 347866 25174
rect 348102 24938 383546 25174
rect 383782 24938 383866 25174
rect 384102 24938 419546 25174
rect 419782 24938 419866 25174
rect 420102 24938 455546 25174
rect 455782 24938 455866 25174
rect 456102 24938 491546 25174
rect 491782 24938 491866 25174
rect 492102 24938 527546 25174
rect 527782 24938 527866 25174
rect 528102 24938 563546 25174
rect 563782 24938 563866 25174
rect 564102 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 23546 24854
rect 23782 24618 23866 24854
rect 24102 24618 59546 24854
rect 59782 24618 59866 24854
rect 60102 24618 95546 24854
rect 95782 24618 95866 24854
rect 96102 24618 131546 24854
rect 131782 24618 131866 24854
rect 132102 24618 167546 24854
rect 167782 24618 167866 24854
rect 168102 24618 203546 24854
rect 203782 24618 203866 24854
rect 204102 24618 239546 24854
rect 239782 24618 239866 24854
rect 240102 24618 275546 24854
rect 275782 24618 275866 24854
rect 276102 24618 311546 24854
rect 311782 24618 311866 24854
rect 312102 24618 347546 24854
rect 347782 24618 347866 24854
rect 348102 24618 383546 24854
rect 383782 24618 383866 24854
rect 384102 24618 419546 24854
rect 419782 24618 419866 24854
rect 420102 24618 455546 24854
rect 455782 24618 455866 24854
rect 456102 24618 491546 24854
rect 491782 24618 491866 24854
rect 492102 24618 527546 24854
rect 527782 24618 527866 24854
rect 528102 24618 563546 24854
rect 563782 24618 563866 24854
rect 564102 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 19826 21454
rect 20062 21218 20146 21454
rect 20382 21218 55826 21454
rect 56062 21218 56146 21454
rect 56382 21218 91826 21454
rect 92062 21218 92146 21454
rect 92382 21218 127826 21454
rect 128062 21218 128146 21454
rect 128382 21218 163826 21454
rect 164062 21218 164146 21454
rect 164382 21218 199826 21454
rect 200062 21218 200146 21454
rect 200382 21218 235826 21454
rect 236062 21218 236146 21454
rect 236382 21218 271826 21454
rect 272062 21218 272146 21454
rect 272382 21218 307826 21454
rect 308062 21218 308146 21454
rect 308382 21218 343826 21454
rect 344062 21218 344146 21454
rect 344382 21218 379826 21454
rect 380062 21218 380146 21454
rect 380382 21218 415826 21454
rect 416062 21218 416146 21454
rect 416382 21218 451826 21454
rect 452062 21218 452146 21454
rect 452382 21218 487826 21454
rect 488062 21218 488146 21454
rect 488382 21218 523826 21454
rect 524062 21218 524146 21454
rect 524382 21218 559826 21454
rect 560062 21218 560146 21454
rect 560382 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 19826 21134
rect 20062 20898 20146 21134
rect 20382 20898 55826 21134
rect 56062 20898 56146 21134
rect 56382 20898 91826 21134
rect 92062 20898 92146 21134
rect 92382 20898 127826 21134
rect 128062 20898 128146 21134
rect 128382 20898 163826 21134
rect 164062 20898 164146 21134
rect 164382 20898 199826 21134
rect 200062 20898 200146 21134
rect 200382 20898 235826 21134
rect 236062 20898 236146 21134
rect 236382 20898 271826 21134
rect 272062 20898 272146 21134
rect 272382 20898 307826 21134
rect 308062 20898 308146 21134
rect 308382 20898 343826 21134
rect 344062 20898 344146 21134
rect 344382 20898 379826 21134
rect 380062 20898 380146 21134
rect 380382 20898 415826 21134
rect 416062 20898 416146 21134
rect 416382 20898 451826 21134
rect 452062 20898 452146 21134
rect 452382 20898 487826 21134
rect 488062 20898 488146 21134
rect 488382 20898 523826 21134
rect 524062 20898 524146 21134
rect 524382 20898 559826 21134
rect 560062 20898 560146 21134
rect 560382 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 12986 14614
rect 13222 14378 13306 14614
rect 13542 14378 48986 14614
rect 49222 14378 49306 14614
rect 49542 14378 84986 14614
rect 85222 14378 85306 14614
rect 85542 14378 120986 14614
rect 121222 14378 121306 14614
rect 121542 14378 156986 14614
rect 157222 14378 157306 14614
rect 157542 14378 192986 14614
rect 193222 14378 193306 14614
rect 193542 14378 228986 14614
rect 229222 14378 229306 14614
rect 229542 14378 264986 14614
rect 265222 14378 265306 14614
rect 265542 14378 300986 14614
rect 301222 14378 301306 14614
rect 301542 14378 336986 14614
rect 337222 14378 337306 14614
rect 337542 14378 372986 14614
rect 373222 14378 373306 14614
rect 373542 14378 408986 14614
rect 409222 14378 409306 14614
rect 409542 14378 444986 14614
rect 445222 14378 445306 14614
rect 445542 14378 480986 14614
rect 481222 14378 481306 14614
rect 481542 14378 516986 14614
rect 517222 14378 517306 14614
rect 517542 14378 552986 14614
rect 553222 14378 553306 14614
rect 553542 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 12986 14294
rect 13222 14058 13306 14294
rect 13542 14058 48986 14294
rect 49222 14058 49306 14294
rect 49542 14058 84986 14294
rect 85222 14058 85306 14294
rect 85542 14058 120986 14294
rect 121222 14058 121306 14294
rect 121542 14058 156986 14294
rect 157222 14058 157306 14294
rect 157542 14058 192986 14294
rect 193222 14058 193306 14294
rect 193542 14058 228986 14294
rect 229222 14058 229306 14294
rect 229542 14058 264986 14294
rect 265222 14058 265306 14294
rect 265542 14058 300986 14294
rect 301222 14058 301306 14294
rect 301542 14058 336986 14294
rect 337222 14058 337306 14294
rect 337542 14058 372986 14294
rect 373222 14058 373306 14294
rect 373542 14058 408986 14294
rect 409222 14058 409306 14294
rect 409542 14058 444986 14294
rect 445222 14058 445306 14294
rect 445542 14058 480986 14294
rect 481222 14058 481306 14294
rect 481542 14058 516986 14294
rect 517222 14058 517306 14294
rect 517542 14058 552986 14294
rect 553222 14058 553306 14294
rect 553542 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 9266 10894
rect 9502 10658 9586 10894
rect 9822 10658 45266 10894
rect 45502 10658 45586 10894
rect 45822 10658 81266 10894
rect 81502 10658 81586 10894
rect 81822 10658 117266 10894
rect 117502 10658 117586 10894
rect 117822 10658 153266 10894
rect 153502 10658 153586 10894
rect 153822 10658 189266 10894
rect 189502 10658 189586 10894
rect 189822 10658 225266 10894
rect 225502 10658 225586 10894
rect 225822 10658 261266 10894
rect 261502 10658 261586 10894
rect 261822 10658 297266 10894
rect 297502 10658 297586 10894
rect 297822 10658 333266 10894
rect 333502 10658 333586 10894
rect 333822 10658 369266 10894
rect 369502 10658 369586 10894
rect 369822 10658 405266 10894
rect 405502 10658 405586 10894
rect 405822 10658 441266 10894
rect 441502 10658 441586 10894
rect 441822 10658 477266 10894
rect 477502 10658 477586 10894
rect 477822 10658 513266 10894
rect 513502 10658 513586 10894
rect 513822 10658 549266 10894
rect 549502 10658 549586 10894
rect 549822 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 9266 10574
rect 9502 10338 9586 10574
rect 9822 10338 45266 10574
rect 45502 10338 45586 10574
rect 45822 10338 81266 10574
rect 81502 10338 81586 10574
rect 81822 10338 117266 10574
rect 117502 10338 117586 10574
rect 117822 10338 153266 10574
rect 153502 10338 153586 10574
rect 153822 10338 189266 10574
rect 189502 10338 189586 10574
rect 189822 10338 225266 10574
rect 225502 10338 225586 10574
rect 225822 10338 261266 10574
rect 261502 10338 261586 10574
rect 261822 10338 297266 10574
rect 297502 10338 297586 10574
rect 297822 10338 333266 10574
rect 333502 10338 333586 10574
rect 333822 10338 369266 10574
rect 369502 10338 369586 10574
rect 369822 10338 405266 10574
rect 405502 10338 405586 10574
rect 405822 10338 441266 10574
rect 441502 10338 441586 10574
rect 441822 10338 477266 10574
rect 477502 10338 477586 10574
rect 477822 10338 513266 10574
rect 513502 10338 513586 10574
rect 513822 10338 549266 10574
rect 549502 10338 549586 10574
rect 549822 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 5546 7174
rect 5782 6938 5866 7174
rect 6102 6938 41546 7174
rect 41782 6938 41866 7174
rect 42102 6938 77546 7174
rect 77782 6938 77866 7174
rect 78102 6938 113546 7174
rect 113782 6938 113866 7174
rect 114102 6938 149546 7174
rect 149782 6938 149866 7174
rect 150102 6938 185546 7174
rect 185782 6938 185866 7174
rect 186102 6938 221546 7174
rect 221782 6938 221866 7174
rect 222102 6938 257546 7174
rect 257782 6938 257866 7174
rect 258102 6938 293546 7174
rect 293782 6938 293866 7174
rect 294102 6938 329546 7174
rect 329782 6938 329866 7174
rect 330102 6938 365546 7174
rect 365782 6938 365866 7174
rect 366102 6938 401546 7174
rect 401782 6938 401866 7174
rect 402102 6938 437546 7174
rect 437782 6938 437866 7174
rect 438102 6938 473546 7174
rect 473782 6938 473866 7174
rect 474102 6938 509546 7174
rect 509782 6938 509866 7174
rect 510102 6938 545546 7174
rect 545782 6938 545866 7174
rect 546102 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 5546 6854
rect 5782 6618 5866 6854
rect 6102 6618 41546 6854
rect 41782 6618 41866 6854
rect 42102 6618 77546 6854
rect 77782 6618 77866 6854
rect 78102 6618 113546 6854
rect 113782 6618 113866 6854
rect 114102 6618 149546 6854
rect 149782 6618 149866 6854
rect 150102 6618 185546 6854
rect 185782 6618 185866 6854
rect 186102 6618 221546 6854
rect 221782 6618 221866 6854
rect 222102 6618 257546 6854
rect 257782 6618 257866 6854
rect 258102 6618 293546 6854
rect 293782 6618 293866 6854
rect 294102 6618 329546 6854
rect 329782 6618 329866 6854
rect 330102 6618 365546 6854
rect 365782 6618 365866 6854
rect 366102 6618 401546 6854
rect 401782 6618 401866 6854
rect 402102 6618 437546 6854
rect 437782 6618 437866 6854
rect 438102 6618 473546 6854
rect 473782 6618 473866 6854
rect 474102 6618 509546 6854
rect 509782 6618 509866 6854
rect 510102 6618 545546 6854
rect 545782 6618 545866 6854
rect 546102 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 1826 3454
rect 2062 3218 2146 3454
rect 2382 3218 37826 3454
rect 38062 3218 38146 3454
rect 38382 3218 73826 3454
rect 74062 3218 74146 3454
rect 74382 3218 109826 3454
rect 110062 3218 110146 3454
rect 110382 3218 145826 3454
rect 146062 3218 146146 3454
rect 146382 3218 181826 3454
rect 182062 3218 182146 3454
rect 182382 3218 217826 3454
rect 218062 3218 218146 3454
rect 218382 3218 253826 3454
rect 254062 3218 254146 3454
rect 254382 3218 289826 3454
rect 290062 3218 290146 3454
rect 290382 3218 325826 3454
rect 326062 3218 326146 3454
rect 326382 3218 361826 3454
rect 362062 3218 362146 3454
rect 362382 3218 397826 3454
rect 398062 3218 398146 3454
rect 398382 3218 433826 3454
rect 434062 3218 434146 3454
rect 434382 3218 469826 3454
rect 470062 3218 470146 3454
rect 470382 3218 505826 3454
rect 506062 3218 506146 3454
rect 506382 3218 541826 3454
rect 542062 3218 542146 3454
rect 542382 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 1826 3134
rect 2062 2898 2146 3134
rect 2382 2898 37826 3134
rect 38062 2898 38146 3134
rect 38382 2898 73826 3134
rect 74062 2898 74146 3134
rect 74382 2898 109826 3134
rect 110062 2898 110146 3134
rect 110382 2898 145826 3134
rect 146062 2898 146146 3134
rect 146382 2898 181826 3134
rect 182062 2898 182146 3134
rect 182382 2898 217826 3134
rect 218062 2898 218146 3134
rect 218382 2898 253826 3134
rect 254062 2898 254146 3134
rect 254382 2898 289826 3134
rect 290062 2898 290146 3134
rect 290382 2898 325826 3134
rect 326062 2898 326146 3134
rect 326382 2898 361826 3134
rect 362062 2898 362146 3134
rect 362382 2898 397826 3134
rect 398062 2898 398146 3134
rect 398382 2898 433826 3134
rect 434062 2898 434146 3134
rect 434382 2898 469826 3134
rect 470062 2898 470146 3134
rect 470382 2898 505826 3134
rect 506062 2898 506146 3134
rect 506382 2898 541826 3134
rect 542062 2898 542146 3134
rect 542382 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 1826 -346
rect 2062 -582 2146 -346
rect 2382 -582 37826 -346
rect 38062 -582 38146 -346
rect 38382 -582 73826 -346
rect 74062 -582 74146 -346
rect 74382 -582 109826 -346
rect 110062 -582 110146 -346
rect 110382 -582 145826 -346
rect 146062 -582 146146 -346
rect 146382 -582 181826 -346
rect 182062 -582 182146 -346
rect 182382 -582 217826 -346
rect 218062 -582 218146 -346
rect 218382 -582 253826 -346
rect 254062 -582 254146 -346
rect 254382 -582 289826 -346
rect 290062 -582 290146 -346
rect 290382 -582 325826 -346
rect 326062 -582 326146 -346
rect 326382 -582 361826 -346
rect 362062 -582 362146 -346
rect 362382 -582 397826 -346
rect 398062 -582 398146 -346
rect 398382 -582 433826 -346
rect 434062 -582 434146 -346
rect 434382 -582 469826 -346
rect 470062 -582 470146 -346
rect 470382 -582 505826 -346
rect 506062 -582 506146 -346
rect 506382 -582 541826 -346
rect 542062 -582 542146 -346
rect 542382 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 1826 -666
rect 2062 -902 2146 -666
rect 2382 -902 37826 -666
rect 38062 -902 38146 -666
rect 38382 -902 73826 -666
rect 74062 -902 74146 -666
rect 74382 -902 109826 -666
rect 110062 -902 110146 -666
rect 110382 -902 145826 -666
rect 146062 -902 146146 -666
rect 146382 -902 181826 -666
rect 182062 -902 182146 -666
rect 182382 -902 217826 -666
rect 218062 -902 218146 -666
rect 218382 -902 253826 -666
rect 254062 -902 254146 -666
rect 254382 -902 289826 -666
rect 290062 -902 290146 -666
rect 290382 -902 325826 -666
rect 326062 -902 326146 -666
rect 326382 -902 361826 -666
rect 362062 -902 362146 -666
rect 362382 -902 397826 -666
rect 398062 -902 398146 -666
rect 398382 -902 433826 -666
rect 434062 -902 434146 -666
rect 434382 -902 469826 -666
rect 470062 -902 470146 -666
rect 470382 -902 505826 -666
rect 506062 -902 506146 -666
rect 506382 -902 541826 -666
rect 542062 -902 542146 -666
rect 542382 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 19826 -1306
rect 20062 -1542 20146 -1306
rect 20382 -1542 55826 -1306
rect 56062 -1542 56146 -1306
rect 56382 -1542 91826 -1306
rect 92062 -1542 92146 -1306
rect 92382 -1542 127826 -1306
rect 128062 -1542 128146 -1306
rect 128382 -1542 163826 -1306
rect 164062 -1542 164146 -1306
rect 164382 -1542 199826 -1306
rect 200062 -1542 200146 -1306
rect 200382 -1542 235826 -1306
rect 236062 -1542 236146 -1306
rect 236382 -1542 271826 -1306
rect 272062 -1542 272146 -1306
rect 272382 -1542 307826 -1306
rect 308062 -1542 308146 -1306
rect 308382 -1542 343826 -1306
rect 344062 -1542 344146 -1306
rect 344382 -1542 379826 -1306
rect 380062 -1542 380146 -1306
rect 380382 -1542 415826 -1306
rect 416062 -1542 416146 -1306
rect 416382 -1542 451826 -1306
rect 452062 -1542 452146 -1306
rect 452382 -1542 487826 -1306
rect 488062 -1542 488146 -1306
rect 488382 -1542 523826 -1306
rect 524062 -1542 524146 -1306
rect 524382 -1542 559826 -1306
rect 560062 -1542 560146 -1306
rect 560382 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 19826 -1626
rect 20062 -1862 20146 -1626
rect 20382 -1862 55826 -1626
rect 56062 -1862 56146 -1626
rect 56382 -1862 91826 -1626
rect 92062 -1862 92146 -1626
rect 92382 -1862 127826 -1626
rect 128062 -1862 128146 -1626
rect 128382 -1862 163826 -1626
rect 164062 -1862 164146 -1626
rect 164382 -1862 199826 -1626
rect 200062 -1862 200146 -1626
rect 200382 -1862 235826 -1626
rect 236062 -1862 236146 -1626
rect 236382 -1862 271826 -1626
rect 272062 -1862 272146 -1626
rect 272382 -1862 307826 -1626
rect 308062 -1862 308146 -1626
rect 308382 -1862 343826 -1626
rect 344062 -1862 344146 -1626
rect 344382 -1862 379826 -1626
rect 380062 -1862 380146 -1626
rect 380382 -1862 415826 -1626
rect 416062 -1862 416146 -1626
rect 416382 -1862 451826 -1626
rect 452062 -1862 452146 -1626
rect 452382 -1862 487826 -1626
rect 488062 -1862 488146 -1626
rect 488382 -1862 523826 -1626
rect 524062 -1862 524146 -1626
rect 524382 -1862 559826 -1626
rect 560062 -1862 560146 -1626
rect 560382 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use sky130_sram_2kbyte_1rw1r_32x512_8  sram1
timestamp 1640322195
transform 1 0 220000 0 1 400000
box 0 0 136620 83308
use sky130_sram_2kbyte_1rw1r_32x512_8  sram
timestamp 1640322195
transform 1 0 60000 0 1 400000
box 0 0 136620 83308
use user_proj  mprj
timestamp 1640322195
transform 1 0 60000 0 1 60000
box 0 0 164780 166924
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 -1894 74414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 -1894 110414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 -1894 146414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 -1894 182414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 -1894 218414 58000 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 228924 74414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 228924 110414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 228924 146414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 228924 182414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 228924 218414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 -1894 254414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 -1894 290414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 -1894 326414 398000 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 -1894 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 -1894 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 485308 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 485308 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 485308 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 485308 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 485308 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 485308 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 485308 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 485308 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 -1894 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 -1894 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 -1894 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 -1894 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 -1894 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 -1894 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 58000 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 228924 78134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 228924 114134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 228924 150134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 228924 186134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 228924 222134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 398000 6 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 485308 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 485308 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 485308 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 485308 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 485308 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 485308 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 485308 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 485308 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 58000 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 228924 81854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 228924 117854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 228924 153854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 228924 189854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 228924 225854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 398000 6 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 485308 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 485308 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 485308 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 485308 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 485308 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 485308 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 485308 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 485308 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 58000 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 228924 85574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 228924 121574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 228924 157574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 228924 193574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 398000 6 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 485308 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 485308 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 485308 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 485308 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 485308 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 485308 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 485308 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 485308 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 58000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 228924 63854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 228924 99854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 228924 135854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 228924 171854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 398000 6 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 485308 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 485308 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 485308 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 485308 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 228924 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 485308 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 485308 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 485308 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 485308 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 58000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 228924 67574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 228924 103574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 228924 139574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 228924 175574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 398000 6 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 485308 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 485308 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 485308 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 485308 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 228924 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 485308 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 485308 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 485308 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 485308 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 -1894 92414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 -1894 128414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 -1894 164414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 -1894 200414 58000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 228924 92414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 228924 128414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 228924 164414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 -1894 236414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 -1894 272414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 -1894 308414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 -1894 344414 398000 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 -1894 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 -1894 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 485308 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 485308 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 485308 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 228924 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 485308 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 485308 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 485308 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 485308 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 -1894 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 -1894 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 -1894 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 -1894 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 -1894 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 -1894 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 58000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 228924 60134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 228924 96134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 228924 132134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 228924 168134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 398000 6 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 485308 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 485308 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 485308 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 485308 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 228924 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 485308 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 485308 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 485308 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 485308 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
