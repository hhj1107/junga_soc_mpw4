magic
tech sky130A
magscale 1 2
timestamp 1640331715
<< obsli1 >>
rect 1104 1649 164743 165563
<< obsm1 >>
rect 382 8 164758 165572
<< metal2 >>
rect 478 166124 534 166924
rect 1398 166124 1454 166924
rect 2318 166124 2374 166924
rect 3238 166124 3294 166924
rect 4158 166124 4214 166924
rect 5078 166124 5134 166924
rect 5998 166124 6054 166924
rect 6918 166124 6974 166924
rect 7838 166124 7894 166924
rect 8758 166124 8814 166924
rect 9678 166124 9734 166924
rect 10598 166124 10654 166924
rect 11518 166124 11574 166924
rect 12438 166124 12494 166924
rect 13358 166124 13414 166924
rect 14278 166124 14334 166924
rect 15198 166124 15254 166924
rect 16210 166124 16266 166924
rect 17130 166124 17186 166924
rect 18050 166124 18106 166924
rect 18970 166124 19026 166924
rect 19890 166124 19946 166924
rect 20810 166124 20866 166924
rect 21730 166124 21786 166924
rect 22650 166124 22706 166924
rect 23570 166124 23626 166924
rect 24490 166124 24546 166924
rect 25410 166124 25466 166924
rect 26330 166124 26386 166924
rect 27250 166124 27306 166924
rect 28170 166124 28226 166924
rect 29090 166124 29146 166924
rect 30010 166124 30066 166924
rect 31022 166124 31078 166924
rect 31942 166124 31998 166924
rect 32862 166124 32918 166924
rect 33782 166124 33838 166924
rect 34702 166124 34758 166924
rect 35622 166124 35678 166924
rect 36542 166124 36598 166924
rect 37462 166124 37518 166924
rect 38382 166124 38438 166924
rect 39302 166124 39358 166924
rect 40222 166124 40278 166924
rect 41142 166124 41198 166924
rect 42062 166124 42118 166924
rect 42982 166124 43038 166924
rect 43902 166124 43958 166924
rect 44822 166124 44878 166924
rect 45834 166124 45890 166924
rect 46754 166124 46810 166924
rect 47674 166124 47730 166924
rect 48594 166124 48650 166924
rect 49514 166124 49570 166924
rect 50434 166124 50490 166924
rect 51354 166124 51410 166924
rect 52274 166124 52330 166924
rect 53194 166124 53250 166924
rect 54114 166124 54170 166924
rect 55034 166124 55090 166924
rect 55954 166124 56010 166924
rect 56874 166124 56930 166924
rect 57794 166124 57850 166924
rect 58714 166124 58770 166924
rect 59634 166124 59690 166924
rect 60646 166124 60702 166924
rect 61566 166124 61622 166924
rect 62486 166124 62542 166924
rect 63406 166124 63462 166924
rect 64326 166124 64382 166924
rect 65246 166124 65302 166924
rect 66166 166124 66222 166924
rect 67086 166124 67142 166924
rect 68006 166124 68062 166924
rect 68926 166124 68982 166924
rect 69846 166124 69902 166924
rect 70766 166124 70822 166924
rect 71686 166124 71742 166924
rect 72606 166124 72662 166924
rect 73526 166124 73582 166924
rect 74446 166124 74502 166924
rect 75458 166124 75514 166924
rect 76378 166124 76434 166924
rect 77298 166124 77354 166924
rect 78218 166124 78274 166924
rect 79138 166124 79194 166924
rect 80058 166124 80114 166924
rect 80978 166124 81034 166924
rect 81898 166124 81954 166924
rect 82818 166124 82874 166924
rect 83738 166124 83794 166924
rect 84658 166124 84714 166924
rect 85578 166124 85634 166924
rect 86498 166124 86554 166924
rect 87418 166124 87474 166924
rect 88338 166124 88394 166924
rect 89258 166124 89314 166924
rect 90178 166124 90234 166924
rect 91190 166124 91246 166924
rect 92110 166124 92166 166924
rect 93030 166124 93086 166924
rect 93950 166124 94006 166924
rect 94870 166124 94926 166924
rect 95790 166124 95846 166924
rect 96710 166124 96766 166924
rect 97630 166124 97686 166924
rect 98550 166124 98606 166924
rect 99470 166124 99526 166924
rect 100390 166124 100446 166924
rect 101310 166124 101366 166924
rect 102230 166124 102286 166924
rect 103150 166124 103206 166924
rect 104070 166124 104126 166924
rect 104990 166124 105046 166924
rect 106002 166124 106058 166924
rect 106922 166124 106978 166924
rect 107842 166124 107898 166924
rect 108762 166124 108818 166924
rect 109682 166124 109738 166924
rect 110602 166124 110658 166924
rect 111522 166124 111578 166924
rect 112442 166124 112498 166924
rect 113362 166124 113418 166924
rect 114282 166124 114338 166924
rect 115202 166124 115258 166924
rect 116122 166124 116178 166924
rect 117042 166124 117098 166924
rect 117962 166124 118018 166924
rect 118882 166124 118938 166924
rect 119802 166124 119858 166924
rect 120814 166124 120870 166924
rect 121734 166124 121790 166924
rect 122654 166124 122710 166924
rect 123574 166124 123630 166924
rect 124494 166124 124550 166924
rect 125414 166124 125470 166924
rect 126334 166124 126390 166924
rect 127254 166124 127310 166924
rect 128174 166124 128230 166924
rect 129094 166124 129150 166924
rect 130014 166124 130070 166924
rect 130934 166124 130990 166924
rect 131854 166124 131910 166924
rect 132774 166124 132830 166924
rect 133694 166124 133750 166924
rect 134614 166124 134670 166924
rect 135626 166124 135682 166924
rect 136546 166124 136602 166924
rect 137466 166124 137522 166924
rect 138386 166124 138442 166924
rect 139306 166124 139362 166924
rect 140226 166124 140282 166924
rect 141146 166124 141202 166924
rect 142066 166124 142122 166924
rect 142986 166124 143042 166924
rect 143906 166124 143962 166924
rect 144826 166124 144882 166924
rect 145746 166124 145802 166924
rect 146666 166124 146722 166924
rect 147586 166124 147642 166924
rect 148506 166124 148562 166924
rect 149426 166124 149482 166924
rect 150438 166124 150494 166924
rect 151358 166124 151414 166924
rect 152278 166124 152334 166924
rect 153198 166124 153254 166924
rect 154118 166124 154174 166924
rect 155038 166124 155094 166924
rect 155958 166124 156014 166924
rect 156878 166124 156934 166924
rect 157798 166124 157854 166924
rect 158718 166124 158774 166924
rect 159638 166124 159694 166924
rect 160558 166124 160614 166924
rect 161478 166124 161534 166924
rect 162398 166124 162454 166924
rect 163318 166124 163374 166924
rect 164238 166124 164294 166924
rect 110 0 166 800
rect 386 0 442 800
rect 662 0 718 800
rect 938 0 994 800
rect 1306 0 1362 800
rect 1582 0 1638 800
rect 1858 0 1914 800
rect 2134 0 2190 800
rect 2502 0 2558 800
rect 2778 0 2834 800
rect 3054 0 3110 800
rect 3330 0 3386 800
rect 3698 0 3754 800
rect 3974 0 4030 800
rect 4250 0 4306 800
rect 4526 0 4582 800
rect 4894 0 4950 800
rect 5170 0 5226 800
rect 5446 0 5502 800
rect 5722 0 5778 800
rect 6090 0 6146 800
rect 6366 0 6422 800
rect 6642 0 6698 800
rect 6918 0 6974 800
rect 7286 0 7342 800
rect 7562 0 7618 800
rect 7838 0 7894 800
rect 8114 0 8170 800
rect 8482 0 8538 800
rect 8758 0 8814 800
rect 9034 0 9090 800
rect 9310 0 9366 800
rect 9678 0 9734 800
rect 9954 0 10010 800
rect 10230 0 10286 800
rect 10506 0 10562 800
rect 10874 0 10930 800
rect 11150 0 11206 800
rect 11426 0 11482 800
rect 11702 0 11758 800
rect 12070 0 12126 800
rect 12346 0 12402 800
rect 12622 0 12678 800
rect 12990 0 13046 800
rect 13266 0 13322 800
rect 13542 0 13598 800
rect 13818 0 13874 800
rect 14186 0 14242 800
rect 14462 0 14518 800
rect 14738 0 14794 800
rect 15014 0 15070 800
rect 15382 0 15438 800
rect 15658 0 15714 800
rect 15934 0 15990 800
rect 16210 0 16266 800
rect 16578 0 16634 800
rect 16854 0 16910 800
rect 17130 0 17186 800
rect 17406 0 17462 800
rect 17774 0 17830 800
rect 18050 0 18106 800
rect 18326 0 18382 800
rect 18602 0 18658 800
rect 18970 0 19026 800
rect 19246 0 19302 800
rect 19522 0 19578 800
rect 19798 0 19854 800
rect 20166 0 20222 800
rect 20442 0 20498 800
rect 20718 0 20774 800
rect 20994 0 21050 800
rect 21362 0 21418 800
rect 21638 0 21694 800
rect 21914 0 21970 800
rect 22190 0 22246 800
rect 22558 0 22614 800
rect 22834 0 22890 800
rect 23110 0 23166 800
rect 23386 0 23442 800
rect 23754 0 23810 800
rect 24030 0 24086 800
rect 24306 0 24362 800
rect 24674 0 24730 800
rect 24950 0 25006 800
rect 25226 0 25282 800
rect 25502 0 25558 800
rect 25870 0 25926 800
rect 26146 0 26202 800
rect 26422 0 26478 800
rect 26698 0 26754 800
rect 27066 0 27122 800
rect 27342 0 27398 800
rect 27618 0 27674 800
rect 27894 0 27950 800
rect 28262 0 28318 800
rect 28538 0 28594 800
rect 28814 0 28870 800
rect 29090 0 29146 800
rect 29458 0 29514 800
rect 29734 0 29790 800
rect 30010 0 30066 800
rect 30286 0 30342 800
rect 30654 0 30710 800
rect 30930 0 30986 800
rect 31206 0 31262 800
rect 31482 0 31538 800
rect 31850 0 31906 800
rect 32126 0 32182 800
rect 32402 0 32458 800
rect 32678 0 32734 800
rect 33046 0 33102 800
rect 33322 0 33378 800
rect 33598 0 33654 800
rect 33874 0 33930 800
rect 34242 0 34298 800
rect 34518 0 34574 800
rect 34794 0 34850 800
rect 35070 0 35126 800
rect 35438 0 35494 800
rect 35714 0 35770 800
rect 35990 0 36046 800
rect 36358 0 36414 800
rect 36634 0 36690 800
rect 36910 0 36966 800
rect 37186 0 37242 800
rect 37554 0 37610 800
rect 37830 0 37886 800
rect 38106 0 38162 800
rect 38382 0 38438 800
rect 38750 0 38806 800
rect 39026 0 39082 800
rect 39302 0 39358 800
rect 39578 0 39634 800
rect 39946 0 40002 800
rect 40222 0 40278 800
rect 40498 0 40554 800
rect 40774 0 40830 800
rect 41142 0 41198 800
rect 41418 0 41474 800
rect 41694 0 41750 800
rect 41970 0 42026 800
rect 42338 0 42394 800
rect 42614 0 42670 800
rect 42890 0 42946 800
rect 43166 0 43222 800
rect 43534 0 43590 800
rect 43810 0 43866 800
rect 44086 0 44142 800
rect 44362 0 44418 800
rect 44730 0 44786 800
rect 45006 0 45062 800
rect 45282 0 45338 800
rect 45558 0 45614 800
rect 45926 0 45982 800
rect 46202 0 46258 800
rect 46478 0 46534 800
rect 46754 0 46810 800
rect 47122 0 47178 800
rect 47398 0 47454 800
rect 47674 0 47730 800
rect 48042 0 48098 800
rect 48318 0 48374 800
rect 48594 0 48650 800
rect 48870 0 48926 800
rect 49238 0 49294 800
rect 49514 0 49570 800
rect 49790 0 49846 800
rect 50066 0 50122 800
rect 50434 0 50490 800
rect 50710 0 50766 800
rect 50986 0 51042 800
rect 51262 0 51318 800
rect 51630 0 51686 800
rect 51906 0 51962 800
rect 52182 0 52238 800
rect 52458 0 52514 800
rect 52826 0 52882 800
rect 53102 0 53158 800
rect 53378 0 53434 800
rect 53654 0 53710 800
rect 54022 0 54078 800
rect 54298 0 54354 800
rect 54574 0 54630 800
rect 54850 0 54906 800
rect 55218 0 55274 800
rect 55494 0 55550 800
rect 55770 0 55826 800
rect 56046 0 56102 800
rect 56414 0 56470 800
rect 56690 0 56746 800
rect 56966 0 57022 800
rect 57242 0 57298 800
rect 57610 0 57666 800
rect 57886 0 57942 800
rect 58162 0 58218 800
rect 58438 0 58494 800
rect 58806 0 58862 800
rect 59082 0 59138 800
rect 59358 0 59414 800
rect 59726 0 59782 800
rect 60002 0 60058 800
rect 60278 0 60334 800
rect 60554 0 60610 800
rect 60922 0 60978 800
rect 61198 0 61254 800
rect 61474 0 61530 800
rect 61750 0 61806 800
rect 62118 0 62174 800
rect 62394 0 62450 800
rect 62670 0 62726 800
rect 62946 0 63002 800
rect 63314 0 63370 800
rect 63590 0 63646 800
rect 63866 0 63922 800
rect 64142 0 64198 800
rect 64510 0 64566 800
rect 64786 0 64842 800
rect 65062 0 65118 800
rect 65338 0 65394 800
rect 65706 0 65762 800
rect 65982 0 66038 800
rect 66258 0 66314 800
rect 66534 0 66590 800
rect 66902 0 66958 800
rect 67178 0 67234 800
rect 67454 0 67510 800
rect 67730 0 67786 800
rect 68098 0 68154 800
rect 68374 0 68430 800
rect 68650 0 68706 800
rect 68926 0 68982 800
rect 69294 0 69350 800
rect 69570 0 69626 800
rect 69846 0 69902 800
rect 70122 0 70178 800
rect 70490 0 70546 800
rect 70766 0 70822 800
rect 71042 0 71098 800
rect 71410 0 71466 800
rect 71686 0 71742 800
rect 71962 0 72018 800
rect 72238 0 72294 800
rect 72606 0 72662 800
rect 72882 0 72938 800
rect 73158 0 73214 800
rect 73434 0 73490 800
rect 73802 0 73858 800
rect 74078 0 74134 800
rect 74354 0 74410 800
rect 74630 0 74686 800
rect 74998 0 75054 800
rect 75274 0 75330 800
rect 75550 0 75606 800
rect 75826 0 75882 800
rect 76194 0 76250 800
rect 76470 0 76526 800
rect 76746 0 76802 800
rect 77022 0 77078 800
rect 77390 0 77446 800
rect 77666 0 77722 800
rect 77942 0 77998 800
rect 78218 0 78274 800
rect 78586 0 78642 800
rect 78862 0 78918 800
rect 79138 0 79194 800
rect 79414 0 79470 800
rect 79782 0 79838 800
rect 80058 0 80114 800
rect 80334 0 80390 800
rect 80610 0 80666 800
rect 80978 0 81034 800
rect 81254 0 81310 800
rect 81530 0 81586 800
rect 81806 0 81862 800
rect 82174 0 82230 800
rect 82450 0 82506 800
rect 82726 0 82782 800
rect 83094 0 83150 800
rect 83370 0 83426 800
rect 83646 0 83702 800
rect 83922 0 83978 800
rect 84290 0 84346 800
rect 84566 0 84622 800
rect 84842 0 84898 800
rect 85118 0 85174 800
rect 85486 0 85542 800
rect 85762 0 85818 800
rect 86038 0 86094 800
rect 86314 0 86370 800
rect 86682 0 86738 800
rect 86958 0 87014 800
rect 87234 0 87290 800
rect 87510 0 87566 800
rect 87878 0 87934 800
rect 88154 0 88210 800
rect 88430 0 88486 800
rect 88706 0 88762 800
rect 89074 0 89130 800
rect 89350 0 89406 800
rect 89626 0 89682 800
rect 89902 0 89958 800
rect 90270 0 90326 800
rect 90546 0 90602 800
rect 90822 0 90878 800
rect 91098 0 91154 800
rect 91466 0 91522 800
rect 91742 0 91798 800
rect 92018 0 92074 800
rect 92294 0 92350 800
rect 92662 0 92718 800
rect 92938 0 92994 800
rect 93214 0 93270 800
rect 93490 0 93546 800
rect 93858 0 93914 800
rect 94134 0 94190 800
rect 94410 0 94466 800
rect 94778 0 94834 800
rect 95054 0 95110 800
rect 95330 0 95386 800
rect 95606 0 95662 800
rect 95974 0 96030 800
rect 96250 0 96306 800
rect 96526 0 96582 800
rect 96802 0 96858 800
rect 97170 0 97226 800
rect 97446 0 97502 800
rect 97722 0 97778 800
rect 97998 0 98054 800
rect 98366 0 98422 800
rect 98642 0 98698 800
rect 98918 0 98974 800
rect 99194 0 99250 800
rect 99562 0 99618 800
rect 99838 0 99894 800
rect 100114 0 100170 800
rect 100390 0 100446 800
rect 100758 0 100814 800
rect 101034 0 101090 800
rect 101310 0 101366 800
rect 101586 0 101642 800
rect 101954 0 102010 800
rect 102230 0 102286 800
rect 102506 0 102562 800
rect 102782 0 102838 800
rect 103150 0 103206 800
rect 103426 0 103482 800
rect 103702 0 103758 800
rect 103978 0 104034 800
rect 104346 0 104402 800
rect 104622 0 104678 800
rect 104898 0 104954 800
rect 105174 0 105230 800
rect 105542 0 105598 800
rect 105818 0 105874 800
rect 106094 0 106150 800
rect 106462 0 106518 800
rect 106738 0 106794 800
rect 107014 0 107070 800
rect 107290 0 107346 800
rect 107658 0 107714 800
rect 107934 0 107990 800
rect 108210 0 108266 800
rect 108486 0 108542 800
rect 108854 0 108910 800
rect 109130 0 109186 800
rect 109406 0 109462 800
rect 109682 0 109738 800
rect 110050 0 110106 800
rect 110326 0 110382 800
rect 110602 0 110658 800
rect 110878 0 110934 800
rect 111246 0 111302 800
rect 111522 0 111578 800
rect 111798 0 111854 800
rect 112074 0 112130 800
rect 112442 0 112498 800
rect 112718 0 112774 800
rect 112994 0 113050 800
rect 113270 0 113326 800
rect 113638 0 113694 800
rect 113914 0 113970 800
rect 114190 0 114246 800
rect 114466 0 114522 800
rect 114834 0 114890 800
rect 115110 0 115166 800
rect 115386 0 115442 800
rect 115662 0 115718 800
rect 116030 0 116086 800
rect 116306 0 116362 800
rect 116582 0 116638 800
rect 116858 0 116914 800
rect 117226 0 117282 800
rect 117502 0 117558 800
rect 117778 0 117834 800
rect 118146 0 118202 800
rect 118422 0 118478 800
rect 118698 0 118754 800
rect 118974 0 119030 800
rect 119342 0 119398 800
rect 119618 0 119674 800
rect 119894 0 119950 800
rect 120170 0 120226 800
rect 120538 0 120594 800
rect 120814 0 120870 800
rect 121090 0 121146 800
rect 121366 0 121422 800
rect 121734 0 121790 800
rect 122010 0 122066 800
rect 122286 0 122342 800
rect 122562 0 122618 800
rect 122930 0 122986 800
rect 123206 0 123262 800
rect 123482 0 123538 800
rect 123758 0 123814 800
rect 124126 0 124182 800
rect 124402 0 124458 800
rect 124678 0 124734 800
rect 124954 0 125010 800
rect 125322 0 125378 800
rect 125598 0 125654 800
rect 125874 0 125930 800
rect 126150 0 126206 800
rect 126518 0 126574 800
rect 126794 0 126850 800
rect 127070 0 127126 800
rect 127346 0 127402 800
rect 127714 0 127770 800
rect 127990 0 128046 800
rect 128266 0 128322 800
rect 128542 0 128598 800
rect 128910 0 128966 800
rect 129186 0 129242 800
rect 129462 0 129518 800
rect 129830 0 129886 800
rect 130106 0 130162 800
rect 130382 0 130438 800
rect 130658 0 130714 800
rect 131026 0 131082 800
rect 131302 0 131358 800
rect 131578 0 131634 800
rect 131854 0 131910 800
rect 132222 0 132278 800
rect 132498 0 132554 800
rect 132774 0 132830 800
rect 133050 0 133106 800
rect 133418 0 133474 800
rect 133694 0 133750 800
rect 133970 0 134026 800
rect 134246 0 134302 800
rect 134614 0 134670 800
rect 134890 0 134946 800
rect 135166 0 135222 800
rect 135442 0 135498 800
rect 135810 0 135866 800
rect 136086 0 136142 800
rect 136362 0 136418 800
rect 136638 0 136694 800
rect 137006 0 137062 800
rect 137282 0 137338 800
rect 137558 0 137614 800
rect 137834 0 137890 800
rect 138202 0 138258 800
rect 138478 0 138534 800
rect 138754 0 138810 800
rect 139030 0 139086 800
rect 139398 0 139454 800
rect 139674 0 139730 800
rect 139950 0 140006 800
rect 140226 0 140282 800
rect 140594 0 140650 800
rect 140870 0 140926 800
rect 141146 0 141202 800
rect 141514 0 141570 800
rect 141790 0 141846 800
rect 142066 0 142122 800
rect 142342 0 142398 800
rect 142710 0 142766 800
rect 142986 0 143042 800
rect 143262 0 143318 800
rect 143538 0 143594 800
rect 143906 0 143962 800
rect 144182 0 144238 800
rect 144458 0 144514 800
rect 144734 0 144790 800
rect 145102 0 145158 800
rect 145378 0 145434 800
rect 145654 0 145710 800
rect 145930 0 145986 800
rect 146298 0 146354 800
rect 146574 0 146630 800
rect 146850 0 146906 800
rect 147126 0 147182 800
rect 147494 0 147550 800
rect 147770 0 147826 800
rect 148046 0 148102 800
rect 148322 0 148378 800
rect 148690 0 148746 800
rect 148966 0 149022 800
rect 149242 0 149298 800
rect 149518 0 149574 800
rect 149886 0 149942 800
rect 150162 0 150218 800
rect 150438 0 150494 800
rect 150714 0 150770 800
rect 151082 0 151138 800
rect 151358 0 151414 800
rect 151634 0 151690 800
rect 151910 0 151966 800
rect 152278 0 152334 800
rect 152554 0 152610 800
rect 152830 0 152886 800
rect 153198 0 153254 800
rect 153474 0 153530 800
rect 153750 0 153806 800
rect 154026 0 154082 800
rect 154394 0 154450 800
rect 154670 0 154726 800
rect 154946 0 155002 800
rect 155222 0 155278 800
rect 155590 0 155646 800
rect 155866 0 155922 800
rect 156142 0 156198 800
rect 156418 0 156474 800
rect 156786 0 156842 800
rect 157062 0 157118 800
rect 157338 0 157394 800
rect 157614 0 157670 800
rect 157982 0 158038 800
rect 158258 0 158314 800
rect 158534 0 158590 800
rect 158810 0 158866 800
rect 159178 0 159234 800
rect 159454 0 159510 800
rect 159730 0 159786 800
rect 160006 0 160062 800
rect 160374 0 160430 800
rect 160650 0 160706 800
rect 160926 0 160982 800
rect 161202 0 161258 800
rect 161570 0 161626 800
rect 161846 0 161902 800
rect 162122 0 162178 800
rect 162398 0 162454 800
rect 162766 0 162822 800
rect 163042 0 163098 800
rect 163318 0 163374 800
rect 163594 0 163650 800
rect 163962 0 164018 800
rect 164238 0 164294 800
rect 164514 0 164570 800
<< obsm2 >>
rect 110 166068 422 166124
rect 590 166068 1342 166124
rect 1510 166068 2262 166124
rect 2430 166068 3182 166124
rect 3350 166068 4102 166124
rect 4270 166068 5022 166124
rect 5190 166068 5942 166124
rect 6110 166068 6862 166124
rect 7030 166068 7782 166124
rect 7950 166068 8702 166124
rect 8870 166068 9622 166124
rect 9790 166068 10542 166124
rect 10710 166068 11462 166124
rect 11630 166068 12382 166124
rect 12550 166068 13302 166124
rect 13470 166068 14222 166124
rect 14390 166068 15142 166124
rect 15310 166068 16154 166124
rect 16322 166068 17074 166124
rect 17242 166068 17994 166124
rect 18162 166068 18914 166124
rect 19082 166068 19834 166124
rect 20002 166068 20754 166124
rect 20922 166068 21674 166124
rect 21842 166068 22594 166124
rect 22762 166068 23514 166124
rect 23682 166068 24434 166124
rect 24602 166068 25354 166124
rect 25522 166068 26274 166124
rect 26442 166068 27194 166124
rect 27362 166068 28114 166124
rect 28282 166068 29034 166124
rect 29202 166068 29954 166124
rect 30122 166068 30966 166124
rect 31134 166068 31886 166124
rect 32054 166068 32806 166124
rect 32974 166068 33726 166124
rect 33894 166068 34646 166124
rect 34814 166068 35566 166124
rect 35734 166068 36486 166124
rect 36654 166068 37406 166124
rect 37574 166068 38326 166124
rect 38494 166068 39246 166124
rect 39414 166068 40166 166124
rect 40334 166068 41086 166124
rect 41254 166068 42006 166124
rect 42174 166068 42926 166124
rect 43094 166068 43846 166124
rect 44014 166068 44766 166124
rect 44934 166068 45778 166124
rect 45946 166068 46698 166124
rect 46866 166068 47618 166124
rect 47786 166068 48538 166124
rect 48706 166068 49458 166124
rect 49626 166068 50378 166124
rect 50546 166068 51298 166124
rect 51466 166068 52218 166124
rect 52386 166068 53138 166124
rect 53306 166068 54058 166124
rect 54226 166068 54978 166124
rect 55146 166068 55898 166124
rect 56066 166068 56818 166124
rect 56986 166068 57738 166124
rect 57906 166068 58658 166124
rect 58826 166068 59578 166124
rect 59746 166068 60590 166124
rect 60758 166068 61510 166124
rect 61678 166068 62430 166124
rect 62598 166068 63350 166124
rect 63518 166068 64270 166124
rect 64438 166068 65190 166124
rect 65358 166068 66110 166124
rect 66278 166068 67030 166124
rect 67198 166068 67950 166124
rect 68118 166068 68870 166124
rect 69038 166068 69790 166124
rect 69958 166068 70710 166124
rect 70878 166068 71630 166124
rect 71798 166068 72550 166124
rect 72718 166068 73470 166124
rect 73638 166068 74390 166124
rect 74558 166068 75402 166124
rect 75570 166068 76322 166124
rect 76490 166068 77242 166124
rect 77410 166068 78162 166124
rect 78330 166068 79082 166124
rect 79250 166068 80002 166124
rect 80170 166068 80922 166124
rect 81090 166068 81842 166124
rect 82010 166068 82762 166124
rect 82930 166068 83682 166124
rect 83850 166068 84602 166124
rect 84770 166068 85522 166124
rect 85690 166068 86442 166124
rect 86610 166068 87362 166124
rect 87530 166068 88282 166124
rect 88450 166068 89202 166124
rect 89370 166068 90122 166124
rect 90290 166068 91134 166124
rect 91302 166068 92054 166124
rect 92222 166068 92974 166124
rect 93142 166068 93894 166124
rect 94062 166068 94814 166124
rect 94982 166068 95734 166124
rect 95902 166068 96654 166124
rect 96822 166068 97574 166124
rect 97742 166068 98494 166124
rect 98662 166068 99414 166124
rect 99582 166068 100334 166124
rect 100502 166068 101254 166124
rect 101422 166068 102174 166124
rect 102342 166068 103094 166124
rect 103262 166068 104014 166124
rect 104182 166068 104934 166124
rect 105102 166068 105946 166124
rect 106114 166068 106866 166124
rect 107034 166068 107786 166124
rect 107954 166068 108706 166124
rect 108874 166068 109626 166124
rect 109794 166068 110546 166124
rect 110714 166068 111466 166124
rect 111634 166068 112386 166124
rect 112554 166068 113306 166124
rect 113474 166068 114226 166124
rect 114394 166068 115146 166124
rect 115314 166068 116066 166124
rect 116234 166068 116986 166124
rect 117154 166068 117906 166124
rect 118074 166068 118826 166124
rect 118994 166068 119746 166124
rect 119914 166068 120758 166124
rect 120926 166068 121678 166124
rect 121846 166068 122598 166124
rect 122766 166068 123518 166124
rect 123686 166068 124438 166124
rect 124606 166068 125358 166124
rect 125526 166068 126278 166124
rect 126446 166068 127198 166124
rect 127366 166068 128118 166124
rect 128286 166068 129038 166124
rect 129206 166068 129958 166124
rect 130126 166068 130878 166124
rect 131046 166068 131798 166124
rect 131966 166068 132718 166124
rect 132886 166068 133638 166124
rect 133806 166068 134558 166124
rect 134726 166068 135570 166124
rect 135738 166068 136490 166124
rect 136658 166068 137410 166124
rect 137578 166068 138330 166124
rect 138498 166068 139250 166124
rect 139418 166068 140170 166124
rect 140338 166068 141090 166124
rect 141258 166068 142010 166124
rect 142178 166068 142930 166124
rect 143098 166068 143850 166124
rect 144018 166068 144770 166124
rect 144938 166068 145690 166124
rect 145858 166068 146610 166124
rect 146778 166068 147530 166124
rect 147698 166068 148450 166124
rect 148618 166068 149370 166124
rect 149538 166068 150382 166124
rect 150550 166068 151302 166124
rect 151470 166068 152222 166124
rect 152390 166068 153142 166124
rect 153310 166068 154062 166124
rect 154230 166068 154982 166124
rect 155150 166068 155902 166124
rect 156070 166068 156822 166124
rect 156990 166068 157742 166124
rect 157910 166068 158662 166124
rect 158830 166068 159582 166124
rect 159750 166068 160502 166124
rect 160670 166068 161422 166124
rect 161590 166068 162342 166124
rect 162510 166068 163262 166124
rect 163430 166068 164182 166124
rect 164350 166068 164754 166124
rect 110 856 164754 166068
rect 222 2 330 856
rect 498 2 606 856
rect 774 2 882 856
rect 1050 2 1250 856
rect 1418 2 1526 856
rect 1694 2 1802 856
rect 1970 2 2078 856
rect 2246 2 2446 856
rect 2614 2 2722 856
rect 2890 2 2998 856
rect 3166 2 3274 856
rect 3442 2 3642 856
rect 3810 2 3918 856
rect 4086 2 4194 856
rect 4362 2 4470 856
rect 4638 2 4838 856
rect 5006 2 5114 856
rect 5282 2 5390 856
rect 5558 2 5666 856
rect 5834 2 6034 856
rect 6202 2 6310 856
rect 6478 2 6586 856
rect 6754 2 6862 856
rect 7030 2 7230 856
rect 7398 2 7506 856
rect 7674 2 7782 856
rect 7950 2 8058 856
rect 8226 2 8426 856
rect 8594 2 8702 856
rect 8870 2 8978 856
rect 9146 2 9254 856
rect 9422 2 9622 856
rect 9790 2 9898 856
rect 10066 2 10174 856
rect 10342 2 10450 856
rect 10618 2 10818 856
rect 10986 2 11094 856
rect 11262 2 11370 856
rect 11538 2 11646 856
rect 11814 2 12014 856
rect 12182 2 12290 856
rect 12458 2 12566 856
rect 12734 2 12934 856
rect 13102 2 13210 856
rect 13378 2 13486 856
rect 13654 2 13762 856
rect 13930 2 14130 856
rect 14298 2 14406 856
rect 14574 2 14682 856
rect 14850 2 14958 856
rect 15126 2 15326 856
rect 15494 2 15602 856
rect 15770 2 15878 856
rect 16046 2 16154 856
rect 16322 2 16522 856
rect 16690 2 16798 856
rect 16966 2 17074 856
rect 17242 2 17350 856
rect 17518 2 17718 856
rect 17886 2 17994 856
rect 18162 2 18270 856
rect 18438 2 18546 856
rect 18714 2 18914 856
rect 19082 2 19190 856
rect 19358 2 19466 856
rect 19634 2 19742 856
rect 19910 2 20110 856
rect 20278 2 20386 856
rect 20554 2 20662 856
rect 20830 2 20938 856
rect 21106 2 21306 856
rect 21474 2 21582 856
rect 21750 2 21858 856
rect 22026 2 22134 856
rect 22302 2 22502 856
rect 22670 2 22778 856
rect 22946 2 23054 856
rect 23222 2 23330 856
rect 23498 2 23698 856
rect 23866 2 23974 856
rect 24142 2 24250 856
rect 24418 2 24618 856
rect 24786 2 24894 856
rect 25062 2 25170 856
rect 25338 2 25446 856
rect 25614 2 25814 856
rect 25982 2 26090 856
rect 26258 2 26366 856
rect 26534 2 26642 856
rect 26810 2 27010 856
rect 27178 2 27286 856
rect 27454 2 27562 856
rect 27730 2 27838 856
rect 28006 2 28206 856
rect 28374 2 28482 856
rect 28650 2 28758 856
rect 28926 2 29034 856
rect 29202 2 29402 856
rect 29570 2 29678 856
rect 29846 2 29954 856
rect 30122 2 30230 856
rect 30398 2 30598 856
rect 30766 2 30874 856
rect 31042 2 31150 856
rect 31318 2 31426 856
rect 31594 2 31794 856
rect 31962 2 32070 856
rect 32238 2 32346 856
rect 32514 2 32622 856
rect 32790 2 32990 856
rect 33158 2 33266 856
rect 33434 2 33542 856
rect 33710 2 33818 856
rect 33986 2 34186 856
rect 34354 2 34462 856
rect 34630 2 34738 856
rect 34906 2 35014 856
rect 35182 2 35382 856
rect 35550 2 35658 856
rect 35826 2 35934 856
rect 36102 2 36302 856
rect 36470 2 36578 856
rect 36746 2 36854 856
rect 37022 2 37130 856
rect 37298 2 37498 856
rect 37666 2 37774 856
rect 37942 2 38050 856
rect 38218 2 38326 856
rect 38494 2 38694 856
rect 38862 2 38970 856
rect 39138 2 39246 856
rect 39414 2 39522 856
rect 39690 2 39890 856
rect 40058 2 40166 856
rect 40334 2 40442 856
rect 40610 2 40718 856
rect 40886 2 41086 856
rect 41254 2 41362 856
rect 41530 2 41638 856
rect 41806 2 41914 856
rect 42082 2 42282 856
rect 42450 2 42558 856
rect 42726 2 42834 856
rect 43002 2 43110 856
rect 43278 2 43478 856
rect 43646 2 43754 856
rect 43922 2 44030 856
rect 44198 2 44306 856
rect 44474 2 44674 856
rect 44842 2 44950 856
rect 45118 2 45226 856
rect 45394 2 45502 856
rect 45670 2 45870 856
rect 46038 2 46146 856
rect 46314 2 46422 856
rect 46590 2 46698 856
rect 46866 2 47066 856
rect 47234 2 47342 856
rect 47510 2 47618 856
rect 47786 2 47986 856
rect 48154 2 48262 856
rect 48430 2 48538 856
rect 48706 2 48814 856
rect 48982 2 49182 856
rect 49350 2 49458 856
rect 49626 2 49734 856
rect 49902 2 50010 856
rect 50178 2 50378 856
rect 50546 2 50654 856
rect 50822 2 50930 856
rect 51098 2 51206 856
rect 51374 2 51574 856
rect 51742 2 51850 856
rect 52018 2 52126 856
rect 52294 2 52402 856
rect 52570 2 52770 856
rect 52938 2 53046 856
rect 53214 2 53322 856
rect 53490 2 53598 856
rect 53766 2 53966 856
rect 54134 2 54242 856
rect 54410 2 54518 856
rect 54686 2 54794 856
rect 54962 2 55162 856
rect 55330 2 55438 856
rect 55606 2 55714 856
rect 55882 2 55990 856
rect 56158 2 56358 856
rect 56526 2 56634 856
rect 56802 2 56910 856
rect 57078 2 57186 856
rect 57354 2 57554 856
rect 57722 2 57830 856
rect 57998 2 58106 856
rect 58274 2 58382 856
rect 58550 2 58750 856
rect 58918 2 59026 856
rect 59194 2 59302 856
rect 59470 2 59670 856
rect 59838 2 59946 856
rect 60114 2 60222 856
rect 60390 2 60498 856
rect 60666 2 60866 856
rect 61034 2 61142 856
rect 61310 2 61418 856
rect 61586 2 61694 856
rect 61862 2 62062 856
rect 62230 2 62338 856
rect 62506 2 62614 856
rect 62782 2 62890 856
rect 63058 2 63258 856
rect 63426 2 63534 856
rect 63702 2 63810 856
rect 63978 2 64086 856
rect 64254 2 64454 856
rect 64622 2 64730 856
rect 64898 2 65006 856
rect 65174 2 65282 856
rect 65450 2 65650 856
rect 65818 2 65926 856
rect 66094 2 66202 856
rect 66370 2 66478 856
rect 66646 2 66846 856
rect 67014 2 67122 856
rect 67290 2 67398 856
rect 67566 2 67674 856
rect 67842 2 68042 856
rect 68210 2 68318 856
rect 68486 2 68594 856
rect 68762 2 68870 856
rect 69038 2 69238 856
rect 69406 2 69514 856
rect 69682 2 69790 856
rect 69958 2 70066 856
rect 70234 2 70434 856
rect 70602 2 70710 856
rect 70878 2 70986 856
rect 71154 2 71354 856
rect 71522 2 71630 856
rect 71798 2 71906 856
rect 72074 2 72182 856
rect 72350 2 72550 856
rect 72718 2 72826 856
rect 72994 2 73102 856
rect 73270 2 73378 856
rect 73546 2 73746 856
rect 73914 2 74022 856
rect 74190 2 74298 856
rect 74466 2 74574 856
rect 74742 2 74942 856
rect 75110 2 75218 856
rect 75386 2 75494 856
rect 75662 2 75770 856
rect 75938 2 76138 856
rect 76306 2 76414 856
rect 76582 2 76690 856
rect 76858 2 76966 856
rect 77134 2 77334 856
rect 77502 2 77610 856
rect 77778 2 77886 856
rect 78054 2 78162 856
rect 78330 2 78530 856
rect 78698 2 78806 856
rect 78974 2 79082 856
rect 79250 2 79358 856
rect 79526 2 79726 856
rect 79894 2 80002 856
rect 80170 2 80278 856
rect 80446 2 80554 856
rect 80722 2 80922 856
rect 81090 2 81198 856
rect 81366 2 81474 856
rect 81642 2 81750 856
rect 81918 2 82118 856
rect 82286 2 82394 856
rect 82562 2 82670 856
rect 82838 2 83038 856
rect 83206 2 83314 856
rect 83482 2 83590 856
rect 83758 2 83866 856
rect 84034 2 84234 856
rect 84402 2 84510 856
rect 84678 2 84786 856
rect 84954 2 85062 856
rect 85230 2 85430 856
rect 85598 2 85706 856
rect 85874 2 85982 856
rect 86150 2 86258 856
rect 86426 2 86626 856
rect 86794 2 86902 856
rect 87070 2 87178 856
rect 87346 2 87454 856
rect 87622 2 87822 856
rect 87990 2 88098 856
rect 88266 2 88374 856
rect 88542 2 88650 856
rect 88818 2 89018 856
rect 89186 2 89294 856
rect 89462 2 89570 856
rect 89738 2 89846 856
rect 90014 2 90214 856
rect 90382 2 90490 856
rect 90658 2 90766 856
rect 90934 2 91042 856
rect 91210 2 91410 856
rect 91578 2 91686 856
rect 91854 2 91962 856
rect 92130 2 92238 856
rect 92406 2 92606 856
rect 92774 2 92882 856
rect 93050 2 93158 856
rect 93326 2 93434 856
rect 93602 2 93802 856
rect 93970 2 94078 856
rect 94246 2 94354 856
rect 94522 2 94722 856
rect 94890 2 94998 856
rect 95166 2 95274 856
rect 95442 2 95550 856
rect 95718 2 95918 856
rect 96086 2 96194 856
rect 96362 2 96470 856
rect 96638 2 96746 856
rect 96914 2 97114 856
rect 97282 2 97390 856
rect 97558 2 97666 856
rect 97834 2 97942 856
rect 98110 2 98310 856
rect 98478 2 98586 856
rect 98754 2 98862 856
rect 99030 2 99138 856
rect 99306 2 99506 856
rect 99674 2 99782 856
rect 99950 2 100058 856
rect 100226 2 100334 856
rect 100502 2 100702 856
rect 100870 2 100978 856
rect 101146 2 101254 856
rect 101422 2 101530 856
rect 101698 2 101898 856
rect 102066 2 102174 856
rect 102342 2 102450 856
rect 102618 2 102726 856
rect 102894 2 103094 856
rect 103262 2 103370 856
rect 103538 2 103646 856
rect 103814 2 103922 856
rect 104090 2 104290 856
rect 104458 2 104566 856
rect 104734 2 104842 856
rect 105010 2 105118 856
rect 105286 2 105486 856
rect 105654 2 105762 856
rect 105930 2 106038 856
rect 106206 2 106406 856
rect 106574 2 106682 856
rect 106850 2 106958 856
rect 107126 2 107234 856
rect 107402 2 107602 856
rect 107770 2 107878 856
rect 108046 2 108154 856
rect 108322 2 108430 856
rect 108598 2 108798 856
rect 108966 2 109074 856
rect 109242 2 109350 856
rect 109518 2 109626 856
rect 109794 2 109994 856
rect 110162 2 110270 856
rect 110438 2 110546 856
rect 110714 2 110822 856
rect 110990 2 111190 856
rect 111358 2 111466 856
rect 111634 2 111742 856
rect 111910 2 112018 856
rect 112186 2 112386 856
rect 112554 2 112662 856
rect 112830 2 112938 856
rect 113106 2 113214 856
rect 113382 2 113582 856
rect 113750 2 113858 856
rect 114026 2 114134 856
rect 114302 2 114410 856
rect 114578 2 114778 856
rect 114946 2 115054 856
rect 115222 2 115330 856
rect 115498 2 115606 856
rect 115774 2 115974 856
rect 116142 2 116250 856
rect 116418 2 116526 856
rect 116694 2 116802 856
rect 116970 2 117170 856
rect 117338 2 117446 856
rect 117614 2 117722 856
rect 117890 2 118090 856
rect 118258 2 118366 856
rect 118534 2 118642 856
rect 118810 2 118918 856
rect 119086 2 119286 856
rect 119454 2 119562 856
rect 119730 2 119838 856
rect 120006 2 120114 856
rect 120282 2 120482 856
rect 120650 2 120758 856
rect 120926 2 121034 856
rect 121202 2 121310 856
rect 121478 2 121678 856
rect 121846 2 121954 856
rect 122122 2 122230 856
rect 122398 2 122506 856
rect 122674 2 122874 856
rect 123042 2 123150 856
rect 123318 2 123426 856
rect 123594 2 123702 856
rect 123870 2 124070 856
rect 124238 2 124346 856
rect 124514 2 124622 856
rect 124790 2 124898 856
rect 125066 2 125266 856
rect 125434 2 125542 856
rect 125710 2 125818 856
rect 125986 2 126094 856
rect 126262 2 126462 856
rect 126630 2 126738 856
rect 126906 2 127014 856
rect 127182 2 127290 856
rect 127458 2 127658 856
rect 127826 2 127934 856
rect 128102 2 128210 856
rect 128378 2 128486 856
rect 128654 2 128854 856
rect 129022 2 129130 856
rect 129298 2 129406 856
rect 129574 2 129774 856
rect 129942 2 130050 856
rect 130218 2 130326 856
rect 130494 2 130602 856
rect 130770 2 130970 856
rect 131138 2 131246 856
rect 131414 2 131522 856
rect 131690 2 131798 856
rect 131966 2 132166 856
rect 132334 2 132442 856
rect 132610 2 132718 856
rect 132886 2 132994 856
rect 133162 2 133362 856
rect 133530 2 133638 856
rect 133806 2 133914 856
rect 134082 2 134190 856
rect 134358 2 134558 856
rect 134726 2 134834 856
rect 135002 2 135110 856
rect 135278 2 135386 856
rect 135554 2 135754 856
rect 135922 2 136030 856
rect 136198 2 136306 856
rect 136474 2 136582 856
rect 136750 2 136950 856
rect 137118 2 137226 856
rect 137394 2 137502 856
rect 137670 2 137778 856
rect 137946 2 138146 856
rect 138314 2 138422 856
rect 138590 2 138698 856
rect 138866 2 138974 856
rect 139142 2 139342 856
rect 139510 2 139618 856
rect 139786 2 139894 856
rect 140062 2 140170 856
rect 140338 2 140538 856
rect 140706 2 140814 856
rect 140982 2 141090 856
rect 141258 2 141458 856
rect 141626 2 141734 856
rect 141902 2 142010 856
rect 142178 2 142286 856
rect 142454 2 142654 856
rect 142822 2 142930 856
rect 143098 2 143206 856
rect 143374 2 143482 856
rect 143650 2 143850 856
rect 144018 2 144126 856
rect 144294 2 144402 856
rect 144570 2 144678 856
rect 144846 2 145046 856
rect 145214 2 145322 856
rect 145490 2 145598 856
rect 145766 2 145874 856
rect 146042 2 146242 856
rect 146410 2 146518 856
rect 146686 2 146794 856
rect 146962 2 147070 856
rect 147238 2 147438 856
rect 147606 2 147714 856
rect 147882 2 147990 856
rect 148158 2 148266 856
rect 148434 2 148634 856
rect 148802 2 148910 856
rect 149078 2 149186 856
rect 149354 2 149462 856
rect 149630 2 149830 856
rect 149998 2 150106 856
rect 150274 2 150382 856
rect 150550 2 150658 856
rect 150826 2 151026 856
rect 151194 2 151302 856
rect 151470 2 151578 856
rect 151746 2 151854 856
rect 152022 2 152222 856
rect 152390 2 152498 856
rect 152666 2 152774 856
rect 152942 2 153142 856
rect 153310 2 153418 856
rect 153586 2 153694 856
rect 153862 2 153970 856
rect 154138 2 154338 856
rect 154506 2 154614 856
rect 154782 2 154890 856
rect 155058 2 155166 856
rect 155334 2 155534 856
rect 155702 2 155810 856
rect 155978 2 156086 856
rect 156254 2 156362 856
rect 156530 2 156730 856
rect 156898 2 157006 856
rect 157174 2 157282 856
rect 157450 2 157558 856
rect 157726 2 157926 856
rect 158094 2 158202 856
rect 158370 2 158478 856
rect 158646 2 158754 856
rect 158922 2 159122 856
rect 159290 2 159398 856
rect 159566 2 159674 856
rect 159842 2 159950 856
rect 160118 2 160318 856
rect 160486 2 160594 856
rect 160762 2 160870 856
rect 161038 2 161146 856
rect 161314 2 161514 856
rect 161682 2 161790 856
rect 161958 2 162066 856
rect 162234 2 162342 856
rect 162510 2 162710 856
rect 162878 2 162986 856
rect 163154 2 163262 856
rect 163430 2 163538 856
rect 163706 2 163906 856
rect 164074 2 164182 856
rect 164350 2 164458 856
rect 164626 2 164754 856
<< metal3 >>
rect 163980 165520 164780 165640
rect 0 165112 800 165232
rect 163980 163072 164780 163192
rect 0 161984 800 162104
rect 163980 160624 164780 160744
rect 0 158856 800 158976
rect 163980 158176 164780 158296
rect 0 155728 800 155848
rect 163980 155728 164780 155848
rect 163980 153280 164780 153400
rect 0 152600 800 152720
rect 163980 150832 164780 150952
rect 0 149472 800 149592
rect 163980 148384 164780 148504
rect 0 146208 800 146328
rect 163980 145936 164780 146056
rect 163980 143488 164780 143608
rect 0 143080 800 143200
rect 163980 141040 164780 141160
rect 0 139952 800 140072
rect 163980 138592 164780 138712
rect 0 136824 800 136944
rect 163980 136144 164780 136264
rect 0 133696 800 133816
rect 163980 133696 164780 133816
rect 163980 131248 164780 131368
rect 0 130568 800 130688
rect 163980 128800 164780 128920
rect 0 127440 800 127560
rect 163980 126352 164780 126472
rect 0 124176 800 124296
rect 163980 123904 164780 124024
rect 163980 121456 164780 121576
rect 0 121048 800 121168
rect 163980 119008 164780 119128
rect 0 117920 800 118040
rect 163980 116560 164780 116680
rect 0 114792 800 114912
rect 163980 114112 164780 114232
rect 0 111664 800 111784
rect 163980 111528 164780 111648
rect 163980 109080 164780 109200
rect 0 108536 800 108656
rect 163980 106632 164780 106752
rect 0 105272 800 105392
rect 163980 104184 164780 104304
rect 0 102144 800 102264
rect 163980 101736 164780 101856
rect 163980 99288 164780 99408
rect 0 99016 800 99136
rect 163980 96840 164780 96960
rect 0 95888 800 96008
rect 163980 94392 164780 94512
rect 0 92760 800 92880
rect 163980 91944 164780 92064
rect 0 89632 800 89752
rect 163980 89496 164780 89616
rect 163980 87048 164780 87168
rect 0 86504 800 86624
rect 163980 84600 164780 84720
rect 0 83240 800 83360
rect 163980 82152 164780 82272
rect 0 80112 800 80232
rect 163980 79704 164780 79824
rect 163980 77256 164780 77376
rect 0 76984 800 77104
rect 163980 74808 164780 74928
rect 0 73856 800 73976
rect 163980 72360 164780 72480
rect 0 70728 800 70848
rect 163980 69912 164780 70032
rect 0 67600 800 67720
rect 163980 67464 164780 67584
rect 163980 65016 164780 65136
rect 0 64472 800 64592
rect 163980 62568 164780 62688
rect 0 61208 800 61328
rect 163980 60120 164780 60240
rect 0 58080 800 58200
rect 163980 57672 164780 57792
rect 0 54952 800 55072
rect 163980 55088 164780 55208
rect 163980 52640 164780 52760
rect 0 51824 800 51944
rect 163980 50192 164780 50312
rect 0 48696 800 48816
rect 163980 47744 164780 47864
rect 0 45568 800 45688
rect 163980 45296 164780 45416
rect 163980 42848 164780 42968
rect 0 42304 800 42424
rect 163980 40400 164780 40520
rect 0 39176 800 39296
rect 163980 37952 164780 38072
rect 0 36048 800 36168
rect 163980 35504 164780 35624
rect 0 32920 800 33040
rect 163980 33056 164780 33176
rect 163980 30608 164780 30728
rect 0 29792 800 29912
rect 163980 28160 164780 28280
rect 0 26664 800 26784
rect 163980 25712 164780 25832
rect 0 23536 800 23656
rect 163980 23264 164780 23384
rect 163980 20816 164780 20936
rect 0 20272 800 20392
rect 163980 18368 164780 18488
rect 0 17144 800 17264
rect 163980 15920 164780 16040
rect 0 14016 800 14136
rect 163980 13472 164780 13592
rect 0 10888 800 11008
rect 163980 11024 164780 11144
rect 163980 8576 164780 8696
rect 0 7760 800 7880
rect 163980 6128 164780 6248
rect 0 4632 800 4752
rect 163980 3680 164780 3800
rect 0 1504 800 1624
rect 163980 1232 164780 1352
<< obsm3 >>
rect 105 165440 163900 165613
rect 105 165312 164759 165440
rect 880 165032 164759 165312
rect 105 163272 164759 165032
rect 105 162992 163900 163272
rect 105 162184 164759 162992
rect 880 161904 164759 162184
rect 105 160824 164759 161904
rect 105 160544 163900 160824
rect 105 159056 164759 160544
rect 880 158776 164759 159056
rect 105 158376 164759 158776
rect 105 158096 163900 158376
rect 105 155928 164759 158096
rect 880 155648 163900 155928
rect 105 153480 164759 155648
rect 105 153200 163900 153480
rect 105 152800 164759 153200
rect 880 152520 164759 152800
rect 105 151032 164759 152520
rect 105 150752 163900 151032
rect 105 149672 164759 150752
rect 880 149392 164759 149672
rect 105 148584 164759 149392
rect 105 148304 163900 148584
rect 105 146408 164759 148304
rect 880 146136 164759 146408
rect 880 146128 163900 146136
rect 105 145856 163900 146128
rect 105 143688 164759 145856
rect 105 143408 163900 143688
rect 105 143280 164759 143408
rect 880 143000 164759 143280
rect 105 141240 164759 143000
rect 105 140960 163900 141240
rect 105 140152 164759 140960
rect 880 139872 164759 140152
rect 105 138792 164759 139872
rect 105 138512 163900 138792
rect 105 137024 164759 138512
rect 880 136744 164759 137024
rect 105 136344 164759 136744
rect 105 136064 163900 136344
rect 105 133896 164759 136064
rect 880 133616 163900 133896
rect 105 131448 164759 133616
rect 105 131168 163900 131448
rect 105 130768 164759 131168
rect 880 130488 164759 130768
rect 105 129000 164759 130488
rect 105 128720 163900 129000
rect 105 127640 164759 128720
rect 880 127360 164759 127640
rect 105 126552 164759 127360
rect 105 126272 163900 126552
rect 105 124376 164759 126272
rect 880 124104 164759 124376
rect 880 124096 163900 124104
rect 105 123824 163900 124096
rect 105 121656 164759 123824
rect 105 121376 163900 121656
rect 105 121248 164759 121376
rect 880 120968 164759 121248
rect 105 119208 164759 120968
rect 105 118928 163900 119208
rect 105 118120 164759 118928
rect 880 117840 164759 118120
rect 105 116760 164759 117840
rect 105 116480 163900 116760
rect 105 114992 164759 116480
rect 880 114712 164759 114992
rect 105 114312 164759 114712
rect 105 114032 163900 114312
rect 105 111864 164759 114032
rect 880 111728 164759 111864
rect 880 111584 163900 111728
rect 105 111448 163900 111584
rect 105 109280 164759 111448
rect 105 109000 163900 109280
rect 105 108736 164759 109000
rect 880 108456 164759 108736
rect 105 106832 164759 108456
rect 105 106552 163900 106832
rect 105 105472 164759 106552
rect 880 105192 164759 105472
rect 105 104384 164759 105192
rect 105 104104 163900 104384
rect 105 102344 164759 104104
rect 880 102064 164759 102344
rect 105 101936 164759 102064
rect 105 101656 163900 101936
rect 105 99488 164759 101656
rect 105 99216 163900 99488
rect 880 99208 163900 99216
rect 880 98936 164759 99208
rect 105 97040 164759 98936
rect 105 96760 163900 97040
rect 105 96088 164759 96760
rect 880 95808 164759 96088
rect 105 94592 164759 95808
rect 105 94312 163900 94592
rect 105 92960 164759 94312
rect 880 92680 164759 92960
rect 105 92144 164759 92680
rect 105 91864 163900 92144
rect 105 89832 164759 91864
rect 880 89696 164759 89832
rect 880 89552 163900 89696
rect 105 89416 163900 89552
rect 105 87248 164759 89416
rect 105 86968 163900 87248
rect 105 86704 164759 86968
rect 880 86424 164759 86704
rect 105 84800 164759 86424
rect 105 84520 163900 84800
rect 105 83440 164759 84520
rect 880 83160 164759 83440
rect 105 82352 164759 83160
rect 105 82072 163900 82352
rect 105 80312 164759 82072
rect 880 80032 164759 80312
rect 105 79904 164759 80032
rect 105 79624 163900 79904
rect 105 77456 164759 79624
rect 105 77184 163900 77456
rect 880 77176 163900 77184
rect 880 76904 164759 77176
rect 105 75008 164759 76904
rect 105 74728 163900 75008
rect 105 74056 164759 74728
rect 880 73776 164759 74056
rect 105 72560 164759 73776
rect 105 72280 163900 72560
rect 105 70928 164759 72280
rect 880 70648 164759 70928
rect 105 70112 164759 70648
rect 105 69832 163900 70112
rect 105 67800 164759 69832
rect 880 67664 164759 67800
rect 880 67520 163900 67664
rect 105 67384 163900 67520
rect 105 65216 164759 67384
rect 105 64936 163900 65216
rect 105 64672 164759 64936
rect 880 64392 164759 64672
rect 105 62768 164759 64392
rect 105 62488 163900 62768
rect 105 61408 164759 62488
rect 880 61128 164759 61408
rect 105 60320 164759 61128
rect 105 60040 163900 60320
rect 105 58280 164759 60040
rect 880 58000 164759 58280
rect 105 57872 164759 58000
rect 105 57592 163900 57872
rect 105 55288 164759 57592
rect 105 55152 163900 55288
rect 880 55008 163900 55152
rect 880 54872 164759 55008
rect 105 52840 164759 54872
rect 105 52560 163900 52840
rect 105 52024 164759 52560
rect 880 51744 164759 52024
rect 105 50392 164759 51744
rect 105 50112 163900 50392
rect 105 48896 164759 50112
rect 880 48616 164759 48896
rect 105 47944 164759 48616
rect 105 47664 163900 47944
rect 105 45768 164759 47664
rect 880 45496 164759 45768
rect 880 45488 163900 45496
rect 105 45216 163900 45488
rect 105 43048 164759 45216
rect 105 42768 163900 43048
rect 105 42504 164759 42768
rect 880 42224 164759 42504
rect 105 40600 164759 42224
rect 105 40320 163900 40600
rect 105 39376 164759 40320
rect 880 39096 164759 39376
rect 105 38152 164759 39096
rect 105 37872 163900 38152
rect 105 36248 164759 37872
rect 880 35968 164759 36248
rect 105 35704 164759 35968
rect 105 35424 163900 35704
rect 105 33256 164759 35424
rect 105 33120 163900 33256
rect 880 32976 163900 33120
rect 880 32840 164759 32976
rect 105 30808 164759 32840
rect 105 30528 163900 30808
rect 105 29992 164759 30528
rect 880 29712 164759 29992
rect 105 28360 164759 29712
rect 105 28080 163900 28360
rect 105 26864 164759 28080
rect 880 26584 164759 26864
rect 105 25912 164759 26584
rect 105 25632 163900 25912
rect 105 23736 164759 25632
rect 880 23464 164759 23736
rect 880 23456 163900 23464
rect 105 23184 163900 23456
rect 105 21016 164759 23184
rect 105 20736 163900 21016
rect 105 20472 164759 20736
rect 880 20192 164759 20472
rect 105 18568 164759 20192
rect 105 18288 163900 18568
rect 105 17344 164759 18288
rect 880 17064 164759 17344
rect 105 16120 164759 17064
rect 105 15840 163900 16120
rect 105 14216 164759 15840
rect 880 13936 164759 14216
rect 105 13672 164759 13936
rect 105 13392 163900 13672
rect 105 11224 164759 13392
rect 105 11088 163900 11224
rect 880 10944 163900 11088
rect 880 10808 164759 10944
rect 105 8776 164759 10808
rect 105 8496 163900 8776
rect 105 7960 164759 8496
rect 880 7680 164759 7960
rect 105 6328 164759 7680
rect 105 6048 163900 6328
rect 105 4832 164759 6048
rect 880 4552 164759 4832
rect 105 3880 164759 4552
rect 105 3600 163900 3880
rect 105 1704 164759 3600
rect 880 1432 164759 1704
rect 880 1424 163900 1432
rect 105 1152 163900 1424
rect 105 307 164759 1152
<< metal4 >>
rect 4208 2128 4528 164336
rect 19568 2128 19888 164336
rect 34928 2128 35248 164336
rect 50288 2128 50608 164336
rect 65648 2128 65968 164336
rect 81008 2128 81328 164336
rect 96368 2128 96688 164336
rect 111728 2128 112048 164336
rect 127088 2128 127408 164336
rect 142448 2128 142768 164336
rect 157808 2128 158128 164336
<< obsm4 >>
rect 1163 2048 4128 156365
rect 4608 2048 19488 156365
rect 19968 2048 34848 156365
rect 35328 2048 50208 156365
rect 50688 2048 65568 156365
rect 66048 2048 80928 156365
rect 81408 2048 96288 156365
rect 96768 2048 111648 156365
rect 112128 2048 127008 156365
rect 127488 2048 142368 156365
rect 142848 2048 157728 156365
rect 158208 2048 163517 156365
rect 1163 579 163517 2048
<< labels >>
rlabel metal2 s 106922 166124 106978 166924 6 i_dout0[0]
port 1 nsew signal input
rlabel metal2 s 125414 166124 125470 166924 6 i_dout0[10]
port 2 nsew signal input
rlabel metal3 s 0 76984 800 77104 6 i_dout0[11]
port 3 nsew signal input
rlabel metal2 s 129094 166124 129150 166924 6 i_dout0[12]
port 4 nsew signal input
rlabel metal3 s 163980 91944 164780 92064 6 i_dout0[13]
port 5 nsew signal input
rlabel metal2 s 159454 0 159510 800 6 i_dout0[14]
port 6 nsew signal input
rlabel metal3 s 163980 104184 164780 104304 6 i_dout0[15]
port 7 nsew signal input
rlabel metal2 s 160374 0 160430 800 6 i_dout0[16]
port 8 nsew signal input
rlabel metal3 s 163980 109080 164780 109200 6 i_dout0[17]
port 9 nsew signal input
rlabel metal2 s 139306 166124 139362 166924 6 i_dout0[18]
port 10 nsew signal input
rlabel metal3 s 163980 119008 164780 119128 6 i_dout0[19]
port 11 nsew signal input
rlabel metal3 s 163980 8576 164780 8696 6 i_dout0[1]
port 12 nsew signal input
rlabel metal2 s 142066 166124 142122 166924 6 i_dout0[20]
port 13 nsew signal input
rlabel metal3 s 163980 126352 164780 126472 6 i_dout0[21]
port 14 nsew signal input
rlabel metal2 s 143906 166124 143962 166924 6 i_dout0[22]
port 15 nsew signal input
rlabel metal3 s 0 124176 800 124296 6 i_dout0[23]
port 16 nsew signal input
rlabel metal2 s 151358 166124 151414 166924 6 i_dout0[24]
port 17 nsew signal input
rlabel metal2 s 153198 166124 153254 166924 6 i_dout0[25]
port 18 nsew signal input
rlabel metal3 s 163980 150832 164780 150952 6 i_dout0[26]
port 19 nsew signal input
rlabel metal3 s 0 146208 800 146328 6 i_dout0[27]
port 20 nsew signal input
rlabel metal3 s 163980 153280 164780 153400 6 i_dout0[28]
port 21 nsew signal input
rlabel metal2 s 157798 166124 157854 166924 6 i_dout0[29]
port 22 nsew signal input
rlabel metal3 s 0 23536 800 23656 6 i_dout0[2]
port 23 nsew signal input
rlabel metal2 s 159638 166124 159694 166924 6 i_dout0[30]
port 24 nsew signal input
rlabel metal2 s 164238 166124 164294 166924 6 i_dout0[31]
port 25 nsew signal input
rlabel metal2 s 151910 0 151966 800 6 i_dout0[3]
port 26 nsew signal input
rlabel metal3 s 163980 45296 164780 45416 6 i_dout0[4]
port 27 nsew signal input
rlabel metal3 s 163980 52640 164780 52760 6 i_dout0[5]
port 28 nsew signal input
rlabel metal3 s 0 48696 800 48816 6 i_dout0[6]
port 29 nsew signal input
rlabel metal2 s 155222 0 155278 800 6 i_dout0[7]
port 30 nsew signal input
rlabel metal3 s 0 61208 800 61328 6 i_dout0[8]
port 31 nsew signal input
rlabel metal2 s 157338 0 157394 800 6 i_dout0[9]
port 32 nsew signal input
rlabel metal2 s 148322 0 148378 800 6 i_dout0_1[0]
port 33 nsew signal input
rlabel metal3 s 163980 79704 164780 79824 6 i_dout0_1[10]
port 34 nsew signal input
rlabel metal3 s 0 73856 800 73976 6 i_dout0_1[11]
port 35 nsew signal input
rlabel metal2 s 158810 0 158866 800 6 i_dout0_1[12]
port 36 nsew signal input
rlabel metal3 s 163980 89496 164780 89616 6 i_dout0_1[13]
port 37 nsew signal input
rlabel metal2 s 130014 166124 130070 166924 6 i_dout0_1[14]
port 38 nsew signal input
rlabel metal2 s 132774 166124 132830 166924 6 i_dout0_1[15]
port 39 nsew signal input
rlabel metal2 s 134614 166124 134670 166924 6 i_dout0_1[16]
port 40 nsew signal input
rlabel metal3 s 0 105272 800 105392 6 i_dout0_1[17]
port 41 nsew signal input
rlabel metal2 s 137466 166124 137522 166924 6 i_dout0_1[18]
port 42 nsew signal input
rlabel metal3 s 163980 114112 164780 114232 6 i_dout0_1[19]
port 43 nsew signal input
rlabel metal2 s 110602 166124 110658 166924 6 i_dout0_1[1]
port 44 nsew signal input
rlabel metal3 s 0 114792 800 114912 6 i_dout0_1[20]
port 45 nsew signal input
rlabel metal2 s 161846 0 161902 800 6 i_dout0_1[21]
port 46 nsew signal input
rlabel metal2 s 162122 0 162178 800 6 i_dout0_1[22]
port 47 nsew signal input
rlabel metal2 s 147586 166124 147642 166924 6 i_dout0_1[23]
port 48 nsew signal input
rlabel metal2 s 150438 166124 150494 166924 6 i_dout0_1[24]
port 49 nsew signal input
rlabel metal3 s 163980 145936 164780 146056 6 i_dout0_1[25]
port 50 nsew signal input
rlabel metal3 s 0 136824 800 136944 6 i_dout0_1[26]
port 51 nsew signal input
rlabel metal2 s 163318 0 163374 800 6 i_dout0_1[27]
port 52 nsew signal input
rlabel metal3 s 0 152600 800 152720 6 i_dout0_1[28]
port 53 nsew signal input
rlabel metal3 s 0 155728 800 155848 6 i_dout0_1[29]
port 54 nsew signal input
rlabel metal2 s 113362 166124 113418 166924 6 i_dout0_1[2]
port 55 nsew signal input
rlabel metal3 s 0 158856 800 158976 6 i_dout0_1[30]
port 56 nsew signal input
rlabel metal2 s 162398 166124 162454 166924 6 i_dout0_1[31]
port 57 nsew signal input
rlabel metal2 s 151634 0 151690 800 6 i_dout0_1[3]
port 58 nsew signal input
rlabel metal3 s 163980 42848 164780 42968 6 i_dout0_1[4]
port 59 nsew signal input
rlabel metal2 s 153198 0 153254 800 6 i_dout0_1[5]
port 60 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 i_dout0_1[6]
port 61 nsew signal input
rlabel metal2 s 154946 0 155002 800 6 i_dout0_1[7]
port 62 nsew signal input
rlabel metal2 s 123574 166124 123630 166924 6 i_dout0_1[8]
port 63 nsew signal input
rlabel metal3 s 0 64472 800 64592 6 i_dout0_1[9]
port 64 nsew signal input
rlabel metal3 s 0 1504 800 1624 6 i_dout1[0]
port 65 nsew signal input
rlabel metal2 s 126334 166124 126390 166924 6 i_dout1[10]
port 66 nsew signal input
rlabel metal2 s 158258 0 158314 800 6 i_dout1[11]
port 67 nsew signal input
rlabel metal3 s 163980 84600 164780 84720 6 i_dout1[12]
port 68 nsew signal input
rlabel metal3 s 163980 94392 164780 94512 6 i_dout1[13]
port 69 nsew signal input
rlabel metal2 s 130934 166124 130990 166924 6 i_dout1[14]
port 70 nsew signal input
rlabel metal3 s 0 92760 800 92880 6 i_dout1[15]
port 71 nsew signal input
rlabel metal3 s 0 99016 800 99136 6 i_dout1[16]
port 72 nsew signal input
rlabel metal3 s 163980 111528 164780 111648 6 i_dout1[17]
port 73 nsew signal input
rlabel metal3 s 0 108536 800 108656 6 i_dout1[18]
port 74 nsew signal input
rlabel metal3 s 163980 121456 164780 121576 6 i_dout1[19]
port 75 nsew signal input
rlabel metal3 s 163980 13472 164780 13592 6 i_dout1[1]
port 76 nsew signal input
rlabel metal3 s 0 121048 800 121168 6 i_dout1[20]
port 77 nsew signal input
rlabel metal3 s 163980 128800 164780 128920 6 i_dout1[21]
port 78 nsew signal input
rlabel metal2 s 144826 166124 144882 166924 6 i_dout1[22]
port 79 nsew signal input
rlabel metal3 s 163980 136144 164780 136264 6 i_dout1[23]
port 80 nsew signal input
rlabel metal2 s 152278 166124 152334 166924 6 i_dout1[24]
port 81 nsew signal input
rlabel metal3 s 0 133696 800 133816 6 i_dout1[25]
port 82 nsew signal input
rlabel metal3 s 0 139952 800 140072 6 i_dout1[26]
port 83 nsew signal input
rlabel metal2 s 155038 166124 155094 166924 6 i_dout1[27]
port 84 nsew signal input
rlabel metal3 s 163980 155728 164780 155848 6 i_dout1[28]
port 85 nsew signal input
rlabel metal2 s 164238 0 164294 800 6 i_dout1[29]
port 86 nsew signal input
rlabel metal3 s 163980 20816 164780 20936 6 i_dout1[2]
port 87 nsew signal input
rlabel metal2 s 160558 166124 160614 166924 6 i_dout1[30]
port 88 nsew signal input
rlabel metal3 s 0 161984 800 162104 6 i_dout1[31]
port 89 nsew signal input
rlabel metal2 s 114282 166124 114338 166924 6 i_dout1[3]
port 90 nsew signal input
rlabel metal3 s 163980 47744 164780 47864 6 i_dout1[4]
port 91 nsew signal input
rlabel metal3 s 163980 55088 164780 55208 6 i_dout1[5]
port 92 nsew signal input
rlabel metal2 s 119802 166124 119858 166924 6 i_dout1[6]
port 93 nsew signal input
rlabel metal3 s 0 51824 800 51944 6 i_dout1[7]
port 94 nsew signal input
rlabel metal2 s 156142 0 156198 800 6 i_dout1[8]
port 95 nsew signal input
rlabel metal3 s 0 70728 800 70848 6 i_dout1[9]
port 96 nsew signal input
rlabel metal2 s 148690 0 148746 800 6 i_dout1_1[0]
port 97 nsew signal input
rlabel metal3 s 163980 82152 164780 82272 6 i_dout1_1[10]
port 98 nsew signal input
rlabel metal2 s 128174 166124 128230 166924 6 i_dout1_1[11]
port 99 nsew signal input
rlabel metal3 s 0 83240 800 83360 6 i_dout1_1[12]
port 100 nsew signal input
rlabel metal3 s 0 86504 800 86624 6 i_dout1_1[13]
port 101 nsew signal input
rlabel metal3 s 163980 99288 164780 99408 6 i_dout1_1[14]
port 102 nsew signal input
rlabel metal2 s 159730 0 159786 800 6 i_dout1_1[15]
port 103 nsew signal input
rlabel metal2 s 160006 0 160062 800 6 i_dout1_1[16]
port 104 nsew signal input
rlabel metal3 s 163980 106632 164780 106752 6 i_dout1_1[17]
port 105 nsew signal input
rlabel metal2 s 138386 166124 138442 166924 6 i_dout1_1[18]
port 106 nsew signal input
rlabel metal3 s 163980 116560 164780 116680 6 i_dout1_1[19]
port 107 nsew signal input
rlabel metal3 s 163980 11024 164780 11144 6 i_dout1_1[1]
port 108 nsew signal input
rlabel metal3 s 0 117920 800 118040 6 i_dout1_1[20]
port 109 nsew signal input
rlabel metal3 s 163980 123904 164780 124024 6 i_dout1_1[21]
port 110 nsew signal input
rlabel metal3 s 163980 133696 164780 133816 6 i_dout1_1[22]
port 111 nsew signal input
rlabel metal2 s 148506 166124 148562 166924 6 i_dout1_1[23]
port 112 nsew signal input
rlabel metal3 s 163980 138592 164780 138712 6 i_dout1_1[24]
port 113 nsew signal input
rlabel metal3 s 0 130568 800 130688 6 i_dout1_1[25]
port 114 nsew signal input
rlabel metal2 s 162766 0 162822 800 6 i_dout1_1[26]
port 115 nsew signal input
rlabel metal2 s 154118 166124 154174 166924 6 i_dout1_1[27]
port 116 nsew signal input
rlabel metal2 s 163962 0 164018 800 6 i_dout1_1[28]
port 117 nsew signal input
rlabel metal2 s 156878 166124 156934 166924 6 i_dout1_1[29]
port 118 nsew signal input
rlabel metal3 s 0 20272 800 20392 6 i_dout1_1[2]
port 119 nsew signal input
rlabel metal2 s 158718 166124 158774 166924 6 i_dout1_1[30]
port 120 nsew signal input
rlabel metal2 s 163318 166124 163374 166924 6 i_dout1_1[31]
port 121 nsew signal input
rlabel metal3 s 163980 28160 164780 28280 6 i_dout1_1[3]
port 122 nsew signal input
rlabel metal3 s 0 32920 800 33040 6 i_dout1_1[4]
port 123 nsew signal input
rlabel metal3 s 0 39176 800 39296 6 i_dout1_1[5]
port 124 nsew signal input
rlabel metal3 s 163980 60120 164780 60240 6 i_dout1_1[6]
port 125 nsew signal input
rlabel metal2 s 122654 166124 122710 166924 6 i_dout1_1[7]
port 126 nsew signal input
rlabel metal3 s 0 58080 800 58200 6 i_dout1_1[8]
port 127 nsew signal input
rlabel metal3 s 0 67600 800 67720 6 i_dout1_1[9]
port 128 nsew signal input
rlabel metal2 s 478 166124 534 166924 6 io_in[0]
port 129 nsew signal input
rlabel metal2 s 28170 166124 28226 166924 6 io_in[10]
port 130 nsew signal input
rlabel metal2 s 31022 166124 31078 166924 6 io_in[11]
port 131 nsew signal input
rlabel metal2 s 33782 166124 33838 166924 6 io_in[12]
port 132 nsew signal input
rlabel metal2 s 36542 166124 36598 166924 6 io_in[13]
port 133 nsew signal input
rlabel metal2 s 39302 166124 39358 166924 6 io_in[14]
port 134 nsew signal input
rlabel metal2 s 42062 166124 42118 166924 6 io_in[15]
port 135 nsew signal input
rlabel metal2 s 44822 166124 44878 166924 6 io_in[16]
port 136 nsew signal input
rlabel metal2 s 47674 166124 47730 166924 6 io_in[17]
port 137 nsew signal input
rlabel metal2 s 50434 166124 50490 166924 6 io_in[18]
port 138 nsew signal input
rlabel metal2 s 53194 166124 53250 166924 6 io_in[19]
port 139 nsew signal input
rlabel metal2 s 3238 166124 3294 166924 6 io_in[1]
port 140 nsew signal input
rlabel metal2 s 55954 166124 56010 166924 6 io_in[20]
port 141 nsew signal input
rlabel metal2 s 58714 166124 58770 166924 6 io_in[21]
port 142 nsew signal input
rlabel metal2 s 61566 166124 61622 166924 6 io_in[22]
port 143 nsew signal input
rlabel metal2 s 64326 166124 64382 166924 6 io_in[23]
port 144 nsew signal input
rlabel metal2 s 67086 166124 67142 166924 6 io_in[24]
port 145 nsew signal input
rlabel metal2 s 69846 166124 69902 166924 6 io_in[25]
port 146 nsew signal input
rlabel metal2 s 72606 166124 72662 166924 6 io_in[26]
port 147 nsew signal input
rlabel metal2 s 75458 166124 75514 166924 6 io_in[27]
port 148 nsew signal input
rlabel metal2 s 78218 166124 78274 166924 6 io_in[28]
port 149 nsew signal input
rlabel metal2 s 80978 166124 81034 166924 6 io_in[29]
port 150 nsew signal input
rlabel metal2 s 5998 166124 6054 166924 6 io_in[2]
port 151 nsew signal input
rlabel metal2 s 83738 166124 83794 166924 6 io_in[30]
port 152 nsew signal input
rlabel metal2 s 86498 166124 86554 166924 6 io_in[31]
port 153 nsew signal input
rlabel metal2 s 89258 166124 89314 166924 6 io_in[32]
port 154 nsew signal input
rlabel metal2 s 92110 166124 92166 166924 6 io_in[33]
port 155 nsew signal input
rlabel metal2 s 94870 166124 94926 166924 6 io_in[34]
port 156 nsew signal input
rlabel metal2 s 97630 166124 97686 166924 6 io_in[35]
port 157 nsew signal input
rlabel metal2 s 100390 166124 100446 166924 6 io_in[36]
port 158 nsew signal input
rlabel metal2 s 103150 166124 103206 166924 6 io_in[37]
port 159 nsew signal input
rlabel metal2 s 8758 166124 8814 166924 6 io_in[3]
port 160 nsew signal input
rlabel metal2 s 11518 166124 11574 166924 6 io_in[4]
port 161 nsew signal input
rlabel metal2 s 14278 166124 14334 166924 6 io_in[5]
port 162 nsew signal input
rlabel metal2 s 17130 166124 17186 166924 6 io_in[6]
port 163 nsew signal input
rlabel metal2 s 19890 166124 19946 166924 6 io_in[7]
port 164 nsew signal input
rlabel metal2 s 22650 166124 22706 166924 6 io_in[8]
port 165 nsew signal input
rlabel metal2 s 25410 166124 25466 166924 6 io_in[9]
port 166 nsew signal input
rlabel metal2 s 1398 166124 1454 166924 6 io_oeb[0]
port 167 nsew signal output
rlabel metal2 s 29090 166124 29146 166924 6 io_oeb[10]
port 168 nsew signal output
rlabel metal2 s 31942 166124 31998 166924 6 io_oeb[11]
port 169 nsew signal output
rlabel metal2 s 34702 166124 34758 166924 6 io_oeb[12]
port 170 nsew signal output
rlabel metal2 s 37462 166124 37518 166924 6 io_oeb[13]
port 171 nsew signal output
rlabel metal2 s 40222 166124 40278 166924 6 io_oeb[14]
port 172 nsew signal output
rlabel metal2 s 42982 166124 43038 166924 6 io_oeb[15]
port 173 nsew signal output
rlabel metal2 s 45834 166124 45890 166924 6 io_oeb[16]
port 174 nsew signal output
rlabel metal2 s 48594 166124 48650 166924 6 io_oeb[17]
port 175 nsew signal output
rlabel metal2 s 51354 166124 51410 166924 6 io_oeb[18]
port 176 nsew signal output
rlabel metal2 s 54114 166124 54170 166924 6 io_oeb[19]
port 177 nsew signal output
rlabel metal2 s 4158 166124 4214 166924 6 io_oeb[1]
port 178 nsew signal output
rlabel metal2 s 56874 166124 56930 166924 6 io_oeb[20]
port 179 nsew signal output
rlabel metal2 s 59634 166124 59690 166924 6 io_oeb[21]
port 180 nsew signal output
rlabel metal2 s 62486 166124 62542 166924 6 io_oeb[22]
port 181 nsew signal output
rlabel metal2 s 65246 166124 65302 166924 6 io_oeb[23]
port 182 nsew signal output
rlabel metal2 s 68006 166124 68062 166924 6 io_oeb[24]
port 183 nsew signal output
rlabel metal2 s 70766 166124 70822 166924 6 io_oeb[25]
port 184 nsew signal output
rlabel metal2 s 73526 166124 73582 166924 6 io_oeb[26]
port 185 nsew signal output
rlabel metal2 s 76378 166124 76434 166924 6 io_oeb[27]
port 186 nsew signal output
rlabel metal2 s 79138 166124 79194 166924 6 io_oeb[28]
port 187 nsew signal output
rlabel metal2 s 81898 166124 81954 166924 6 io_oeb[29]
port 188 nsew signal output
rlabel metal2 s 6918 166124 6974 166924 6 io_oeb[2]
port 189 nsew signal output
rlabel metal2 s 84658 166124 84714 166924 6 io_oeb[30]
port 190 nsew signal output
rlabel metal2 s 87418 166124 87474 166924 6 io_oeb[31]
port 191 nsew signal output
rlabel metal2 s 90178 166124 90234 166924 6 io_oeb[32]
port 192 nsew signal output
rlabel metal2 s 93030 166124 93086 166924 6 io_oeb[33]
port 193 nsew signal output
rlabel metal2 s 95790 166124 95846 166924 6 io_oeb[34]
port 194 nsew signal output
rlabel metal2 s 98550 166124 98606 166924 6 io_oeb[35]
port 195 nsew signal output
rlabel metal2 s 101310 166124 101366 166924 6 io_oeb[36]
port 196 nsew signal output
rlabel metal2 s 104070 166124 104126 166924 6 io_oeb[37]
port 197 nsew signal output
rlabel metal2 s 9678 166124 9734 166924 6 io_oeb[3]
port 198 nsew signal output
rlabel metal2 s 12438 166124 12494 166924 6 io_oeb[4]
port 199 nsew signal output
rlabel metal2 s 15198 166124 15254 166924 6 io_oeb[5]
port 200 nsew signal output
rlabel metal2 s 18050 166124 18106 166924 6 io_oeb[6]
port 201 nsew signal output
rlabel metal2 s 20810 166124 20866 166924 6 io_oeb[7]
port 202 nsew signal output
rlabel metal2 s 23570 166124 23626 166924 6 io_oeb[8]
port 203 nsew signal output
rlabel metal2 s 26330 166124 26386 166924 6 io_oeb[9]
port 204 nsew signal output
rlabel metal2 s 2318 166124 2374 166924 6 io_out[0]
port 205 nsew signal output
rlabel metal2 s 30010 166124 30066 166924 6 io_out[10]
port 206 nsew signal output
rlabel metal2 s 32862 166124 32918 166924 6 io_out[11]
port 207 nsew signal output
rlabel metal2 s 35622 166124 35678 166924 6 io_out[12]
port 208 nsew signal output
rlabel metal2 s 38382 166124 38438 166924 6 io_out[13]
port 209 nsew signal output
rlabel metal2 s 41142 166124 41198 166924 6 io_out[14]
port 210 nsew signal output
rlabel metal2 s 43902 166124 43958 166924 6 io_out[15]
port 211 nsew signal output
rlabel metal2 s 46754 166124 46810 166924 6 io_out[16]
port 212 nsew signal output
rlabel metal2 s 49514 166124 49570 166924 6 io_out[17]
port 213 nsew signal output
rlabel metal2 s 52274 166124 52330 166924 6 io_out[18]
port 214 nsew signal output
rlabel metal2 s 55034 166124 55090 166924 6 io_out[19]
port 215 nsew signal output
rlabel metal2 s 5078 166124 5134 166924 6 io_out[1]
port 216 nsew signal output
rlabel metal2 s 57794 166124 57850 166924 6 io_out[20]
port 217 nsew signal output
rlabel metal2 s 60646 166124 60702 166924 6 io_out[21]
port 218 nsew signal output
rlabel metal2 s 63406 166124 63462 166924 6 io_out[22]
port 219 nsew signal output
rlabel metal2 s 66166 166124 66222 166924 6 io_out[23]
port 220 nsew signal output
rlabel metal2 s 68926 166124 68982 166924 6 io_out[24]
port 221 nsew signal output
rlabel metal2 s 71686 166124 71742 166924 6 io_out[25]
port 222 nsew signal output
rlabel metal2 s 74446 166124 74502 166924 6 io_out[26]
port 223 nsew signal output
rlabel metal2 s 77298 166124 77354 166924 6 io_out[27]
port 224 nsew signal output
rlabel metal2 s 80058 166124 80114 166924 6 io_out[28]
port 225 nsew signal output
rlabel metal2 s 82818 166124 82874 166924 6 io_out[29]
port 226 nsew signal output
rlabel metal2 s 7838 166124 7894 166924 6 io_out[2]
port 227 nsew signal output
rlabel metal2 s 85578 166124 85634 166924 6 io_out[30]
port 228 nsew signal output
rlabel metal2 s 88338 166124 88394 166924 6 io_out[31]
port 229 nsew signal output
rlabel metal2 s 91190 166124 91246 166924 6 io_out[32]
port 230 nsew signal output
rlabel metal2 s 93950 166124 94006 166924 6 io_out[33]
port 231 nsew signal output
rlabel metal2 s 96710 166124 96766 166924 6 io_out[34]
port 232 nsew signal output
rlabel metal2 s 99470 166124 99526 166924 6 io_out[35]
port 233 nsew signal output
rlabel metal2 s 102230 166124 102286 166924 6 io_out[36]
port 234 nsew signal output
rlabel metal2 s 104990 166124 105046 166924 6 io_out[37]
port 235 nsew signal output
rlabel metal2 s 10598 166124 10654 166924 6 io_out[3]
port 236 nsew signal output
rlabel metal2 s 13358 166124 13414 166924 6 io_out[4]
port 237 nsew signal output
rlabel metal2 s 16210 166124 16266 166924 6 io_out[5]
port 238 nsew signal output
rlabel metal2 s 18970 166124 19026 166924 6 io_out[6]
port 239 nsew signal output
rlabel metal2 s 21730 166124 21786 166924 6 io_out[7]
port 240 nsew signal output
rlabel metal2 s 24490 166124 24546 166924 6 io_out[8]
port 241 nsew signal output
rlabel metal2 s 27250 166124 27306 166924 6 io_out[9]
port 242 nsew signal output
rlabel metal2 s 146850 0 146906 800 6 irq[0]
port 243 nsew signal output
rlabel metal2 s 147126 0 147182 800 6 irq[1]
port 244 nsew signal output
rlabel metal2 s 147494 0 147550 800 6 irq[2]
port 245 nsew signal output
rlabel metal2 s 31850 0 31906 800 6 la_data_in[0]
port 246 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 la_data_in[100]
port 247 nsew signal input
rlabel metal2 s 122562 0 122618 800 6 la_data_in[101]
port 248 nsew signal input
rlabel metal2 s 123482 0 123538 800 6 la_data_in[102]
port 249 nsew signal input
rlabel metal2 s 124402 0 124458 800 6 la_data_in[103]
port 250 nsew signal input
rlabel metal2 s 125322 0 125378 800 6 la_data_in[104]
port 251 nsew signal input
rlabel metal2 s 126150 0 126206 800 6 la_data_in[105]
port 252 nsew signal input
rlabel metal2 s 127070 0 127126 800 6 la_data_in[106]
port 253 nsew signal input
rlabel metal2 s 127990 0 128046 800 6 la_data_in[107]
port 254 nsew signal input
rlabel metal2 s 128910 0 128966 800 6 la_data_in[108]
port 255 nsew signal input
rlabel metal2 s 129830 0 129886 800 6 la_data_in[109]
port 256 nsew signal input
rlabel metal2 s 40774 0 40830 800 6 la_data_in[10]
port 257 nsew signal input
rlabel metal2 s 130658 0 130714 800 6 la_data_in[110]
port 258 nsew signal input
rlabel metal2 s 131578 0 131634 800 6 la_data_in[111]
port 259 nsew signal input
rlabel metal2 s 132498 0 132554 800 6 la_data_in[112]
port 260 nsew signal input
rlabel metal2 s 133418 0 133474 800 6 la_data_in[113]
port 261 nsew signal input
rlabel metal2 s 134246 0 134302 800 6 la_data_in[114]
port 262 nsew signal input
rlabel metal2 s 135166 0 135222 800 6 la_data_in[115]
port 263 nsew signal input
rlabel metal2 s 136086 0 136142 800 6 la_data_in[116]
port 264 nsew signal input
rlabel metal2 s 137006 0 137062 800 6 la_data_in[117]
port 265 nsew signal input
rlabel metal2 s 137834 0 137890 800 6 la_data_in[118]
port 266 nsew signal input
rlabel metal2 s 138754 0 138810 800 6 la_data_in[119]
port 267 nsew signal input
rlabel metal2 s 41694 0 41750 800 6 la_data_in[11]
port 268 nsew signal input
rlabel metal2 s 139674 0 139730 800 6 la_data_in[120]
port 269 nsew signal input
rlabel metal2 s 140594 0 140650 800 6 la_data_in[121]
port 270 nsew signal input
rlabel metal2 s 141514 0 141570 800 6 la_data_in[122]
port 271 nsew signal input
rlabel metal2 s 142342 0 142398 800 6 la_data_in[123]
port 272 nsew signal input
rlabel metal2 s 143262 0 143318 800 6 la_data_in[124]
port 273 nsew signal input
rlabel metal2 s 144182 0 144238 800 6 la_data_in[125]
port 274 nsew signal input
rlabel metal2 s 145102 0 145158 800 6 la_data_in[126]
port 275 nsew signal input
rlabel metal2 s 145930 0 145986 800 6 la_data_in[127]
port 276 nsew signal input
rlabel metal2 s 42614 0 42670 800 6 la_data_in[12]
port 277 nsew signal input
rlabel metal2 s 43534 0 43590 800 6 la_data_in[13]
port 278 nsew signal input
rlabel metal2 s 44362 0 44418 800 6 la_data_in[14]
port 279 nsew signal input
rlabel metal2 s 45282 0 45338 800 6 la_data_in[15]
port 280 nsew signal input
rlabel metal2 s 46202 0 46258 800 6 la_data_in[16]
port 281 nsew signal input
rlabel metal2 s 47122 0 47178 800 6 la_data_in[17]
port 282 nsew signal input
rlabel metal2 s 48042 0 48098 800 6 la_data_in[18]
port 283 nsew signal input
rlabel metal2 s 48870 0 48926 800 6 la_data_in[19]
port 284 nsew signal input
rlabel metal2 s 32678 0 32734 800 6 la_data_in[1]
port 285 nsew signal input
rlabel metal2 s 49790 0 49846 800 6 la_data_in[20]
port 286 nsew signal input
rlabel metal2 s 50710 0 50766 800 6 la_data_in[21]
port 287 nsew signal input
rlabel metal2 s 51630 0 51686 800 6 la_data_in[22]
port 288 nsew signal input
rlabel metal2 s 52458 0 52514 800 6 la_data_in[23]
port 289 nsew signal input
rlabel metal2 s 53378 0 53434 800 6 la_data_in[24]
port 290 nsew signal input
rlabel metal2 s 54298 0 54354 800 6 la_data_in[25]
port 291 nsew signal input
rlabel metal2 s 55218 0 55274 800 6 la_data_in[26]
port 292 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 la_data_in[27]
port 293 nsew signal input
rlabel metal2 s 56966 0 57022 800 6 la_data_in[28]
port 294 nsew signal input
rlabel metal2 s 57886 0 57942 800 6 la_data_in[29]
port 295 nsew signal input
rlabel metal2 s 33598 0 33654 800 6 la_data_in[2]
port 296 nsew signal input
rlabel metal2 s 58806 0 58862 800 6 la_data_in[30]
port 297 nsew signal input
rlabel metal2 s 59726 0 59782 800 6 la_data_in[31]
port 298 nsew signal input
rlabel metal2 s 60554 0 60610 800 6 la_data_in[32]
port 299 nsew signal input
rlabel metal2 s 61474 0 61530 800 6 la_data_in[33]
port 300 nsew signal input
rlabel metal2 s 62394 0 62450 800 6 la_data_in[34]
port 301 nsew signal input
rlabel metal2 s 63314 0 63370 800 6 la_data_in[35]
port 302 nsew signal input
rlabel metal2 s 64142 0 64198 800 6 la_data_in[36]
port 303 nsew signal input
rlabel metal2 s 65062 0 65118 800 6 la_data_in[37]
port 304 nsew signal input
rlabel metal2 s 65982 0 66038 800 6 la_data_in[38]
port 305 nsew signal input
rlabel metal2 s 66902 0 66958 800 6 la_data_in[39]
port 306 nsew signal input
rlabel metal2 s 34518 0 34574 800 6 la_data_in[3]
port 307 nsew signal input
rlabel metal2 s 67730 0 67786 800 6 la_data_in[40]
port 308 nsew signal input
rlabel metal2 s 68650 0 68706 800 6 la_data_in[41]
port 309 nsew signal input
rlabel metal2 s 69570 0 69626 800 6 la_data_in[42]
port 310 nsew signal input
rlabel metal2 s 70490 0 70546 800 6 la_data_in[43]
port 311 nsew signal input
rlabel metal2 s 71410 0 71466 800 6 la_data_in[44]
port 312 nsew signal input
rlabel metal2 s 72238 0 72294 800 6 la_data_in[45]
port 313 nsew signal input
rlabel metal2 s 73158 0 73214 800 6 la_data_in[46]
port 314 nsew signal input
rlabel metal2 s 74078 0 74134 800 6 la_data_in[47]
port 315 nsew signal input
rlabel metal2 s 74998 0 75054 800 6 la_data_in[48]
port 316 nsew signal input
rlabel metal2 s 75826 0 75882 800 6 la_data_in[49]
port 317 nsew signal input
rlabel metal2 s 35438 0 35494 800 6 la_data_in[4]
port 318 nsew signal input
rlabel metal2 s 76746 0 76802 800 6 la_data_in[50]
port 319 nsew signal input
rlabel metal2 s 77666 0 77722 800 6 la_data_in[51]
port 320 nsew signal input
rlabel metal2 s 78586 0 78642 800 6 la_data_in[52]
port 321 nsew signal input
rlabel metal2 s 79414 0 79470 800 6 la_data_in[53]
port 322 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 la_data_in[54]
port 323 nsew signal input
rlabel metal2 s 81254 0 81310 800 6 la_data_in[55]
port 324 nsew signal input
rlabel metal2 s 82174 0 82230 800 6 la_data_in[56]
port 325 nsew signal input
rlabel metal2 s 83094 0 83150 800 6 la_data_in[57]
port 326 nsew signal input
rlabel metal2 s 83922 0 83978 800 6 la_data_in[58]
port 327 nsew signal input
rlabel metal2 s 84842 0 84898 800 6 la_data_in[59]
port 328 nsew signal input
rlabel metal2 s 36358 0 36414 800 6 la_data_in[5]
port 329 nsew signal input
rlabel metal2 s 85762 0 85818 800 6 la_data_in[60]
port 330 nsew signal input
rlabel metal2 s 86682 0 86738 800 6 la_data_in[61]
port 331 nsew signal input
rlabel metal2 s 87510 0 87566 800 6 la_data_in[62]
port 332 nsew signal input
rlabel metal2 s 88430 0 88486 800 6 la_data_in[63]
port 333 nsew signal input
rlabel metal2 s 89350 0 89406 800 6 la_data_in[64]
port 334 nsew signal input
rlabel metal2 s 90270 0 90326 800 6 la_data_in[65]
port 335 nsew signal input
rlabel metal2 s 91098 0 91154 800 6 la_data_in[66]
port 336 nsew signal input
rlabel metal2 s 92018 0 92074 800 6 la_data_in[67]
port 337 nsew signal input
rlabel metal2 s 92938 0 92994 800 6 la_data_in[68]
port 338 nsew signal input
rlabel metal2 s 93858 0 93914 800 6 la_data_in[69]
port 339 nsew signal input
rlabel metal2 s 37186 0 37242 800 6 la_data_in[6]
port 340 nsew signal input
rlabel metal2 s 94778 0 94834 800 6 la_data_in[70]
port 341 nsew signal input
rlabel metal2 s 95606 0 95662 800 6 la_data_in[71]
port 342 nsew signal input
rlabel metal2 s 96526 0 96582 800 6 la_data_in[72]
port 343 nsew signal input
rlabel metal2 s 97446 0 97502 800 6 la_data_in[73]
port 344 nsew signal input
rlabel metal2 s 98366 0 98422 800 6 la_data_in[74]
port 345 nsew signal input
rlabel metal2 s 99194 0 99250 800 6 la_data_in[75]
port 346 nsew signal input
rlabel metal2 s 100114 0 100170 800 6 la_data_in[76]
port 347 nsew signal input
rlabel metal2 s 101034 0 101090 800 6 la_data_in[77]
port 348 nsew signal input
rlabel metal2 s 101954 0 102010 800 6 la_data_in[78]
port 349 nsew signal input
rlabel metal2 s 102782 0 102838 800 6 la_data_in[79]
port 350 nsew signal input
rlabel metal2 s 38106 0 38162 800 6 la_data_in[7]
port 351 nsew signal input
rlabel metal2 s 103702 0 103758 800 6 la_data_in[80]
port 352 nsew signal input
rlabel metal2 s 104622 0 104678 800 6 la_data_in[81]
port 353 nsew signal input
rlabel metal2 s 105542 0 105598 800 6 la_data_in[82]
port 354 nsew signal input
rlabel metal2 s 106462 0 106518 800 6 la_data_in[83]
port 355 nsew signal input
rlabel metal2 s 107290 0 107346 800 6 la_data_in[84]
port 356 nsew signal input
rlabel metal2 s 108210 0 108266 800 6 la_data_in[85]
port 357 nsew signal input
rlabel metal2 s 109130 0 109186 800 6 la_data_in[86]
port 358 nsew signal input
rlabel metal2 s 110050 0 110106 800 6 la_data_in[87]
port 359 nsew signal input
rlabel metal2 s 110878 0 110934 800 6 la_data_in[88]
port 360 nsew signal input
rlabel metal2 s 111798 0 111854 800 6 la_data_in[89]
port 361 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 la_data_in[8]
port 362 nsew signal input
rlabel metal2 s 112718 0 112774 800 6 la_data_in[90]
port 363 nsew signal input
rlabel metal2 s 113638 0 113694 800 6 la_data_in[91]
port 364 nsew signal input
rlabel metal2 s 114466 0 114522 800 6 la_data_in[92]
port 365 nsew signal input
rlabel metal2 s 115386 0 115442 800 6 la_data_in[93]
port 366 nsew signal input
rlabel metal2 s 116306 0 116362 800 6 la_data_in[94]
port 367 nsew signal input
rlabel metal2 s 117226 0 117282 800 6 la_data_in[95]
port 368 nsew signal input
rlabel metal2 s 118146 0 118202 800 6 la_data_in[96]
port 369 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 la_data_in[97]
port 370 nsew signal input
rlabel metal2 s 119894 0 119950 800 6 la_data_in[98]
port 371 nsew signal input
rlabel metal2 s 120814 0 120870 800 6 la_data_in[99]
port 372 nsew signal input
rlabel metal2 s 39946 0 40002 800 6 la_data_in[9]
port 373 nsew signal input
rlabel metal2 s 32126 0 32182 800 6 la_data_out[0]
port 374 nsew signal output
rlabel metal2 s 122010 0 122066 800 6 la_data_out[100]
port 375 nsew signal output
rlabel metal2 s 122930 0 122986 800 6 la_data_out[101]
port 376 nsew signal output
rlabel metal2 s 123758 0 123814 800 6 la_data_out[102]
port 377 nsew signal output
rlabel metal2 s 124678 0 124734 800 6 la_data_out[103]
port 378 nsew signal output
rlabel metal2 s 125598 0 125654 800 6 la_data_out[104]
port 379 nsew signal output
rlabel metal2 s 126518 0 126574 800 6 la_data_out[105]
port 380 nsew signal output
rlabel metal2 s 127346 0 127402 800 6 la_data_out[106]
port 381 nsew signal output
rlabel metal2 s 128266 0 128322 800 6 la_data_out[107]
port 382 nsew signal output
rlabel metal2 s 129186 0 129242 800 6 la_data_out[108]
port 383 nsew signal output
rlabel metal2 s 130106 0 130162 800 6 la_data_out[109]
port 384 nsew signal output
rlabel metal2 s 41142 0 41198 800 6 la_data_out[10]
port 385 nsew signal output
rlabel metal2 s 131026 0 131082 800 6 la_data_out[110]
port 386 nsew signal output
rlabel metal2 s 131854 0 131910 800 6 la_data_out[111]
port 387 nsew signal output
rlabel metal2 s 132774 0 132830 800 6 la_data_out[112]
port 388 nsew signal output
rlabel metal2 s 133694 0 133750 800 6 la_data_out[113]
port 389 nsew signal output
rlabel metal2 s 134614 0 134670 800 6 la_data_out[114]
port 390 nsew signal output
rlabel metal2 s 135442 0 135498 800 6 la_data_out[115]
port 391 nsew signal output
rlabel metal2 s 136362 0 136418 800 6 la_data_out[116]
port 392 nsew signal output
rlabel metal2 s 137282 0 137338 800 6 la_data_out[117]
port 393 nsew signal output
rlabel metal2 s 138202 0 138258 800 6 la_data_out[118]
port 394 nsew signal output
rlabel metal2 s 139030 0 139086 800 6 la_data_out[119]
port 395 nsew signal output
rlabel metal2 s 41970 0 42026 800 6 la_data_out[11]
port 396 nsew signal output
rlabel metal2 s 139950 0 140006 800 6 la_data_out[120]
port 397 nsew signal output
rlabel metal2 s 140870 0 140926 800 6 la_data_out[121]
port 398 nsew signal output
rlabel metal2 s 141790 0 141846 800 6 la_data_out[122]
port 399 nsew signal output
rlabel metal2 s 142710 0 142766 800 6 la_data_out[123]
port 400 nsew signal output
rlabel metal2 s 143538 0 143594 800 6 la_data_out[124]
port 401 nsew signal output
rlabel metal2 s 144458 0 144514 800 6 la_data_out[125]
port 402 nsew signal output
rlabel metal2 s 145378 0 145434 800 6 la_data_out[126]
port 403 nsew signal output
rlabel metal2 s 146298 0 146354 800 6 la_data_out[127]
port 404 nsew signal output
rlabel metal2 s 42890 0 42946 800 6 la_data_out[12]
port 405 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 la_data_out[13]
port 406 nsew signal output
rlabel metal2 s 44730 0 44786 800 6 la_data_out[14]
port 407 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 la_data_out[15]
port 408 nsew signal output
rlabel metal2 s 46478 0 46534 800 6 la_data_out[16]
port 409 nsew signal output
rlabel metal2 s 47398 0 47454 800 6 la_data_out[17]
port 410 nsew signal output
rlabel metal2 s 48318 0 48374 800 6 la_data_out[18]
port 411 nsew signal output
rlabel metal2 s 49238 0 49294 800 6 la_data_out[19]
port 412 nsew signal output
rlabel metal2 s 33046 0 33102 800 6 la_data_out[1]
port 413 nsew signal output
rlabel metal2 s 50066 0 50122 800 6 la_data_out[20]
port 414 nsew signal output
rlabel metal2 s 50986 0 51042 800 6 la_data_out[21]
port 415 nsew signal output
rlabel metal2 s 51906 0 51962 800 6 la_data_out[22]
port 416 nsew signal output
rlabel metal2 s 52826 0 52882 800 6 la_data_out[23]
port 417 nsew signal output
rlabel metal2 s 53654 0 53710 800 6 la_data_out[24]
port 418 nsew signal output
rlabel metal2 s 54574 0 54630 800 6 la_data_out[25]
port 419 nsew signal output
rlabel metal2 s 55494 0 55550 800 6 la_data_out[26]
port 420 nsew signal output
rlabel metal2 s 56414 0 56470 800 6 la_data_out[27]
port 421 nsew signal output
rlabel metal2 s 57242 0 57298 800 6 la_data_out[28]
port 422 nsew signal output
rlabel metal2 s 58162 0 58218 800 6 la_data_out[29]
port 423 nsew signal output
rlabel metal2 s 33874 0 33930 800 6 la_data_out[2]
port 424 nsew signal output
rlabel metal2 s 59082 0 59138 800 6 la_data_out[30]
port 425 nsew signal output
rlabel metal2 s 60002 0 60058 800 6 la_data_out[31]
port 426 nsew signal output
rlabel metal2 s 60922 0 60978 800 6 la_data_out[32]
port 427 nsew signal output
rlabel metal2 s 61750 0 61806 800 6 la_data_out[33]
port 428 nsew signal output
rlabel metal2 s 62670 0 62726 800 6 la_data_out[34]
port 429 nsew signal output
rlabel metal2 s 63590 0 63646 800 6 la_data_out[35]
port 430 nsew signal output
rlabel metal2 s 64510 0 64566 800 6 la_data_out[36]
port 431 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 la_data_out[37]
port 432 nsew signal output
rlabel metal2 s 66258 0 66314 800 6 la_data_out[38]
port 433 nsew signal output
rlabel metal2 s 67178 0 67234 800 6 la_data_out[39]
port 434 nsew signal output
rlabel metal2 s 34794 0 34850 800 6 la_data_out[3]
port 435 nsew signal output
rlabel metal2 s 68098 0 68154 800 6 la_data_out[40]
port 436 nsew signal output
rlabel metal2 s 68926 0 68982 800 6 la_data_out[41]
port 437 nsew signal output
rlabel metal2 s 69846 0 69902 800 6 la_data_out[42]
port 438 nsew signal output
rlabel metal2 s 70766 0 70822 800 6 la_data_out[43]
port 439 nsew signal output
rlabel metal2 s 71686 0 71742 800 6 la_data_out[44]
port 440 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 la_data_out[45]
port 441 nsew signal output
rlabel metal2 s 73434 0 73490 800 6 la_data_out[46]
port 442 nsew signal output
rlabel metal2 s 74354 0 74410 800 6 la_data_out[47]
port 443 nsew signal output
rlabel metal2 s 75274 0 75330 800 6 la_data_out[48]
port 444 nsew signal output
rlabel metal2 s 76194 0 76250 800 6 la_data_out[49]
port 445 nsew signal output
rlabel metal2 s 35714 0 35770 800 6 la_data_out[4]
port 446 nsew signal output
rlabel metal2 s 77022 0 77078 800 6 la_data_out[50]
port 447 nsew signal output
rlabel metal2 s 77942 0 77998 800 6 la_data_out[51]
port 448 nsew signal output
rlabel metal2 s 78862 0 78918 800 6 la_data_out[52]
port 449 nsew signal output
rlabel metal2 s 79782 0 79838 800 6 la_data_out[53]
port 450 nsew signal output
rlabel metal2 s 80610 0 80666 800 6 la_data_out[54]
port 451 nsew signal output
rlabel metal2 s 81530 0 81586 800 6 la_data_out[55]
port 452 nsew signal output
rlabel metal2 s 82450 0 82506 800 6 la_data_out[56]
port 453 nsew signal output
rlabel metal2 s 83370 0 83426 800 6 la_data_out[57]
port 454 nsew signal output
rlabel metal2 s 84290 0 84346 800 6 la_data_out[58]
port 455 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 la_data_out[59]
port 456 nsew signal output
rlabel metal2 s 36634 0 36690 800 6 la_data_out[5]
port 457 nsew signal output
rlabel metal2 s 86038 0 86094 800 6 la_data_out[60]
port 458 nsew signal output
rlabel metal2 s 86958 0 87014 800 6 la_data_out[61]
port 459 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 la_data_out[62]
port 460 nsew signal output
rlabel metal2 s 88706 0 88762 800 6 la_data_out[63]
port 461 nsew signal output
rlabel metal2 s 89626 0 89682 800 6 la_data_out[64]
port 462 nsew signal output
rlabel metal2 s 90546 0 90602 800 6 la_data_out[65]
port 463 nsew signal output
rlabel metal2 s 91466 0 91522 800 6 la_data_out[66]
port 464 nsew signal output
rlabel metal2 s 92294 0 92350 800 6 la_data_out[67]
port 465 nsew signal output
rlabel metal2 s 93214 0 93270 800 6 la_data_out[68]
port 466 nsew signal output
rlabel metal2 s 94134 0 94190 800 6 la_data_out[69]
port 467 nsew signal output
rlabel metal2 s 37554 0 37610 800 6 la_data_out[6]
port 468 nsew signal output
rlabel metal2 s 95054 0 95110 800 6 la_data_out[70]
port 469 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 la_data_out[71]
port 470 nsew signal output
rlabel metal2 s 96802 0 96858 800 6 la_data_out[72]
port 471 nsew signal output
rlabel metal2 s 97722 0 97778 800 6 la_data_out[73]
port 472 nsew signal output
rlabel metal2 s 98642 0 98698 800 6 la_data_out[74]
port 473 nsew signal output
rlabel metal2 s 99562 0 99618 800 6 la_data_out[75]
port 474 nsew signal output
rlabel metal2 s 100390 0 100446 800 6 la_data_out[76]
port 475 nsew signal output
rlabel metal2 s 101310 0 101366 800 6 la_data_out[77]
port 476 nsew signal output
rlabel metal2 s 102230 0 102286 800 6 la_data_out[78]
port 477 nsew signal output
rlabel metal2 s 103150 0 103206 800 6 la_data_out[79]
port 478 nsew signal output
rlabel metal2 s 38382 0 38438 800 6 la_data_out[7]
port 479 nsew signal output
rlabel metal2 s 103978 0 104034 800 6 la_data_out[80]
port 480 nsew signal output
rlabel metal2 s 104898 0 104954 800 6 la_data_out[81]
port 481 nsew signal output
rlabel metal2 s 105818 0 105874 800 6 la_data_out[82]
port 482 nsew signal output
rlabel metal2 s 106738 0 106794 800 6 la_data_out[83]
port 483 nsew signal output
rlabel metal2 s 107658 0 107714 800 6 la_data_out[84]
port 484 nsew signal output
rlabel metal2 s 108486 0 108542 800 6 la_data_out[85]
port 485 nsew signal output
rlabel metal2 s 109406 0 109462 800 6 la_data_out[86]
port 486 nsew signal output
rlabel metal2 s 110326 0 110382 800 6 la_data_out[87]
port 487 nsew signal output
rlabel metal2 s 111246 0 111302 800 6 la_data_out[88]
port 488 nsew signal output
rlabel metal2 s 112074 0 112130 800 6 la_data_out[89]
port 489 nsew signal output
rlabel metal2 s 39302 0 39358 800 6 la_data_out[8]
port 490 nsew signal output
rlabel metal2 s 112994 0 113050 800 6 la_data_out[90]
port 491 nsew signal output
rlabel metal2 s 113914 0 113970 800 6 la_data_out[91]
port 492 nsew signal output
rlabel metal2 s 114834 0 114890 800 6 la_data_out[92]
port 493 nsew signal output
rlabel metal2 s 115662 0 115718 800 6 la_data_out[93]
port 494 nsew signal output
rlabel metal2 s 116582 0 116638 800 6 la_data_out[94]
port 495 nsew signal output
rlabel metal2 s 117502 0 117558 800 6 la_data_out[95]
port 496 nsew signal output
rlabel metal2 s 118422 0 118478 800 6 la_data_out[96]
port 497 nsew signal output
rlabel metal2 s 119342 0 119398 800 6 la_data_out[97]
port 498 nsew signal output
rlabel metal2 s 120170 0 120226 800 6 la_data_out[98]
port 499 nsew signal output
rlabel metal2 s 121090 0 121146 800 6 la_data_out[99]
port 500 nsew signal output
rlabel metal2 s 40222 0 40278 800 6 la_data_out[9]
port 501 nsew signal output
rlabel metal2 s 32402 0 32458 800 6 la_oenb[0]
port 502 nsew signal input
rlabel metal2 s 122286 0 122342 800 6 la_oenb[100]
port 503 nsew signal input
rlabel metal2 s 123206 0 123262 800 6 la_oenb[101]
port 504 nsew signal input
rlabel metal2 s 124126 0 124182 800 6 la_oenb[102]
port 505 nsew signal input
rlabel metal2 s 124954 0 125010 800 6 la_oenb[103]
port 506 nsew signal input
rlabel metal2 s 125874 0 125930 800 6 la_oenb[104]
port 507 nsew signal input
rlabel metal2 s 126794 0 126850 800 6 la_oenb[105]
port 508 nsew signal input
rlabel metal2 s 127714 0 127770 800 6 la_oenb[106]
port 509 nsew signal input
rlabel metal2 s 128542 0 128598 800 6 la_oenb[107]
port 510 nsew signal input
rlabel metal2 s 129462 0 129518 800 6 la_oenb[108]
port 511 nsew signal input
rlabel metal2 s 130382 0 130438 800 6 la_oenb[109]
port 512 nsew signal input
rlabel metal2 s 41418 0 41474 800 6 la_oenb[10]
port 513 nsew signal input
rlabel metal2 s 131302 0 131358 800 6 la_oenb[110]
port 514 nsew signal input
rlabel metal2 s 132222 0 132278 800 6 la_oenb[111]
port 515 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 la_oenb[112]
port 516 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 la_oenb[113]
port 517 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 la_oenb[114]
port 518 nsew signal input
rlabel metal2 s 135810 0 135866 800 6 la_oenb[115]
port 519 nsew signal input
rlabel metal2 s 136638 0 136694 800 6 la_oenb[116]
port 520 nsew signal input
rlabel metal2 s 137558 0 137614 800 6 la_oenb[117]
port 521 nsew signal input
rlabel metal2 s 138478 0 138534 800 6 la_oenb[118]
port 522 nsew signal input
rlabel metal2 s 139398 0 139454 800 6 la_oenb[119]
port 523 nsew signal input
rlabel metal2 s 42338 0 42394 800 6 la_oenb[11]
port 524 nsew signal input
rlabel metal2 s 140226 0 140282 800 6 la_oenb[120]
port 525 nsew signal input
rlabel metal2 s 141146 0 141202 800 6 la_oenb[121]
port 526 nsew signal input
rlabel metal2 s 142066 0 142122 800 6 la_oenb[122]
port 527 nsew signal input
rlabel metal2 s 142986 0 143042 800 6 la_oenb[123]
port 528 nsew signal input
rlabel metal2 s 143906 0 143962 800 6 la_oenb[124]
port 529 nsew signal input
rlabel metal2 s 144734 0 144790 800 6 la_oenb[125]
port 530 nsew signal input
rlabel metal2 s 145654 0 145710 800 6 la_oenb[126]
port 531 nsew signal input
rlabel metal2 s 146574 0 146630 800 6 la_oenb[127]
port 532 nsew signal input
rlabel metal2 s 43166 0 43222 800 6 la_oenb[12]
port 533 nsew signal input
rlabel metal2 s 44086 0 44142 800 6 la_oenb[13]
port 534 nsew signal input
rlabel metal2 s 45006 0 45062 800 6 la_oenb[14]
port 535 nsew signal input
rlabel metal2 s 45926 0 45982 800 6 la_oenb[15]
port 536 nsew signal input
rlabel metal2 s 46754 0 46810 800 6 la_oenb[16]
port 537 nsew signal input
rlabel metal2 s 47674 0 47730 800 6 la_oenb[17]
port 538 nsew signal input
rlabel metal2 s 48594 0 48650 800 6 la_oenb[18]
port 539 nsew signal input
rlabel metal2 s 49514 0 49570 800 6 la_oenb[19]
port 540 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 la_oenb[1]
port 541 nsew signal input
rlabel metal2 s 50434 0 50490 800 6 la_oenb[20]
port 542 nsew signal input
rlabel metal2 s 51262 0 51318 800 6 la_oenb[21]
port 543 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 la_oenb[22]
port 544 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 la_oenb[23]
port 545 nsew signal input
rlabel metal2 s 54022 0 54078 800 6 la_oenb[24]
port 546 nsew signal input
rlabel metal2 s 54850 0 54906 800 6 la_oenb[25]
port 547 nsew signal input
rlabel metal2 s 55770 0 55826 800 6 la_oenb[26]
port 548 nsew signal input
rlabel metal2 s 56690 0 56746 800 6 la_oenb[27]
port 549 nsew signal input
rlabel metal2 s 57610 0 57666 800 6 la_oenb[28]
port 550 nsew signal input
rlabel metal2 s 58438 0 58494 800 6 la_oenb[29]
port 551 nsew signal input
rlabel metal2 s 34242 0 34298 800 6 la_oenb[2]
port 552 nsew signal input
rlabel metal2 s 59358 0 59414 800 6 la_oenb[30]
port 553 nsew signal input
rlabel metal2 s 60278 0 60334 800 6 la_oenb[31]
port 554 nsew signal input
rlabel metal2 s 61198 0 61254 800 6 la_oenb[32]
port 555 nsew signal input
rlabel metal2 s 62118 0 62174 800 6 la_oenb[33]
port 556 nsew signal input
rlabel metal2 s 62946 0 63002 800 6 la_oenb[34]
port 557 nsew signal input
rlabel metal2 s 63866 0 63922 800 6 la_oenb[35]
port 558 nsew signal input
rlabel metal2 s 64786 0 64842 800 6 la_oenb[36]
port 559 nsew signal input
rlabel metal2 s 65706 0 65762 800 6 la_oenb[37]
port 560 nsew signal input
rlabel metal2 s 66534 0 66590 800 6 la_oenb[38]
port 561 nsew signal input
rlabel metal2 s 67454 0 67510 800 6 la_oenb[39]
port 562 nsew signal input
rlabel metal2 s 35070 0 35126 800 6 la_oenb[3]
port 563 nsew signal input
rlabel metal2 s 68374 0 68430 800 6 la_oenb[40]
port 564 nsew signal input
rlabel metal2 s 69294 0 69350 800 6 la_oenb[41]
port 565 nsew signal input
rlabel metal2 s 70122 0 70178 800 6 la_oenb[42]
port 566 nsew signal input
rlabel metal2 s 71042 0 71098 800 6 la_oenb[43]
port 567 nsew signal input
rlabel metal2 s 71962 0 72018 800 6 la_oenb[44]
port 568 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 la_oenb[45]
port 569 nsew signal input
rlabel metal2 s 73802 0 73858 800 6 la_oenb[46]
port 570 nsew signal input
rlabel metal2 s 74630 0 74686 800 6 la_oenb[47]
port 571 nsew signal input
rlabel metal2 s 75550 0 75606 800 6 la_oenb[48]
port 572 nsew signal input
rlabel metal2 s 76470 0 76526 800 6 la_oenb[49]
port 573 nsew signal input
rlabel metal2 s 35990 0 36046 800 6 la_oenb[4]
port 574 nsew signal input
rlabel metal2 s 77390 0 77446 800 6 la_oenb[50]
port 575 nsew signal input
rlabel metal2 s 78218 0 78274 800 6 la_oenb[51]
port 576 nsew signal input
rlabel metal2 s 79138 0 79194 800 6 la_oenb[52]
port 577 nsew signal input
rlabel metal2 s 80058 0 80114 800 6 la_oenb[53]
port 578 nsew signal input
rlabel metal2 s 80978 0 81034 800 6 la_oenb[54]
port 579 nsew signal input
rlabel metal2 s 81806 0 81862 800 6 la_oenb[55]
port 580 nsew signal input
rlabel metal2 s 82726 0 82782 800 6 la_oenb[56]
port 581 nsew signal input
rlabel metal2 s 83646 0 83702 800 6 la_oenb[57]
port 582 nsew signal input
rlabel metal2 s 84566 0 84622 800 6 la_oenb[58]
port 583 nsew signal input
rlabel metal2 s 85486 0 85542 800 6 la_oenb[59]
port 584 nsew signal input
rlabel metal2 s 36910 0 36966 800 6 la_oenb[5]
port 585 nsew signal input
rlabel metal2 s 86314 0 86370 800 6 la_oenb[60]
port 586 nsew signal input
rlabel metal2 s 87234 0 87290 800 6 la_oenb[61]
port 587 nsew signal input
rlabel metal2 s 88154 0 88210 800 6 la_oenb[62]
port 588 nsew signal input
rlabel metal2 s 89074 0 89130 800 6 la_oenb[63]
port 589 nsew signal input
rlabel metal2 s 89902 0 89958 800 6 la_oenb[64]
port 590 nsew signal input
rlabel metal2 s 90822 0 90878 800 6 la_oenb[65]
port 591 nsew signal input
rlabel metal2 s 91742 0 91798 800 6 la_oenb[66]
port 592 nsew signal input
rlabel metal2 s 92662 0 92718 800 6 la_oenb[67]
port 593 nsew signal input
rlabel metal2 s 93490 0 93546 800 6 la_oenb[68]
port 594 nsew signal input
rlabel metal2 s 94410 0 94466 800 6 la_oenb[69]
port 595 nsew signal input
rlabel metal2 s 37830 0 37886 800 6 la_oenb[6]
port 596 nsew signal input
rlabel metal2 s 95330 0 95386 800 6 la_oenb[70]
port 597 nsew signal input
rlabel metal2 s 96250 0 96306 800 6 la_oenb[71]
port 598 nsew signal input
rlabel metal2 s 97170 0 97226 800 6 la_oenb[72]
port 599 nsew signal input
rlabel metal2 s 97998 0 98054 800 6 la_oenb[73]
port 600 nsew signal input
rlabel metal2 s 98918 0 98974 800 6 la_oenb[74]
port 601 nsew signal input
rlabel metal2 s 99838 0 99894 800 6 la_oenb[75]
port 602 nsew signal input
rlabel metal2 s 100758 0 100814 800 6 la_oenb[76]
port 603 nsew signal input
rlabel metal2 s 101586 0 101642 800 6 la_oenb[77]
port 604 nsew signal input
rlabel metal2 s 102506 0 102562 800 6 la_oenb[78]
port 605 nsew signal input
rlabel metal2 s 103426 0 103482 800 6 la_oenb[79]
port 606 nsew signal input
rlabel metal2 s 38750 0 38806 800 6 la_oenb[7]
port 607 nsew signal input
rlabel metal2 s 104346 0 104402 800 6 la_oenb[80]
port 608 nsew signal input
rlabel metal2 s 105174 0 105230 800 6 la_oenb[81]
port 609 nsew signal input
rlabel metal2 s 106094 0 106150 800 6 la_oenb[82]
port 610 nsew signal input
rlabel metal2 s 107014 0 107070 800 6 la_oenb[83]
port 611 nsew signal input
rlabel metal2 s 107934 0 107990 800 6 la_oenb[84]
port 612 nsew signal input
rlabel metal2 s 108854 0 108910 800 6 la_oenb[85]
port 613 nsew signal input
rlabel metal2 s 109682 0 109738 800 6 la_oenb[86]
port 614 nsew signal input
rlabel metal2 s 110602 0 110658 800 6 la_oenb[87]
port 615 nsew signal input
rlabel metal2 s 111522 0 111578 800 6 la_oenb[88]
port 616 nsew signal input
rlabel metal2 s 112442 0 112498 800 6 la_oenb[89]
port 617 nsew signal input
rlabel metal2 s 39578 0 39634 800 6 la_oenb[8]
port 618 nsew signal input
rlabel metal2 s 113270 0 113326 800 6 la_oenb[90]
port 619 nsew signal input
rlabel metal2 s 114190 0 114246 800 6 la_oenb[91]
port 620 nsew signal input
rlabel metal2 s 115110 0 115166 800 6 la_oenb[92]
port 621 nsew signal input
rlabel metal2 s 116030 0 116086 800 6 la_oenb[93]
port 622 nsew signal input
rlabel metal2 s 116858 0 116914 800 6 la_oenb[94]
port 623 nsew signal input
rlabel metal2 s 117778 0 117834 800 6 la_oenb[95]
port 624 nsew signal input
rlabel metal2 s 118698 0 118754 800 6 la_oenb[96]
port 625 nsew signal input
rlabel metal2 s 119618 0 119674 800 6 la_oenb[97]
port 626 nsew signal input
rlabel metal2 s 120538 0 120594 800 6 la_oenb[98]
port 627 nsew signal input
rlabel metal2 s 121366 0 121422 800 6 la_oenb[99]
port 628 nsew signal input
rlabel metal2 s 40498 0 40554 800 6 la_oenb[9]
port 629 nsew signal input
rlabel metal2 s 107842 166124 107898 166924 6 o_addr1[0]
port 630 nsew signal output
rlabel metal2 s 111522 166124 111578 166924 6 o_addr1[1]
port 631 nsew signal output
rlabel metal2 s 150438 0 150494 800 6 o_addr1[2]
port 632 nsew signal output
rlabel metal3 s 0 29792 800 29912 6 o_addr1[3]
port 633 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 o_addr1[4]
port 634 nsew signal output
rlabel metal2 s 153474 0 153530 800 6 o_addr1[5]
port 635 nsew signal output
rlabel metal2 s 154026 0 154082 800 6 o_addr1[6]
port 636 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 o_addr1[7]
port 637 nsew signal output
rlabel metal2 s 156786 0 156842 800 6 o_addr1[8]
port 638 nsew signal output
rlabel metal3 s 0 4632 800 4752 6 o_addr1_1[0]
port 639 nsew signal output
rlabel metal3 s 163980 15920 164780 16040 6 o_addr1_1[1]
port 640 nsew signal output
rlabel metal2 s 150162 0 150218 800 6 o_addr1_1[2]
port 641 nsew signal output
rlabel metal3 s 163980 30608 164780 30728 6 o_addr1_1[3]
port 642 nsew signal output
rlabel metal2 s 152554 0 152610 800 6 o_addr1_1[4]
port 643 nsew signal output
rlabel metal3 s 0 42304 800 42424 6 o_addr1_1[5]
port 644 nsew signal output
rlabel metal2 s 120814 166124 120870 166924 6 o_addr1_1[6]
port 645 nsew signal output
rlabel metal2 s 155590 0 155646 800 6 o_addr1_1[7]
port 646 nsew signal output
rlabel metal2 s 156418 0 156474 800 6 o_addr1_1[8]
port 647 nsew signal output
rlabel metal3 s 163980 1232 164780 1352 6 o_csb0
port 648 nsew signal output
rlabel metal2 s 147770 0 147826 800 6 o_csb0_1
port 649 nsew signal output
rlabel metal2 s 148046 0 148102 800 6 o_csb1
port 650 nsew signal output
rlabel metal3 s 163980 3680 164780 3800 6 o_csb1_1
port 651 nsew signal output
rlabel metal3 s 0 7760 800 7880 6 o_din0[0]
port 652 nsew signal output
rlabel metal2 s 157982 0 158038 800 6 o_din0[10]
port 653 nsew signal output
rlabel metal3 s 0 80112 800 80232 6 o_din0[11]
port 654 nsew signal output
rlabel metal3 s 163980 87048 164780 87168 6 o_din0[12]
port 655 nsew signal output
rlabel metal3 s 0 89632 800 89752 6 o_din0[13]
port 656 nsew signal output
rlabel metal3 s 163980 101736 164780 101856 6 o_din0[14]
port 657 nsew signal output
rlabel metal2 s 133694 166124 133750 166924 6 o_din0[15]
port 658 nsew signal output
rlabel metal3 s 0 102144 800 102264 6 o_din0[16]
port 659 nsew signal output
rlabel metal2 s 136546 166124 136602 166924 6 o_din0[17]
port 660 nsew signal output
rlabel metal2 s 160926 0 160982 800 6 o_din0[18]
port 661 nsew signal output
rlabel metal2 s 141146 166124 141202 166924 6 o_din0[19]
port 662 nsew signal output
rlabel metal3 s 163980 18368 164780 18488 6 o_din0[1]
port 663 nsew signal output
rlabel metal2 s 161570 0 161626 800 6 o_din0[20]
port 664 nsew signal output
rlabel metal2 s 142986 166124 143042 166924 6 o_din0[21]
port 665 nsew signal output
rlabel metal2 s 146666 166124 146722 166924 6 o_din0[22]
port 666 nsew signal output
rlabel metal3 s 0 127440 800 127560 6 o_din0[23]
port 667 nsew signal output
rlabel metal3 s 163980 143488 164780 143608 6 o_din0[24]
port 668 nsew signal output
rlabel metal2 s 162398 0 162454 800 6 o_din0[25]
port 669 nsew signal output
rlabel metal2 s 163042 0 163098 800 6 o_din0[26]
port 670 nsew signal output
rlabel metal3 s 0 149472 800 149592 6 o_din0[27]
port 671 nsew signal output
rlabel metal3 s 163980 158176 164780 158296 6 o_din0[28]
port 672 nsew signal output
rlabel metal3 s 163980 160624 164780 160744 6 o_din0[29]
port 673 nsew signal output
rlabel metal2 s 150714 0 150770 800 6 o_din0[2]
port 674 nsew signal output
rlabel metal3 s 163980 163072 164780 163192 6 o_din0[30]
port 675 nsew signal output
rlabel metal3 s 163980 165520 164780 165640 6 o_din0[31]
port 676 nsew signal output
rlabel metal3 s 163980 33056 164780 33176 6 o_din0[3]
port 677 nsew signal output
rlabel metal2 s 116122 166124 116178 166924 6 o_din0[4]
port 678 nsew signal output
rlabel metal2 s 118882 166124 118938 166924 6 o_din0[5]
port 679 nsew signal output
rlabel metal2 s 154394 0 154450 800 6 o_din0[6]
port 680 nsew signal output
rlabel metal2 s 155866 0 155922 800 6 o_din0[7]
port 681 nsew signal output
rlabel metal3 s 163980 74808 164780 74928 6 o_din0[8]
port 682 nsew signal output
rlabel metal2 s 157614 0 157670 800 6 o_din0[9]
port 683 nsew signal output
rlabel metal3 s 0 10888 800 11008 6 o_din0_1[0]
port 684 nsew signal output
rlabel metal2 s 127254 166124 127310 166924 6 o_din0_1[10]
port 685 nsew signal output
rlabel metal2 s 158534 0 158590 800 6 o_din0_1[11]
port 686 nsew signal output
rlabel metal2 s 159178 0 159234 800 6 o_din0_1[12]
port 687 nsew signal output
rlabel metal3 s 163980 96840 164780 96960 6 o_din0_1[13]
port 688 nsew signal output
rlabel metal2 s 131854 166124 131910 166924 6 o_din0_1[14]
port 689 nsew signal output
rlabel metal3 s 0 95888 800 96008 6 o_din0_1[15]
port 690 nsew signal output
rlabel metal2 s 160650 0 160706 800 6 o_din0_1[16]
port 691 nsew signal output
rlabel metal2 s 135626 166124 135682 166924 6 o_din0_1[17]
port 692 nsew signal output
rlabel metal2 s 140226 166124 140282 166924 6 o_din0_1[18]
port 693 nsew signal output
rlabel metal3 s 0 111664 800 111784 6 o_din0_1[19]
port 694 nsew signal output
rlabel metal2 s 149518 0 149574 800 6 o_din0_1[1]
port 695 nsew signal output
rlabel metal2 s 161202 0 161258 800 6 o_din0_1[20]
port 696 nsew signal output
rlabel metal3 s 163980 131248 164780 131368 6 o_din0_1[21]
port 697 nsew signal output
rlabel metal2 s 145746 166124 145802 166924 6 o_din0_1[22]
port 698 nsew signal output
rlabel metal2 s 149426 166124 149482 166924 6 o_din0_1[23]
port 699 nsew signal output
rlabel metal3 s 163980 141040 164780 141160 6 o_din0_1[24]
port 700 nsew signal output
rlabel metal3 s 163980 148384 164780 148504 6 o_din0_1[25]
port 701 nsew signal output
rlabel metal3 s 0 143080 800 143200 6 o_din0_1[26]
port 702 nsew signal output
rlabel metal2 s 163594 0 163650 800 6 o_din0_1[27]
port 703 nsew signal output
rlabel metal2 s 155958 166124 156014 166924 6 o_din0_1[28]
port 704 nsew signal output
rlabel metal2 s 164514 0 164570 800 6 o_din0_1[29]
port 705 nsew signal output
rlabel metal3 s 163980 23264 164780 23384 6 o_din0_1[2]
port 706 nsew signal output
rlabel metal2 s 161478 166124 161534 166924 6 o_din0_1[30]
port 707 nsew signal output
rlabel metal3 s 0 165112 800 165232 6 o_din0_1[31]
port 708 nsew signal output
rlabel metal2 s 152278 0 152334 800 6 o_din0_1[3]
port 709 nsew signal output
rlabel metal3 s 163980 50192 164780 50312 6 o_din0_1[4]
port 710 nsew signal output
rlabel metal2 s 117962 166124 118018 166924 6 o_din0_1[5]
port 711 nsew signal output
rlabel metal2 s 121734 166124 121790 166924 6 o_din0_1[6]
port 712 nsew signal output
rlabel metal3 s 163980 65016 164780 65136 6 o_din0_1[7]
port 713 nsew signal output
rlabel metal3 s 163980 72360 164780 72480 6 o_din0_1[8]
port 714 nsew signal output
rlabel metal2 s 124494 166124 124550 166924 6 o_din0_1[9]
port 715 nsew signal output
rlabel metal2 s 108762 166124 108818 166924 6 o_waddr0[0]
port 716 nsew signal output
rlabel metal3 s 0 14016 800 14136 6 o_waddr0[1]
port 717 nsew signal output
rlabel metal2 s 151082 0 151138 800 6 o_waddr0[2]
port 718 nsew signal output
rlabel metal3 s 163980 37952 164780 38072 6 o_waddr0[3]
port 719 nsew signal output
rlabel metal2 s 152830 0 152886 800 6 o_waddr0[4]
port 720 nsew signal output
rlabel metal3 s 0 45568 800 45688 6 o_waddr0[5]
port 721 nsew signal output
rlabel metal3 s 163980 62568 164780 62688 6 o_waddr0[6]
port 722 nsew signal output
rlabel metal3 s 163980 69912 164780 70032 6 o_waddr0[7]
port 723 nsew signal output
rlabel metal2 s 157062 0 157118 800 6 o_waddr0[8]
port 724 nsew signal output
rlabel metal2 s 148966 0 149022 800 6 o_waddr0_1[0]
port 725 nsew signal output
rlabel metal2 s 112442 166124 112498 166924 6 o_waddr0_1[1]
port 726 nsew signal output
rlabel metal3 s 163980 25712 164780 25832 6 o_waddr0_1[2]
port 727 nsew signal output
rlabel metal3 s 163980 35504 164780 35624 6 o_waddr0_1[3]
port 728 nsew signal output
rlabel metal2 s 117042 166124 117098 166924 6 o_waddr0_1[4]
port 729 nsew signal output
rlabel metal3 s 163980 57672 164780 57792 6 o_waddr0_1[5]
port 730 nsew signal output
rlabel metal2 s 154670 0 154726 800 6 o_waddr0_1[6]
port 731 nsew signal output
rlabel metal3 s 163980 67464 164780 67584 6 o_waddr0_1[7]
port 732 nsew signal output
rlabel metal3 s 163980 77256 164780 77376 6 o_waddr0_1[8]
port 733 nsew signal output
rlabel metal2 s 106002 166124 106058 166924 6 o_web0
port 734 nsew signal output
rlabel metal3 s 163980 6128 164780 6248 6 o_web0_1
port 735 nsew signal output
rlabel metal2 s 109682 166124 109738 166924 6 o_wmask0[0]
port 736 nsew signal output
rlabel metal2 s 149886 0 149942 800 6 o_wmask0[1]
port 737 nsew signal output
rlabel metal3 s 0 26664 800 26784 6 o_wmask0[2]
port 738 nsew signal output
rlabel metal2 s 115202 166124 115258 166924 6 o_wmask0[3]
port 739 nsew signal output
rlabel metal2 s 149242 0 149298 800 6 o_wmask0_1[0]
port 740 nsew signal output
rlabel metal3 s 0 17144 800 17264 6 o_wmask0_1[1]
port 741 nsew signal output
rlabel metal2 s 151358 0 151414 800 6 o_wmask0_1[2]
port 742 nsew signal output
rlabel metal3 s 163980 40400 164780 40520 6 o_wmask0_1[3]
port 743 nsew signal output
rlabel metal4 s 4208 2128 4528 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 34928 2128 35248 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 65648 2128 65968 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 96368 2128 96688 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 127088 2128 127408 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 157808 2128 158128 164336 6 vccd1
port 744 nsew power input
rlabel metal4 s 19568 2128 19888 164336 6 vssd1
port 745 nsew ground input
rlabel metal4 s 50288 2128 50608 164336 6 vssd1
port 745 nsew ground input
rlabel metal4 s 81008 2128 81328 164336 6 vssd1
port 745 nsew ground input
rlabel metal4 s 111728 2128 112048 164336 6 vssd1
port 745 nsew ground input
rlabel metal4 s 142448 2128 142768 164336 6 vssd1
port 745 nsew ground input
rlabel metal2 s 110 0 166 800 6 wb_clk_i
port 746 nsew signal input
rlabel metal2 s 386 0 442 800 6 wb_rst_i
port 747 nsew signal input
rlabel metal2 s 662 0 718 800 6 wbs_ack_o
port 748 nsew signal output
rlabel metal2 s 1858 0 1914 800 6 wbs_adr_i[0]
port 749 nsew signal input
rlabel metal2 s 12070 0 12126 800 6 wbs_adr_i[10]
port 750 nsew signal input
rlabel metal2 s 12990 0 13046 800 6 wbs_adr_i[11]
port 751 nsew signal input
rlabel metal2 s 13818 0 13874 800 6 wbs_adr_i[12]
port 752 nsew signal input
rlabel metal2 s 14738 0 14794 800 6 wbs_adr_i[13]
port 753 nsew signal input
rlabel metal2 s 15658 0 15714 800 6 wbs_adr_i[14]
port 754 nsew signal input
rlabel metal2 s 16578 0 16634 800 6 wbs_adr_i[15]
port 755 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[16]
port 756 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_adr_i[17]
port 757 nsew signal input
rlabel metal2 s 19246 0 19302 800 6 wbs_adr_i[18]
port 758 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_adr_i[19]
port 759 nsew signal input
rlabel metal2 s 3054 0 3110 800 6 wbs_adr_i[1]
port 760 nsew signal input
rlabel metal2 s 20994 0 21050 800 6 wbs_adr_i[20]
port 761 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 wbs_adr_i[21]
port 762 nsew signal input
rlabel metal2 s 22834 0 22890 800 6 wbs_adr_i[22]
port 763 nsew signal input
rlabel metal2 s 23754 0 23810 800 6 wbs_adr_i[23]
port 764 nsew signal input
rlabel metal2 s 24674 0 24730 800 6 wbs_adr_i[24]
port 765 nsew signal input
rlabel metal2 s 25502 0 25558 800 6 wbs_adr_i[25]
port 766 nsew signal input
rlabel metal2 s 26422 0 26478 800 6 wbs_adr_i[26]
port 767 nsew signal input
rlabel metal2 s 27342 0 27398 800 6 wbs_adr_i[27]
port 768 nsew signal input
rlabel metal2 s 28262 0 28318 800 6 wbs_adr_i[28]
port 769 nsew signal input
rlabel metal2 s 29090 0 29146 800 6 wbs_adr_i[29]
port 770 nsew signal input
rlabel metal2 s 4250 0 4306 800 6 wbs_adr_i[2]
port 771 nsew signal input
rlabel metal2 s 30010 0 30066 800 6 wbs_adr_i[30]
port 772 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 wbs_adr_i[31]
port 773 nsew signal input
rlabel metal2 s 5446 0 5502 800 6 wbs_adr_i[3]
port 774 nsew signal input
rlabel metal2 s 6642 0 6698 800 6 wbs_adr_i[4]
port 775 nsew signal input
rlabel metal2 s 7562 0 7618 800 6 wbs_adr_i[5]
port 776 nsew signal input
rlabel metal2 s 8482 0 8538 800 6 wbs_adr_i[6]
port 777 nsew signal input
rlabel metal2 s 9310 0 9366 800 6 wbs_adr_i[7]
port 778 nsew signal input
rlabel metal2 s 10230 0 10286 800 6 wbs_adr_i[8]
port 779 nsew signal input
rlabel metal2 s 11150 0 11206 800 6 wbs_adr_i[9]
port 780 nsew signal input
rlabel metal2 s 938 0 994 800 6 wbs_cyc_i
port 781 nsew signal input
rlabel metal2 s 2134 0 2190 800 6 wbs_dat_i[0]
port 782 nsew signal input
rlabel metal2 s 12346 0 12402 800 6 wbs_dat_i[10]
port 783 nsew signal input
rlabel metal2 s 13266 0 13322 800 6 wbs_dat_i[11]
port 784 nsew signal input
rlabel metal2 s 14186 0 14242 800 6 wbs_dat_i[12]
port 785 nsew signal input
rlabel metal2 s 15014 0 15070 800 6 wbs_dat_i[13]
port 786 nsew signal input
rlabel metal2 s 15934 0 15990 800 6 wbs_dat_i[14]
port 787 nsew signal input
rlabel metal2 s 16854 0 16910 800 6 wbs_dat_i[15]
port 788 nsew signal input
rlabel metal2 s 17774 0 17830 800 6 wbs_dat_i[16]
port 789 nsew signal input
rlabel metal2 s 18602 0 18658 800 6 wbs_dat_i[17]
port 790 nsew signal input
rlabel metal2 s 19522 0 19578 800 6 wbs_dat_i[18]
port 791 nsew signal input
rlabel metal2 s 20442 0 20498 800 6 wbs_dat_i[19]
port 792 nsew signal input
rlabel metal2 s 3330 0 3386 800 6 wbs_dat_i[1]
port 793 nsew signal input
rlabel metal2 s 21362 0 21418 800 6 wbs_dat_i[20]
port 794 nsew signal input
rlabel metal2 s 22190 0 22246 800 6 wbs_dat_i[21]
port 795 nsew signal input
rlabel metal2 s 23110 0 23166 800 6 wbs_dat_i[22]
port 796 nsew signal input
rlabel metal2 s 24030 0 24086 800 6 wbs_dat_i[23]
port 797 nsew signal input
rlabel metal2 s 24950 0 25006 800 6 wbs_dat_i[24]
port 798 nsew signal input
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_i[25]
port 799 nsew signal input
rlabel metal2 s 26698 0 26754 800 6 wbs_dat_i[26]
port 800 nsew signal input
rlabel metal2 s 27618 0 27674 800 6 wbs_dat_i[27]
port 801 nsew signal input
rlabel metal2 s 28538 0 28594 800 6 wbs_dat_i[28]
port 802 nsew signal input
rlabel metal2 s 29458 0 29514 800 6 wbs_dat_i[29]
port 803 nsew signal input
rlabel metal2 s 4526 0 4582 800 6 wbs_dat_i[2]
port 804 nsew signal input
rlabel metal2 s 30286 0 30342 800 6 wbs_dat_i[30]
port 805 nsew signal input
rlabel metal2 s 31206 0 31262 800 6 wbs_dat_i[31]
port 806 nsew signal input
rlabel metal2 s 5722 0 5778 800 6 wbs_dat_i[3]
port 807 nsew signal input
rlabel metal2 s 6918 0 6974 800 6 wbs_dat_i[4]
port 808 nsew signal input
rlabel metal2 s 7838 0 7894 800 6 wbs_dat_i[5]
port 809 nsew signal input
rlabel metal2 s 8758 0 8814 800 6 wbs_dat_i[6]
port 810 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 wbs_dat_i[7]
port 811 nsew signal input
rlabel metal2 s 10506 0 10562 800 6 wbs_dat_i[8]
port 812 nsew signal input
rlabel metal2 s 11426 0 11482 800 6 wbs_dat_i[9]
port 813 nsew signal input
rlabel metal2 s 2502 0 2558 800 6 wbs_dat_o[0]
port 814 nsew signal output
rlabel metal2 s 12622 0 12678 800 6 wbs_dat_o[10]
port 815 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 wbs_dat_o[11]
port 816 nsew signal output
rlabel metal2 s 14462 0 14518 800 6 wbs_dat_o[12]
port 817 nsew signal output
rlabel metal2 s 15382 0 15438 800 6 wbs_dat_o[13]
port 818 nsew signal output
rlabel metal2 s 16210 0 16266 800 6 wbs_dat_o[14]
port 819 nsew signal output
rlabel metal2 s 17130 0 17186 800 6 wbs_dat_o[15]
port 820 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 wbs_dat_o[16]
port 821 nsew signal output
rlabel metal2 s 18970 0 19026 800 6 wbs_dat_o[17]
port 822 nsew signal output
rlabel metal2 s 19798 0 19854 800 6 wbs_dat_o[18]
port 823 nsew signal output
rlabel metal2 s 20718 0 20774 800 6 wbs_dat_o[19]
port 824 nsew signal output
rlabel metal2 s 3698 0 3754 800 6 wbs_dat_o[1]
port 825 nsew signal output
rlabel metal2 s 21638 0 21694 800 6 wbs_dat_o[20]
port 826 nsew signal output
rlabel metal2 s 22558 0 22614 800 6 wbs_dat_o[21]
port 827 nsew signal output
rlabel metal2 s 23386 0 23442 800 6 wbs_dat_o[22]
port 828 nsew signal output
rlabel metal2 s 24306 0 24362 800 6 wbs_dat_o[23]
port 829 nsew signal output
rlabel metal2 s 25226 0 25282 800 6 wbs_dat_o[24]
port 830 nsew signal output
rlabel metal2 s 26146 0 26202 800 6 wbs_dat_o[25]
port 831 nsew signal output
rlabel metal2 s 27066 0 27122 800 6 wbs_dat_o[26]
port 832 nsew signal output
rlabel metal2 s 27894 0 27950 800 6 wbs_dat_o[27]
port 833 nsew signal output
rlabel metal2 s 28814 0 28870 800 6 wbs_dat_o[28]
port 834 nsew signal output
rlabel metal2 s 29734 0 29790 800 6 wbs_dat_o[29]
port 835 nsew signal output
rlabel metal2 s 4894 0 4950 800 6 wbs_dat_o[2]
port 836 nsew signal output
rlabel metal2 s 30654 0 30710 800 6 wbs_dat_o[30]
port 837 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_o[31]
port 838 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 wbs_dat_o[3]
port 839 nsew signal output
rlabel metal2 s 7286 0 7342 800 6 wbs_dat_o[4]
port 840 nsew signal output
rlabel metal2 s 8114 0 8170 800 6 wbs_dat_o[5]
port 841 nsew signal output
rlabel metal2 s 9034 0 9090 800 6 wbs_dat_o[6]
port 842 nsew signal output
rlabel metal2 s 9954 0 10010 800 6 wbs_dat_o[7]
port 843 nsew signal output
rlabel metal2 s 10874 0 10930 800 6 wbs_dat_o[8]
port 844 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[9]
port 845 nsew signal output
rlabel metal2 s 2778 0 2834 800 6 wbs_sel_i[0]
port 846 nsew signal input
rlabel metal2 s 3974 0 4030 800 6 wbs_sel_i[1]
port 847 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_sel_i[2]
port 848 nsew signal input
rlabel metal2 s 6366 0 6422 800 6 wbs_sel_i[3]
port 849 nsew signal input
rlabel metal2 s 1306 0 1362 800 6 wbs_stb_i
port 850 nsew signal input
rlabel metal2 s 1582 0 1638 800 6 wbs_we_i
port 851 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 164780 166924
string LEFview TRUE
string GDS_FILE /local/caravel_user_project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 82295346
string GDS_START 1378666
<< end >>

