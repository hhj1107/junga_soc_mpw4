magic
tech sky130A
magscale 1 2
timestamp 1640663083
<< obsli1 >>
rect 1409 2261 163731 164203
<< obsm1 >>
rect 290 8 163743 164336
<< metal2 >>
rect 478 165957 534 166757
rect 1398 165957 1454 166757
rect 2410 165957 2466 166757
rect 3330 165957 3386 166757
rect 4342 165957 4398 166757
rect 5262 165957 5318 166757
rect 6274 165957 6330 166757
rect 7286 165957 7342 166757
rect 8206 165957 8262 166757
rect 9218 165957 9274 166757
rect 10138 165957 10194 166757
rect 11150 165957 11206 166757
rect 12162 165957 12218 166757
rect 13082 165957 13138 166757
rect 14094 165957 14150 166757
rect 15014 165957 15070 166757
rect 16026 165957 16082 166757
rect 16946 165957 17002 166757
rect 17958 165957 18014 166757
rect 18970 165957 19026 166757
rect 19890 165957 19946 166757
rect 20902 165957 20958 166757
rect 21822 165957 21878 166757
rect 22834 165957 22890 166757
rect 23846 165957 23902 166757
rect 24766 165957 24822 166757
rect 25778 165957 25834 166757
rect 26698 165957 26754 166757
rect 27710 165957 27766 166757
rect 28630 165957 28686 166757
rect 29642 165957 29698 166757
rect 30654 165957 30710 166757
rect 31574 165957 31630 166757
rect 32586 165957 32642 166757
rect 33506 165957 33562 166757
rect 34518 165957 34574 166757
rect 35530 165957 35586 166757
rect 36450 165957 36506 166757
rect 37462 165957 37518 166757
rect 38382 165957 38438 166757
rect 39394 165957 39450 166757
rect 40406 165957 40462 166757
rect 41326 165957 41382 166757
rect 42338 165957 42394 166757
rect 43258 165957 43314 166757
rect 44270 165957 44326 166757
rect 45190 165957 45246 166757
rect 46202 165957 46258 166757
rect 47214 165957 47270 166757
rect 48134 165957 48190 166757
rect 49146 165957 49202 166757
rect 50066 165957 50122 166757
rect 51078 165957 51134 166757
rect 52090 165957 52146 166757
rect 53010 165957 53066 166757
rect 54022 165957 54078 166757
rect 54942 165957 54998 166757
rect 55954 165957 56010 166757
rect 56874 165957 56930 166757
rect 57886 165957 57942 166757
rect 58898 165957 58954 166757
rect 59818 165957 59874 166757
rect 60830 165957 60886 166757
rect 61750 165957 61806 166757
rect 62762 165957 62818 166757
rect 63774 165957 63830 166757
rect 64694 165957 64750 166757
rect 65706 165957 65762 166757
rect 66626 165957 66682 166757
rect 67638 165957 67694 166757
rect 68650 165957 68706 166757
rect 69570 165957 69626 166757
rect 70582 165957 70638 166757
rect 71502 165957 71558 166757
rect 72514 165957 72570 166757
rect 73434 165957 73490 166757
rect 74446 165957 74502 166757
rect 75458 165957 75514 166757
rect 76378 165957 76434 166757
rect 77390 165957 77446 166757
rect 78310 165957 78366 166757
rect 79322 165957 79378 166757
rect 80334 165957 80390 166757
rect 81254 165957 81310 166757
rect 82266 165957 82322 166757
rect 83186 165957 83242 166757
rect 84198 165957 84254 166757
rect 85118 165957 85174 166757
rect 86130 165957 86186 166757
rect 87142 165957 87198 166757
rect 88062 165957 88118 166757
rect 89074 165957 89130 166757
rect 89994 165957 90050 166757
rect 91006 165957 91062 166757
rect 92018 165957 92074 166757
rect 92938 165957 92994 166757
rect 93950 165957 94006 166757
rect 94870 165957 94926 166757
rect 95882 165957 95938 166757
rect 96802 165957 96858 166757
rect 97814 165957 97870 166757
rect 98826 165957 98882 166757
rect 99746 165957 99802 166757
rect 100758 165957 100814 166757
rect 101678 165957 101734 166757
rect 102690 165957 102746 166757
rect 103702 165957 103758 166757
rect 104622 165957 104678 166757
rect 105634 165957 105690 166757
rect 106554 165957 106610 166757
rect 107566 165957 107622 166757
rect 108578 165957 108634 166757
rect 109498 165957 109554 166757
rect 110510 165957 110566 166757
rect 111430 165957 111486 166757
rect 112442 165957 112498 166757
rect 113362 165957 113418 166757
rect 114374 165957 114430 166757
rect 115386 165957 115442 166757
rect 116306 165957 116362 166757
rect 117318 165957 117374 166757
rect 118238 165957 118294 166757
rect 119250 165957 119306 166757
rect 120262 165957 120318 166757
rect 121182 165957 121238 166757
rect 122194 165957 122250 166757
rect 123114 165957 123170 166757
rect 124126 165957 124182 166757
rect 125046 165957 125102 166757
rect 126058 165957 126114 166757
rect 127070 165957 127126 166757
rect 127990 165957 128046 166757
rect 129002 165957 129058 166757
rect 129922 165957 129978 166757
rect 130934 165957 130990 166757
rect 131946 165957 132002 166757
rect 132866 165957 132922 166757
rect 133878 165957 133934 166757
rect 134798 165957 134854 166757
rect 135810 165957 135866 166757
rect 136822 165957 136878 166757
rect 137742 165957 137798 166757
rect 138754 165957 138810 166757
rect 139674 165957 139730 166757
rect 140686 165957 140742 166757
rect 141606 165957 141662 166757
rect 142618 165957 142674 166757
rect 143630 165957 143686 166757
rect 144550 165957 144606 166757
rect 145562 165957 145618 166757
rect 146482 165957 146538 166757
rect 147494 165957 147550 166757
rect 148506 165957 148562 166757
rect 149426 165957 149482 166757
rect 150438 165957 150494 166757
rect 151358 165957 151414 166757
rect 152370 165957 152426 166757
rect 153290 165957 153346 166757
rect 154302 165957 154358 166757
rect 155314 165957 155370 166757
rect 156234 165957 156290 166757
rect 157246 165957 157302 166757
rect 158166 165957 158222 166757
rect 159178 165957 159234 166757
rect 160190 165957 160246 166757
rect 161110 165957 161166 166757
rect 162122 165957 162178 166757
rect 163042 165957 163098 166757
rect 164054 165957 164110 166757
rect 478 0 534 800
rect 1398 0 1454 800
rect 2318 0 2374 800
rect 3238 0 3294 800
rect 4158 0 4214 800
rect 5170 0 5226 800
rect 6090 0 6146 800
rect 7010 0 7066 800
rect 7930 0 7986 800
rect 8942 0 8998 800
rect 9862 0 9918 800
rect 10782 0 10838 800
rect 11702 0 11758 800
rect 12622 0 12678 800
rect 13634 0 13690 800
rect 14554 0 14610 800
rect 15474 0 15530 800
rect 16394 0 16450 800
rect 17406 0 17462 800
rect 18326 0 18382 800
rect 19246 0 19302 800
rect 20166 0 20222 800
rect 21086 0 21142 800
rect 22098 0 22154 800
rect 23018 0 23074 800
rect 23938 0 23994 800
rect 24858 0 24914 800
rect 25870 0 25926 800
rect 26790 0 26846 800
rect 27710 0 27766 800
rect 28630 0 28686 800
rect 29550 0 29606 800
rect 30562 0 30618 800
rect 31482 0 31538 800
rect 32402 0 32458 800
rect 33322 0 33378 800
rect 34334 0 34390 800
rect 35254 0 35310 800
rect 36174 0 36230 800
rect 37094 0 37150 800
rect 38014 0 38070 800
rect 39026 0 39082 800
rect 39946 0 40002 800
rect 40866 0 40922 800
rect 41786 0 41842 800
rect 42798 0 42854 800
rect 43718 0 43774 800
rect 44638 0 44694 800
rect 45558 0 45614 800
rect 46478 0 46534 800
rect 47490 0 47546 800
rect 48410 0 48466 800
rect 49330 0 49386 800
rect 50250 0 50306 800
rect 51262 0 51318 800
rect 52182 0 52238 800
rect 53102 0 53158 800
rect 54022 0 54078 800
rect 54942 0 54998 800
rect 55954 0 56010 800
rect 56874 0 56930 800
rect 57794 0 57850 800
rect 58714 0 58770 800
rect 59726 0 59782 800
rect 60646 0 60702 800
rect 61566 0 61622 800
rect 62486 0 62542 800
rect 63406 0 63462 800
rect 64418 0 64474 800
rect 65338 0 65394 800
rect 66258 0 66314 800
rect 67178 0 67234 800
rect 68190 0 68246 800
rect 69110 0 69166 800
rect 70030 0 70086 800
rect 70950 0 71006 800
rect 71870 0 71926 800
rect 72882 0 72938 800
rect 73802 0 73858 800
rect 74722 0 74778 800
rect 75642 0 75698 800
rect 76654 0 76710 800
rect 77574 0 77630 800
rect 78494 0 78550 800
rect 79414 0 79470 800
rect 80334 0 80390 800
rect 81346 0 81402 800
rect 82266 0 82322 800
rect 83186 0 83242 800
rect 84106 0 84162 800
rect 85118 0 85174 800
rect 86038 0 86094 800
rect 86958 0 87014 800
rect 87878 0 87934 800
rect 88798 0 88854 800
rect 89810 0 89866 800
rect 90730 0 90786 800
rect 91650 0 91706 800
rect 92570 0 92626 800
rect 93582 0 93638 800
rect 94502 0 94558 800
rect 95422 0 95478 800
rect 96342 0 96398 800
rect 97262 0 97318 800
rect 98274 0 98330 800
rect 99194 0 99250 800
rect 100114 0 100170 800
rect 101034 0 101090 800
rect 102046 0 102102 800
rect 102966 0 103022 800
rect 103886 0 103942 800
rect 104806 0 104862 800
rect 105726 0 105782 800
rect 106738 0 106794 800
rect 107658 0 107714 800
rect 108578 0 108634 800
rect 109498 0 109554 800
rect 110510 0 110566 800
rect 111430 0 111486 800
rect 112350 0 112406 800
rect 113270 0 113326 800
rect 114190 0 114246 800
rect 115202 0 115258 800
rect 116122 0 116178 800
rect 117042 0 117098 800
rect 117962 0 118018 800
rect 118974 0 119030 800
rect 119894 0 119950 800
rect 120814 0 120870 800
rect 121734 0 121790 800
rect 122654 0 122710 800
rect 123666 0 123722 800
rect 124586 0 124642 800
rect 125506 0 125562 800
rect 126426 0 126482 800
rect 127438 0 127494 800
rect 128358 0 128414 800
rect 129278 0 129334 800
rect 130198 0 130254 800
rect 131118 0 131174 800
rect 132130 0 132186 800
rect 133050 0 133106 800
rect 133970 0 134026 800
rect 134890 0 134946 800
rect 135902 0 135958 800
rect 136822 0 136878 800
rect 137742 0 137798 800
rect 138662 0 138718 800
rect 139582 0 139638 800
rect 140594 0 140650 800
rect 141514 0 141570 800
rect 142434 0 142490 800
rect 143354 0 143410 800
rect 144366 0 144422 800
rect 145286 0 145342 800
rect 146206 0 146262 800
rect 147126 0 147182 800
rect 148046 0 148102 800
rect 149058 0 149114 800
rect 149978 0 150034 800
rect 150898 0 150954 800
rect 151818 0 151874 800
rect 152830 0 152886 800
rect 153750 0 153806 800
rect 154670 0 154726 800
rect 155590 0 155646 800
rect 156510 0 156566 800
rect 157522 0 157578 800
rect 158442 0 158498 800
rect 159362 0 159418 800
rect 160282 0 160338 800
rect 161294 0 161350 800
rect 162214 0 162270 800
rect 163134 0 163190 800
rect 164054 0 164110 800
<< obsm2 >>
rect 294 165901 422 166002
rect 590 165901 1342 166002
rect 1510 165901 2354 166002
rect 2522 165901 3274 166002
rect 3442 165901 4286 166002
rect 4454 165901 5206 166002
rect 5374 165901 6218 166002
rect 6386 165901 7230 166002
rect 7398 165901 8150 166002
rect 8318 165901 9162 166002
rect 9330 165901 10082 166002
rect 10250 165901 11094 166002
rect 11262 165901 12106 166002
rect 12274 165901 13026 166002
rect 13194 165901 14038 166002
rect 14206 165901 14958 166002
rect 15126 165901 15970 166002
rect 16138 165901 16890 166002
rect 17058 165901 17902 166002
rect 18070 165901 18914 166002
rect 19082 165901 19834 166002
rect 20002 165901 20846 166002
rect 21014 165901 21766 166002
rect 21934 165901 22778 166002
rect 22946 165901 23790 166002
rect 23958 165901 24710 166002
rect 24878 165901 25722 166002
rect 25890 165901 26642 166002
rect 26810 165901 27654 166002
rect 27822 165901 28574 166002
rect 28742 165901 29586 166002
rect 29754 165901 30598 166002
rect 30766 165901 31518 166002
rect 31686 165901 32530 166002
rect 32698 165901 33450 166002
rect 33618 165901 34462 166002
rect 34630 165901 35474 166002
rect 35642 165901 36394 166002
rect 36562 165901 37406 166002
rect 37574 165901 38326 166002
rect 38494 165901 39338 166002
rect 39506 165901 40350 166002
rect 40518 165901 41270 166002
rect 41438 165901 42282 166002
rect 42450 165901 43202 166002
rect 43370 165901 44214 166002
rect 44382 165901 45134 166002
rect 45302 165901 46146 166002
rect 46314 165901 47158 166002
rect 47326 165901 48078 166002
rect 48246 165901 49090 166002
rect 49258 165901 50010 166002
rect 50178 165901 51022 166002
rect 51190 165901 52034 166002
rect 52202 165901 52954 166002
rect 53122 165901 53966 166002
rect 54134 165901 54886 166002
rect 55054 165901 55898 166002
rect 56066 165901 56818 166002
rect 56986 165901 57830 166002
rect 57998 165901 58842 166002
rect 59010 165901 59762 166002
rect 59930 165901 60774 166002
rect 60942 165901 61694 166002
rect 61862 165901 62706 166002
rect 62874 165901 63718 166002
rect 63886 165901 64638 166002
rect 64806 165901 65650 166002
rect 65818 165901 66570 166002
rect 66738 165901 67582 166002
rect 67750 165901 68594 166002
rect 68762 165901 69514 166002
rect 69682 165901 70526 166002
rect 70694 165901 71446 166002
rect 71614 165901 72458 166002
rect 72626 165901 73378 166002
rect 73546 165901 74390 166002
rect 74558 165901 75402 166002
rect 75570 165901 76322 166002
rect 76490 165901 77334 166002
rect 77502 165901 78254 166002
rect 78422 165901 79266 166002
rect 79434 165901 80278 166002
rect 80446 165901 81198 166002
rect 81366 165901 82210 166002
rect 82378 165901 83130 166002
rect 83298 165901 84142 166002
rect 84310 165901 85062 166002
rect 85230 165901 86074 166002
rect 86242 165901 87086 166002
rect 87254 165901 88006 166002
rect 88174 165901 89018 166002
rect 89186 165901 89938 166002
rect 90106 165901 90950 166002
rect 91118 165901 91962 166002
rect 92130 165901 92882 166002
rect 93050 165901 93894 166002
rect 94062 165901 94814 166002
rect 94982 165901 95826 166002
rect 95994 165901 96746 166002
rect 96914 165901 97758 166002
rect 97926 165901 98770 166002
rect 98938 165901 99690 166002
rect 99858 165901 100702 166002
rect 100870 165901 101622 166002
rect 101790 165901 102634 166002
rect 102802 165901 103646 166002
rect 103814 165901 104566 166002
rect 104734 165901 105578 166002
rect 105746 165901 106498 166002
rect 106666 165901 107510 166002
rect 107678 165901 108522 166002
rect 108690 165901 109442 166002
rect 109610 165901 110454 166002
rect 110622 165901 111374 166002
rect 111542 165901 112386 166002
rect 112554 165901 113306 166002
rect 113474 165901 114318 166002
rect 114486 165901 115330 166002
rect 115498 165901 116250 166002
rect 116418 165901 117262 166002
rect 117430 165901 118182 166002
rect 118350 165901 119194 166002
rect 119362 165901 120206 166002
rect 120374 165901 121126 166002
rect 121294 165901 122138 166002
rect 122306 165901 123058 166002
rect 123226 165901 124070 166002
rect 124238 165901 124990 166002
rect 125158 165901 126002 166002
rect 126170 165901 127014 166002
rect 127182 165901 127934 166002
rect 128102 165901 128946 166002
rect 129114 165901 129866 166002
rect 130034 165901 130878 166002
rect 131046 165901 131890 166002
rect 132058 165901 132810 166002
rect 132978 165901 133822 166002
rect 133990 165901 134742 166002
rect 134910 165901 135754 166002
rect 135922 165901 136766 166002
rect 136934 165901 137686 166002
rect 137854 165901 138698 166002
rect 138866 165901 139618 166002
rect 139786 165901 140630 166002
rect 140798 165901 141550 166002
rect 141718 165901 142562 166002
rect 142730 165901 143574 166002
rect 143742 165901 144494 166002
rect 144662 165901 145506 166002
rect 145674 165901 146426 166002
rect 146594 165901 147438 166002
rect 147606 165901 148450 166002
rect 148618 165901 149370 166002
rect 149538 165901 150382 166002
rect 150550 165901 151302 166002
rect 151470 165901 152314 166002
rect 152482 165901 153234 166002
rect 153402 165901 154246 166002
rect 154414 165901 155258 166002
rect 155426 165901 156178 166002
rect 156346 165901 157190 166002
rect 157358 165901 158110 166002
rect 158278 165901 159122 166002
rect 159290 165901 160134 166002
rect 160302 165901 161054 166002
rect 161222 165901 162066 166002
rect 162234 165901 162986 166002
rect 294 856 163006 165901
rect 294 2 422 856
rect 590 2 1342 856
rect 1510 2 2262 856
rect 2430 2 3182 856
rect 3350 2 4102 856
rect 4270 2 5114 856
rect 5282 2 6034 856
rect 6202 2 6954 856
rect 7122 2 7874 856
rect 8042 2 8886 856
rect 9054 2 9806 856
rect 9974 2 10726 856
rect 10894 2 11646 856
rect 11814 2 12566 856
rect 12734 2 13578 856
rect 13746 2 14498 856
rect 14666 2 15418 856
rect 15586 2 16338 856
rect 16506 2 17350 856
rect 17518 2 18270 856
rect 18438 2 19190 856
rect 19358 2 20110 856
rect 20278 2 21030 856
rect 21198 2 22042 856
rect 22210 2 22962 856
rect 23130 2 23882 856
rect 24050 2 24802 856
rect 24970 2 25814 856
rect 25982 2 26734 856
rect 26902 2 27654 856
rect 27822 2 28574 856
rect 28742 2 29494 856
rect 29662 2 30506 856
rect 30674 2 31426 856
rect 31594 2 32346 856
rect 32514 2 33266 856
rect 33434 2 34278 856
rect 34446 2 35198 856
rect 35366 2 36118 856
rect 36286 2 37038 856
rect 37206 2 37958 856
rect 38126 2 38970 856
rect 39138 2 39890 856
rect 40058 2 40810 856
rect 40978 2 41730 856
rect 41898 2 42742 856
rect 42910 2 43662 856
rect 43830 2 44582 856
rect 44750 2 45502 856
rect 45670 2 46422 856
rect 46590 2 47434 856
rect 47602 2 48354 856
rect 48522 2 49274 856
rect 49442 2 50194 856
rect 50362 2 51206 856
rect 51374 2 52126 856
rect 52294 2 53046 856
rect 53214 2 53966 856
rect 54134 2 54886 856
rect 55054 2 55898 856
rect 56066 2 56818 856
rect 56986 2 57738 856
rect 57906 2 58658 856
rect 58826 2 59670 856
rect 59838 2 60590 856
rect 60758 2 61510 856
rect 61678 2 62430 856
rect 62598 2 63350 856
rect 63518 2 64362 856
rect 64530 2 65282 856
rect 65450 2 66202 856
rect 66370 2 67122 856
rect 67290 2 68134 856
rect 68302 2 69054 856
rect 69222 2 69974 856
rect 70142 2 70894 856
rect 71062 2 71814 856
rect 71982 2 72826 856
rect 72994 2 73746 856
rect 73914 2 74666 856
rect 74834 2 75586 856
rect 75754 2 76598 856
rect 76766 2 77518 856
rect 77686 2 78438 856
rect 78606 2 79358 856
rect 79526 2 80278 856
rect 80446 2 81290 856
rect 81458 2 82210 856
rect 82378 2 83130 856
rect 83298 2 84050 856
rect 84218 2 85062 856
rect 85230 2 85982 856
rect 86150 2 86902 856
rect 87070 2 87822 856
rect 87990 2 88742 856
rect 88910 2 89754 856
rect 89922 2 90674 856
rect 90842 2 91594 856
rect 91762 2 92514 856
rect 92682 2 93526 856
rect 93694 2 94446 856
rect 94614 2 95366 856
rect 95534 2 96286 856
rect 96454 2 97206 856
rect 97374 2 98218 856
rect 98386 2 99138 856
rect 99306 2 100058 856
rect 100226 2 100978 856
rect 101146 2 101990 856
rect 102158 2 102910 856
rect 103078 2 103830 856
rect 103998 2 104750 856
rect 104918 2 105670 856
rect 105838 2 106682 856
rect 106850 2 107602 856
rect 107770 2 108522 856
rect 108690 2 109442 856
rect 109610 2 110454 856
rect 110622 2 111374 856
rect 111542 2 112294 856
rect 112462 2 113214 856
rect 113382 2 114134 856
rect 114302 2 115146 856
rect 115314 2 116066 856
rect 116234 2 116986 856
rect 117154 2 117906 856
rect 118074 2 118918 856
rect 119086 2 119838 856
rect 120006 2 120758 856
rect 120926 2 121678 856
rect 121846 2 122598 856
rect 122766 2 123610 856
rect 123778 2 124530 856
rect 124698 2 125450 856
rect 125618 2 126370 856
rect 126538 2 127382 856
rect 127550 2 128302 856
rect 128470 2 129222 856
rect 129390 2 130142 856
rect 130310 2 131062 856
rect 131230 2 132074 856
rect 132242 2 132994 856
rect 133162 2 133914 856
rect 134082 2 134834 856
rect 135002 2 135846 856
rect 136014 2 136766 856
rect 136934 2 137686 856
rect 137854 2 138606 856
rect 138774 2 139526 856
rect 139694 2 140538 856
rect 140706 2 141458 856
rect 141626 2 142378 856
rect 142546 2 143298 856
rect 143466 2 144310 856
rect 144478 2 145230 856
rect 145398 2 146150 856
rect 146318 2 147070 856
rect 147238 2 147990 856
rect 148158 2 149002 856
rect 149170 2 149922 856
rect 150090 2 150842 856
rect 151010 2 151762 856
rect 151930 2 152774 856
rect 152942 2 153694 856
rect 153862 2 154614 856
rect 154782 2 155534 856
rect 155702 2 156454 856
rect 156622 2 157466 856
rect 157634 2 158386 856
rect 158554 2 159306 856
rect 159474 2 160226 856
rect 160394 2 161238 856
rect 161406 2 162158 856
rect 162326 2 163006 856
<< metal3 >>
rect 0 165248 800 165368
rect 163813 165248 164613 165368
rect 0 162392 800 162512
rect 163813 162528 164613 162648
rect 163813 159808 164613 159928
rect 0 159536 800 159656
rect 163813 157088 164613 157208
rect 0 156680 800 156800
rect 163813 154504 164613 154624
rect 0 153960 800 154080
rect 163813 151784 164613 151904
rect 0 151104 800 151224
rect 163813 149064 164613 149184
rect 0 148248 800 148368
rect 163813 146344 164613 146464
rect 0 145392 800 145512
rect 163813 143760 164613 143880
rect 0 142536 800 142656
rect 163813 141040 164613 141160
rect 0 139816 800 139936
rect 163813 138320 164613 138440
rect 0 136960 800 137080
rect 163813 135600 164613 135720
rect 0 134104 800 134224
rect 163813 132880 164613 133000
rect 0 131248 800 131368
rect 163813 130296 164613 130416
rect 0 128528 800 128648
rect 163813 127576 164613 127696
rect 0 125672 800 125792
rect 163813 124856 164613 124976
rect 0 122816 800 122936
rect 163813 122136 164613 122256
rect 0 119960 800 120080
rect 163813 119552 164613 119672
rect 0 117104 800 117224
rect 163813 116832 164613 116952
rect 0 114384 800 114504
rect 163813 114112 164613 114232
rect 0 111528 800 111648
rect 163813 111392 164613 111512
rect 0 108672 800 108792
rect 163813 108672 164613 108792
rect 163813 106088 164613 106208
rect 0 105816 800 105936
rect 163813 103368 164613 103488
rect 0 103096 800 103216
rect 163813 100648 164613 100768
rect 0 100240 800 100360
rect 163813 97928 164613 98048
rect 0 97384 800 97504
rect 163813 95344 164613 95464
rect 0 94528 800 94648
rect 163813 92624 164613 92744
rect 0 91672 800 91792
rect 163813 89904 164613 90024
rect 0 88952 800 89072
rect 163813 87184 164613 87304
rect 0 86096 800 86216
rect 163813 84600 164613 84720
rect 0 83240 800 83360
rect 163813 81880 164613 82000
rect 0 80384 800 80504
rect 163813 79160 164613 79280
rect 0 77664 800 77784
rect 163813 76440 164613 76560
rect 0 74808 800 74928
rect 163813 73720 164613 73840
rect 0 71952 800 72072
rect 163813 71136 164613 71256
rect 0 69096 800 69216
rect 163813 68416 164613 68536
rect 0 66240 800 66360
rect 163813 65696 164613 65816
rect 0 63520 800 63640
rect 163813 62976 164613 63096
rect 0 60664 800 60784
rect 163813 60392 164613 60512
rect 0 57808 800 57928
rect 163813 57672 164613 57792
rect 0 54952 800 55072
rect 163813 54952 164613 55072
rect 0 52232 800 52352
rect 163813 52232 164613 52352
rect 0 49376 800 49496
rect 163813 49512 164613 49632
rect 163813 46928 164613 47048
rect 0 46520 800 46640
rect 163813 44208 164613 44328
rect 0 43664 800 43784
rect 163813 41488 164613 41608
rect 0 40808 800 40928
rect 163813 38768 164613 38888
rect 0 38088 800 38208
rect 163813 36184 164613 36304
rect 0 35232 800 35352
rect 163813 33464 164613 33584
rect 0 32376 800 32496
rect 163813 30744 164613 30864
rect 0 29520 800 29640
rect 163813 28024 164613 28144
rect 0 26800 800 26920
rect 163813 25304 164613 25424
rect 0 23944 800 24064
rect 163813 22720 164613 22840
rect 0 21088 800 21208
rect 163813 20000 164613 20120
rect 0 18232 800 18352
rect 163813 17280 164613 17400
rect 0 15376 800 15496
rect 163813 14560 164613 14680
rect 0 12656 800 12776
rect 163813 11976 164613 12096
rect 0 9800 800 9920
rect 163813 9256 164613 9376
rect 0 6944 800 7064
rect 163813 6536 164613 6656
rect 0 4088 800 4208
rect 163813 3816 164613 3936
rect 0 1368 800 1488
rect 163813 1232 164613 1352
<< obsm3 >>
rect 880 165168 163733 165341
rect 238 162728 163813 165168
rect 238 162592 163733 162728
rect 880 162448 163733 162592
rect 880 162312 163813 162448
rect 238 160008 163813 162312
rect 238 159736 163733 160008
rect 880 159728 163733 159736
rect 880 159456 163813 159728
rect 238 157288 163813 159456
rect 238 157008 163733 157288
rect 238 156880 163813 157008
rect 880 156600 163813 156880
rect 238 154704 163813 156600
rect 238 154424 163733 154704
rect 238 154160 163813 154424
rect 880 153880 163813 154160
rect 238 151984 163813 153880
rect 238 151704 163733 151984
rect 238 151304 163813 151704
rect 880 151024 163813 151304
rect 238 149264 163813 151024
rect 238 148984 163733 149264
rect 238 148448 163813 148984
rect 880 148168 163813 148448
rect 238 146544 163813 148168
rect 238 146264 163733 146544
rect 238 145592 163813 146264
rect 880 145312 163813 145592
rect 238 143960 163813 145312
rect 238 143680 163733 143960
rect 238 142736 163813 143680
rect 880 142456 163813 142736
rect 238 141240 163813 142456
rect 238 140960 163733 141240
rect 238 140016 163813 140960
rect 880 139736 163813 140016
rect 238 138520 163813 139736
rect 238 138240 163733 138520
rect 238 137160 163813 138240
rect 880 136880 163813 137160
rect 238 135800 163813 136880
rect 238 135520 163733 135800
rect 238 134304 163813 135520
rect 880 134024 163813 134304
rect 238 133080 163813 134024
rect 238 132800 163733 133080
rect 238 131448 163813 132800
rect 880 131168 163813 131448
rect 238 130496 163813 131168
rect 238 130216 163733 130496
rect 238 128728 163813 130216
rect 880 128448 163813 128728
rect 238 127776 163813 128448
rect 238 127496 163733 127776
rect 238 125872 163813 127496
rect 880 125592 163813 125872
rect 238 125056 163813 125592
rect 238 124776 163733 125056
rect 238 123016 163813 124776
rect 880 122736 163813 123016
rect 238 122336 163813 122736
rect 238 122056 163733 122336
rect 238 120160 163813 122056
rect 880 119880 163813 120160
rect 238 119752 163813 119880
rect 238 119472 163733 119752
rect 238 117304 163813 119472
rect 880 117032 163813 117304
rect 880 117024 163733 117032
rect 238 116752 163733 117024
rect 238 114584 163813 116752
rect 880 114312 163813 114584
rect 880 114304 163733 114312
rect 238 114032 163733 114304
rect 238 111728 163813 114032
rect 880 111592 163813 111728
rect 880 111448 163733 111592
rect 238 111312 163733 111448
rect 238 108872 163813 111312
rect 880 108592 163733 108872
rect 238 106288 163813 108592
rect 238 106016 163733 106288
rect 880 106008 163733 106016
rect 880 105736 163813 106008
rect 238 103568 163813 105736
rect 238 103296 163733 103568
rect 880 103288 163733 103296
rect 880 103016 163813 103288
rect 238 100848 163813 103016
rect 238 100568 163733 100848
rect 238 100440 163813 100568
rect 880 100160 163813 100440
rect 238 98128 163813 100160
rect 238 97848 163733 98128
rect 238 97584 163813 97848
rect 880 97304 163813 97584
rect 238 95544 163813 97304
rect 238 95264 163733 95544
rect 238 94728 163813 95264
rect 880 94448 163813 94728
rect 238 92824 163813 94448
rect 238 92544 163733 92824
rect 238 91872 163813 92544
rect 880 91592 163813 91872
rect 238 90104 163813 91592
rect 238 89824 163733 90104
rect 238 89152 163813 89824
rect 880 88872 163813 89152
rect 238 87384 163813 88872
rect 238 87104 163733 87384
rect 238 86296 163813 87104
rect 880 86016 163813 86296
rect 238 84800 163813 86016
rect 238 84520 163733 84800
rect 238 83440 163813 84520
rect 880 83160 163813 83440
rect 238 82080 163813 83160
rect 238 81800 163733 82080
rect 238 80584 163813 81800
rect 880 80304 163813 80584
rect 238 79360 163813 80304
rect 238 79080 163733 79360
rect 238 77864 163813 79080
rect 880 77584 163813 77864
rect 238 76640 163813 77584
rect 238 76360 163733 76640
rect 238 75008 163813 76360
rect 880 74728 163813 75008
rect 238 73920 163813 74728
rect 238 73640 163733 73920
rect 238 72152 163813 73640
rect 880 71872 163813 72152
rect 238 71336 163813 71872
rect 238 71056 163733 71336
rect 238 69296 163813 71056
rect 880 69016 163813 69296
rect 238 68616 163813 69016
rect 238 68336 163733 68616
rect 238 66440 163813 68336
rect 880 66160 163813 66440
rect 238 65896 163813 66160
rect 238 65616 163733 65896
rect 238 63720 163813 65616
rect 880 63440 163813 63720
rect 238 63176 163813 63440
rect 238 62896 163733 63176
rect 238 60864 163813 62896
rect 880 60592 163813 60864
rect 880 60584 163733 60592
rect 238 60312 163733 60584
rect 238 58008 163813 60312
rect 880 57872 163813 58008
rect 880 57728 163733 57872
rect 238 57592 163733 57728
rect 238 55152 163813 57592
rect 880 54872 163733 55152
rect 238 52432 163813 54872
rect 880 52152 163733 52432
rect 238 49712 163813 52152
rect 238 49576 163733 49712
rect 880 49432 163733 49576
rect 880 49296 163813 49432
rect 238 47128 163813 49296
rect 238 46848 163733 47128
rect 238 46720 163813 46848
rect 880 46440 163813 46720
rect 238 44408 163813 46440
rect 238 44128 163733 44408
rect 238 43864 163813 44128
rect 880 43584 163813 43864
rect 238 41688 163813 43584
rect 238 41408 163733 41688
rect 238 41008 163813 41408
rect 880 40728 163813 41008
rect 238 38968 163813 40728
rect 238 38688 163733 38968
rect 238 38288 163813 38688
rect 880 38008 163813 38288
rect 238 36384 163813 38008
rect 238 36104 163733 36384
rect 238 35432 163813 36104
rect 880 35152 163813 35432
rect 238 33664 163813 35152
rect 238 33384 163733 33664
rect 238 32576 163813 33384
rect 880 32296 163813 32576
rect 238 30944 163813 32296
rect 238 30664 163733 30944
rect 238 29720 163813 30664
rect 880 29440 163813 29720
rect 238 28224 163813 29440
rect 238 27944 163733 28224
rect 238 27000 163813 27944
rect 880 26720 163813 27000
rect 238 25504 163813 26720
rect 238 25224 163733 25504
rect 238 24144 163813 25224
rect 880 23864 163813 24144
rect 238 22920 163813 23864
rect 238 22640 163733 22920
rect 238 21288 163813 22640
rect 880 21008 163813 21288
rect 238 20200 163813 21008
rect 238 19920 163733 20200
rect 238 18432 163813 19920
rect 880 18152 163813 18432
rect 238 17480 163813 18152
rect 238 17200 163733 17480
rect 238 15576 163813 17200
rect 880 15296 163813 15576
rect 238 14760 163813 15296
rect 238 14480 163733 14760
rect 238 12856 163813 14480
rect 880 12576 163813 12856
rect 238 12176 163813 12576
rect 238 11896 163733 12176
rect 238 10000 163813 11896
rect 880 9720 163813 10000
rect 238 9456 163813 9720
rect 238 9176 163733 9456
rect 238 7144 163813 9176
rect 880 6864 163813 7144
rect 238 6736 163813 6864
rect 238 6456 163733 6736
rect 238 4288 163813 6456
rect 880 4016 163813 4288
rect 880 4008 163733 4016
rect 238 3736 163733 4008
rect 238 1568 163813 3736
rect 880 1432 163813 1568
rect 880 1288 163733 1432
rect 238 1152 163733 1288
rect 238 35 163813 1152
<< metal4 >>
rect 4208 2128 4528 164336
rect 19568 2128 19888 164336
rect 34928 2128 35248 164336
rect 50288 2128 50608 164336
rect 65648 2128 65968 164336
rect 81008 2128 81328 164336
rect 96368 2128 96688 164336
rect 111728 2128 112048 164336
rect 127088 2128 127408 164336
rect 142448 2128 142768 164336
rect 157808 2128 158128 164336
<< obsm4 >>
rect 243 2048 4128 164117
rect 4608 2048 19488 164117
rect 19968 2048 34848 164117
rect 35328 2048 50208 164117
rect 50688 2048 65568 164117
rect 66048 2048 80928 164117
rect 81408 2048 96288 164117
rect 96768 2048 111648 164117
rect 112128 2048 127008 164117
rect 127488 2048 141069 164117
rect 243 443 141069 2048
<< labels >>
rlabel metal3 s 0 1368 800 1488 6 i_dout0[0]
port 1 nsew signal input
rlabel metal2 s 133970 0 134026 800 6 i_dout0[10]
port 2 nsew signal input
rlabel metal3 s 163813 89904 164613 90024 6 i_dout0[11]
port 3 nsew signal input
rlabel metal2 s 135810 165957 135866 166757 6 i_dout0[12]
port 4 nsew signal input
rlabel metal3 s 163813 100648 164613 100768 6 i_dout0[13]
port 5 nsew signal input
rlabel metal3 s 0 86096 800 86216 6 i_dout0[14]
port 6 nsew signal input
rlabel metal2 s 139674 165957 139730 166757 6 i_dout0[15]
port 7 nsew signal input
rlabel metal3 s 163813 111392 164613 111512 6 i_dout0[16]
port 8 nsew signal input
rlabel metal2 s 142434 0 142490 800 6 i_dout0[17]
port 9 nsew signal input
rlabel metal2 s 142618 165957 142674 166757 6 i_dout0[18]
port 10 nsew signal input
rlabel metal2 s 144550 165957 144606 166757 6 i_dout0[19]
port 11 nsew signal input
rlabel metal2 s 114374 165957 114430 166757 6 i_dout0[1]
port 12 nsew signal input
rlabel metal2 s 146482 165957 146538 166757 6 i_dout0[20]
port 13 nsew signal input
rlabel metal3 s 0 119960 800 120080 6 i_dout0[21]
port 14 nsew signal input
rlabel metal3 s 0 122816 800 122936 6 i_dout0[22]
port 15 nsew signal input
rlabel metal2 s 149978 0 150034 800 6 i_dout0[23]
port 16 nsew signal input
rlabel metal3 s 0 131248 800 131368 6 i_dout0[24]
port 17 nsew signal input
rlabel metal3 s 163813 141040 164613 141160 6 i_dout0[25]
port 18 nsew signal input
rlabel metal2 s 153750 0 153806 800 6 i_dout0[26]
port 19 nsew signal input
rlabel metal3 s 0 142536 800 142656 6 i_dout0[27]
port 20 nsew signal input
rlabel metal2 s 157522 0 157578 800 6 i_dout0[28]
port 21 nsew signal input
rlabel metal2 s 158442 0 158498 800 6 i_dout0[29]
port 22 nsew signal input
rlabel metal3 s 163813 22720 164613 22840 6 i_dout0[2]
port 23 nsew signal input
rlabel metal3 s 163813 162528 164613 162648 6 i_dout0[30]
port 24 nsew signal input
rlabel metal3 s 0 162392 800 162512 6 i_dout0[31]
port 25 nsew signal input
rlabel metal3 s 0 26800 800 26920 6 i_dout0[3]
port 26 nsew signal input
rlabel metal2 s 121734 0 121790 800 6 i_dout0[4]
port 27 nsew signal input
rlabel metal3 s 163813 49512 164613 49632 6 i_dout0[5]
port 28 nsew signal input
rlabel metal2 s 128358 0 128414 800 6 i_dout0[6]
port 29 nsew signal input
rlabel metal2 s 125046 165957 125102 166757 6 i_dout0[7]
port 30 nsew signal input
rlabel metal3 s 0 60664 800 60784 6 i_dout0[8]
port 31 nsew signal input
rlabel metal3 s 163813 79160 164613 79280 6 i_dout0[9]
port 32 nsew signal input
rlabel metal3 s 163813 3816 164613 3936 6 i_dout0_1[0]
port 33 nsew signal input
rlabel metal2 s 133050 0 133106 800 6 i_dout0_1[10]
port 34 nsew signal input
rlabel metal3 s 163813 87184 164613 87304 6 i_dout0_1[11]
port 35 nsew signal input
rlabel metal2 s 134798 165957 134854 166757 6 i_dout0_1[12]
port 36 nsew signal input
rlabel metal3 s 163813 97928 164613 98048 6 i_dout0_1[13]
port 37 nsew signal input
rlabel metal2 s 138662 0 138718 800 6 i_dout0_1[14]
port 38 nsew signal input
rlabel metal3 s 0 91672 800 91792 6 i_dout0_1[15]
port 39 nsew signal input
rlabel metal3 s 163813 108672 164613 108792 6 i_dout0_1[16]
port 40 nsew signal input
rlabel metal3 s 0 100240 800 100360 6 i_dout0_1[17]
port 41 nsew signal input
rlabel metal3 s 0 105816 800 105936 6 i_dout0_1[18]
port 42 nsew signal input
rlabel metal2 s 145286 0 145342 800 6 i_dout0_1[19]
port 43 nsew signal input
rlabel metal2 s 110510 0 110566 800 6 i_dout0_1[1]
port 44 nsew signal input
rlabel metal2 s 147126 0 147182 800 6 i_dout0_1[20]
port 45 nsew signal input
rlabel metal3 s 163813 124856 164613 124976 6 i_dout0_1[21]
port 46 nsew signal input
rlabel metal3 s 163813 130296 164613 130416 6 i_dout0_1[22]
port 47 nsew signal input
rlabel metal2 s 149058 0 149114 800 6 i_dout0_1[23]
port 48 nsew signal input
rlabel metal2 s 155314 165957 155370 166757 6 i_dout0_1[24]
port 49 nsew signal input
rlabel metal3 s 163813 138320 164613 138440 6 i_dout0_1[25]
port 50 nsew signal input
rlabel metal3 s 163813 146344 164613 146464 6 i_dout0_1[26]
port 51 nsew signal input
rlabel metal2 s 155590 0 155646 800 6 i_dout0_1[27]
port 52 nsew signal input
rlabel metal3 s 0 148248 800 148368 6 i_dout0_1[28]
port 53 nsew signal input
rlabel metal2 s 162122 165957 162178 166757 6 i_dout0_1[29]
port 54 nsew signal input
rlabel metal3 s 163813 20000 164613 20120 6 i_dout0_1[2]
port 55 nsew signal input
rlabel metal3 s 163813 159808 164613 159928 6 i_dout0_1[30]
port 56 nsew signal input
rlabel metal2 s 163134 0 163190 800 6 i_dout0_1[31]
port 57 nsew signal input
rlabel metal3 s 0 23944 800 24064 6 i_dout0_1[3]
port 58 nsew signal input
rlabel metal3 s 163813 38768 164613 38888 6 i_dout0_1[4]
port 59 nsew signal input
rlabel metal2 s 120262 165957 120318 166757 6 i_dout0_1[5]
port 60 nsew signal input
rlabel metal2 s 122194 165957 122250 166757 6 i_dout0_1[6]
port 61 nsew signal input
rlabel metal3 s 163813 65696 164613 65816 6 i_dout0_1[7]
port 62 nsew signal input
rlabel metal2 s 131118 0 131174 800 6 i_dout0_1[8]
port 63 nsew signal input
rlabel metal2 s 129002 165957 129058 166757 6 i_dout0_1[9]
port 64 nsew signal input
rlabel metal2 s 112442 165957 112498 166757 6 i_dout1[0]
port 65 nsew signal input
rlabel metal3 s 0 77664 800 77784 6 i_dout1[10]
port 66 nsew signal input
rlabel metal3 s 163813 92624 164613 92744 6 i_dout1[11]
port 67 nsew signal input
rlabel metal2 s 135902 0 135958 800 6 i_dout1[12]
port 68 nsew signal input
rlabel metal2 s 136822 0 136878 800 6 i_dout1[13]
port 69 nsew signal input
rlabel metal3 s 0 88952 800 89072 6 i_dout1[14]
port 70 nsew signal input
rlabel metal2 s 140686 165957 140742 166757 6 i_dout1[15]
port 71 nsew signal input
rlabel metal3 s 0 97384 800 97504 6 i_dout1[16]
port 72 nsew signal input
rlabel metal2 s 143354 0 143410 800 6 i_dout1[17]
port 73 nsew signal input
rlabel metal3 s 0 108672 800 108792 6 i_dout1[18]
port 74 nsew signal input
rlabel metal2 s 146206 0 146262 800 6 i_dout1[19]
port 75 nsew signal input
rlabel metal3 s 163813 11976 164613 12096 6 i_dout1[1]
port 76 nsew signal input
rlabel metal2 s 147494 165957 147550 166757 6 i_dout1[20]
port 77 nsew signal input
rlabel metal2 s 148046 0 148102 800 6 i_dout1[21]
port 78 nsew signal input
rlabel metal3 s 163813 132880 164613 133000 6 i_dout1[22]
port 79 nsew signal input
rlabel metal3 s 0 128528 800 128648 6 i_dout1[23]
port 80 nsew signal input
rlabel metal3 s 0 134104 800 134224 6 i_dout1[24]
port 81 nsew signal input
rlabel metal3 s 0 136960 800 137080 6 i_dout1[25]
port 82 nsew signal input
rlabel metal2 s 158166 165957 158222 166757 6 i_dout1[26]
port 83 nsew signal input
rlabel metal3 s 163813 154504 164613 154624 6 i_dout1[27]
port 84 nsew signal input
rlabel metal3 s 0 151104 800 151224 6 i_dout1[28]
port 85 nsew signal input
rlabel metal2 s 163042 165957 163098 166757 6 i_dout1[29]
port 86 nsew signal input
rlabel metal3 s 0 15376 800 15496 6 i_dout1[2]
port 87 nsew signal input
rlabel metal2 s 164054 165957 164110 166757 6 i_dout1[30]
port 88 nsew signal input
rlabel metal2 s 164054 0 164110 800 6 i_dout1[31]
port 89 nsew signal input
rlabel metal2 s 118974 0 119030 800 6 i_dout1[3]
port 90 nsew signal input
rlabel metal3 s 163813 44208 164613 44328 6 i_dout1[4]
port 91 nsew signal input
rlabel metal3 s 163813 52232 164613 52352 6 i_dout1[5]
port 92 nsew signal input
rlabel metal2 s 123114 165957 123170 166757 6 i_dout1[6]
port 93 nsew signal input
rlabel metal2 s 126058 165957 126114 166757 6 i_dout1[7]
port 94 nsew signal input
rlabel metal3 s 163813 71136 164613 71256 6 i_dout1[8]
port 95 nsew signal input
rlabel metal2 s 130934 165957 130990 166757 6 i_dout1[9]
port 96 nsew signal input
rlabel metal3 s 0 4088 800 4208 6 i_dout1_1[0]
port 97 nsew signal input
rlabel metal3 s 0 74808 800 74928 6 i_dout1_1[10]
port 98 nsew signal input
rlabel metal2 s 132866 165957 132922 166757 6 i_dout1_1[11]
port 99 nsew signal input
rlabel metal2 s 134890 0 134946 800 6 i_dout1_1[12]
port 100 nsew signal input
rlabel metal2 s 136822 165957 136878 166757 6 i_dout1_1[13]
port 101 nsew signal input
rlabel metal3 s 163813 103368 164613 103488 6 i_dout1_1[14]
port 102 nsew signal input
rlabel metal3 s 163813 106088 164613 106208 6 i_dout1_1[15]
port 103 nsew signal input
rlabel metal3 s 0 94528 800 94648 6 i_dout1_1[16]
port 104 nsew signal input
rlabel metal3 s 0 103096 800 103216 6 i_dout1_1[17]
port 105 nsew signal input
rlabel metal3 s 163813 119552 164613 119672 6 i_dout1_1[18]
port 106 nsew signal input
rlabel metal3 s 0 114384 800 114504 6 i_dout1_1[19]
port 107 nsew signal input
rlabel metal3 s 0 9800 800 9920 6 i_dout1_1[1]
port 108 nsew signal input
rlabel metal3 s 0 117104 800 117224 6 i_dout1_1[20]
port 109 nsew signal input
rlabel metal3 s 163813 127576 164613 127696 6 i_dout1_1[21]
port 110 nsew signal input
rlabel metal2 s 152370 165957 152426 166757 6 i_dout1_1[22]
port 111 nsew signal input
rlabel metal3 s 0 125672 800 125792 6 i_dout1_1[23]
port 112 nsew signal input
rlabel metal3 s 163813 135600 164613 135720 6 i_dout1_1[24]
port 113 nsew signal input
rlabel metal2 s 152830 0 152886 800 6 i_dout1_1[25]
port 114 nsew signal input
rlabel metal3 s 163813 149064 164613 149184 6 i_dout1_1[26]
port 115 nsew signal input
rlabel metal3 s 163813 151784 164613 151904 6 i_dout1_1[27]
port 116 nsew signal input
rlabel metal2 s 160190 165957 160246 166757 6 i_dout1_1[28]
port 117 nsew signal input
rlabel metal3 s 163813 157088 164613 157208 6 i_dout1_1[29]
port 118 nsew signal input
rlabel metal2 s 116122 0 116178 800 6 i_dout1_1[2]
port 119 nsew signal input
rlabel metal2 s 161294 0 161350 800 6 i_dout1_1[30]
port 120 nsew signal input
rlabel metal3 s 0 159536 800 159656 6 i_dout1_1[31]
port 121 nsew signal input
rlabel metal2 s 117962 0 118018 800 6 i_dout1_1[3]
port 122 nsew signal input
rlabel metal3 s 163813 41488 164613 41608 6 i_dout1_1[4]
port 123 nsew signal input
rlabel metal3 s 0 38088 800 38208 6 i_dout1_1[5]
port 124 nsew signal input
rlabel metal3 s 0 43664 800 43784 6 i_dout1_1[6]
port 125 nsew signal input
rlabel metal3 s 0 52232 800 52352 6 i_dout1_1[7]
port 126 nsew signal input
rlabel metal2 s 132130 0 132186 800 6 i_dout1_1[8]
port 127 nsew signal input
rlabel metal2 s 129922 165957 129978 166757 6 i_dout1_1[9]
port 128 nsew signal input
rlabel metal2 s 478 165957 534 166757 6 io_in[0]
port 129 nsew signal input
rlabel metal2 s 29642 165957 29698 166757 6 io_in[10]
port 130 nsew signal input
rlabel metal2 s 32586 165957 32642 166757 6 io_in[11]
port 131 nsew signal input
rlabel metal2 s 35530 165957 35586 166757 6 io_in[12]
port 132 nsew signal input
rlabel metal2 s 38382 165957 38438 166757 6 io_in[13]
port 133 nsew signal input
rlabel metal2 s 41326 165957 41382 166757 6 io_in[14]
port 134 nsew signal input
rlabel metal2 s 44270 165957 44326 166757 6 io_in[15]
port 135 nsew signal input
rlabel metal2 s 47214 165957 47270 166757 6 io_in[16]
port 136 nsew signal input
rlabel metal2 s 50066 165957 50122 166757 6 io_in[17]
port 137 nsew signal input
rlabel metal2 s 53010 165957 53066 166757 6 io_in[18]
port 138 nsew signal input
rlabel metal2 s 55954 165957 56010 166757 6 io_in[19]
port 139 nsew signal input
rlabel metal2 s 3330 165957 3386 166757 6 io_in[1]
port 140 nsew signal input
rlabel metal2 s 58898 165957 58954 166757 6 io_in[20]
port 141 nsew signal input
rlabel metal2 s 61750 165957 61806 166757 6 io_in[21]
port 142 nsew signal input
rlabel metal2 s 64694 165957 64750 166757 6 io_in[22]
port 143 nsew signal input
rlabel metal2 s 67638 165957 67694 166757 6 io_in[23]
port 144 nsew signal input
rlabel metal2 s 70582 165957 70638 166757 6 io_in[24]
port 145 nsew signal input
rlabel metal2 s 73434 165957 73490 166757 6 io_in[25]
port 146 nsew signal input
rlabel metal2 s 76378 165957 76434 166757 6 io_in[26]
port 147 nsew signal input
rlabel metal2 s 79322 165957 79378 166757 6 io_in[27]
port 148 nsew signal input
rlabel metal2 s 82266 165957 82322 166757 6 io_in[28]
port 149 nsew signal input
rlabel metal2 s 85118 165957 85174 166757 6 io_in[29]
port 150 nsew signal input
rlabel metal2 s 6274 165957 6330 166757 6 io_in[2]
port 151 nsew signal input
rlabel metal2 s 88062 165957 88118 166757 6 io_in[30]
port 152 nsew signal input
rlabel metal2 s 91006 165957 91062 166757 6 io_in[31]
port 153 nsew signal input
rlabel metal2 s 93950 165957 94006 166757 6 io_in[32]
port 154 nsew signal input
rlabel metal2 s 96802 165957 96858 166757 6 io_in[33]
port 155 nsew signal input
rlabel metal2 s 99746 165957 99802 166757 6 io_in[34]
port 156 nsew signal input
rlabel metal2 s 102690 165957 102746 166757 6 io_in[35]
port 157 nsew signal input
rlabel metal2 s 105634 165957 105690 166757 6 io_in[36]
port 158 nsew signal input
rlabel metal2 s 108578 165957 108634 166757 6 io_in[37]
port 159 nsew signal input
rlabel metal2 s 9218 165957 9274 166757 6 io_in[3]
port 160 nsew signal input
rlabel metal2 s 12162 165957 12218 166757 6 io_in[4]
port 161 nsew signal input
rlabel metal2 s 15014 165957 15070 166757 6 io_in[5]
port 162 nsew signal input
rlabel metal2 s 17958 165957 18014 166757 6 io_in[6]
port 163 nsew signal input
rlabel metal2 s 20902 165957 20958 166757 6 io_in[7]
port 164 nsew signal input
rlabel metal2 s 23846 165957 23902 166757 6 io_in[8]
port 165 nsew signal input
rlabel metal2 s 26698 165957 26754 166757 6 io_in[9]
port 166 nsew signal input
rlabel metal2 s 1398 165957 1454 166757 6 io_oeb[0]
port 167 nsew signal output
rlabel metal2 s 30654 165957 30710 166757 6 io_oeb[10]
port 168 nsew signal output
rlabel metal2 s 33506 165957 33562 166757 6 io_oeb[11]
port 169 nsew signal output
rlabel metal2 s 36450 165957 36506 166757 6 io_oeb[12]
port 170 nsew signal output
rlabel metal2 s 39394 165957 39450 166757 6 io_oeb[13]
port 171 nsew signal output
rlabel metal2 s 42338 165957 42394 166757 6 io_oeb[14]
port 172 nsew signal output
rlabel metal2 s 45190 165957 45246 166757 6 io_oeb[15]
port 173 nsew signal output
rlabel metal2 s 48134 165957 48190 166757 6 io_oeb[16]
port 174 nsew signal output
rlabel metal2 s 51078 165957 51134 166757 6 io_oeb[17]
port 175 nsew signal output
rlabel metal2 s 54022 165957 54078 166757 6 io_oeb[18]
port 176 nsew signal output
rlabel metal2 s 56874 165957 56930 166757 6 io_oeb[19]
port 177 nsew signal output
rlabel metal2 s 4342 165957 4398 166757 6 io_oeb[1]
port 178 nsew signal output
rlabel metal2 s 59818 165957 59874 166757 6 io_oeb[20]
port 179 nsew signal output
rlabel metal2 s 62762 165957 62818 166757 6 io_oeb[21]
port 180 nsew signal output
rlabel metal2 s 65706 165957 65762 166757 6 io_oeb[22]
port 181 nsew signal output
rlabel metal2 s 68650 165957 68706 166757 6 io_oeb[23]
port 182 nsew signal output
rlabel metal2 s 71502 165957 71558 166757 6 io_oeb[24]
port 183 nsew signal output
rlabel metal2 s 74446 165957 74502 166757 6 io_oeb[25]
port 184 nsew signal output
rlabel metal2 s 77390 165957 77446 166757 6 io_oeb[26]
port 185 nsew signal output
rlabel metal2 s 80334 165957 80390 166757 6 io_oeb[27]
port 186 nsew signal output
rlabel metal2 s 83186 165957 83242 166757 6 io_oeb[28]
port 187 nsew signal output
rlabel metal2 s 86130 165957 86186 166757 6 io_oeb[29]
port 188 nsew signal output
rlabel metal2 s 7286 165957 7342 166757 6 io_oeb[2]
port 189 nsew signal output
rlabel metal2 s 89074 165957 89130 166757 6 io_oeb[30]
port 190 nsew signal output
rlabel metal2 s 92018 165957 92074 166757 6 io_oeb[31]
port 191 nsew signal output
rlabel metal2 s 94870 165957 94926 166757 6 io_oeb[32]
port 192 nsew signal output
rlabel metal2 s 97814 165957 97870 166757 6 io_oeb[33]
port 193 nsew signal output
rlabel metal2 s 100758 165957 100814 166757 6 io_oeb[34]
port 194 nsew signal output
rlabel metal2 s 103702 165957 103758 166757 6 io_oeb[35]
port 195 nsew signal output
rlabel metal2 s 106554 165957 106610 166757 6 io_oeb[36]
port 196 nsew signal output
rlabel metal2 s 109498 165957 109554 166757 6 io_oeb[37]
port 197 nsew signal output
rlabel metal2 s 10138 165957 10194 166757 6 io_oeb[3]
port 198 nsew signal output
rlabel metal2 s 13082 165957 13138 166757 6 io_oeb[4]
port 199 nsew signal output
rlabel metal2 s 16026 165957 16082 166757 6 io_oeb[5]
port 200 nsew signal output
rlabel metal2 s 18970 165957 19026 166757 6 io_oeb[6]
port 201 nsew signal output
rlabel metal2 s 21822 165957 21878 166757 6 io_oeb[7]
port 202 nsew signal output
rlabel metal2 s 24766 165957 24822 166757 6 io_oeb[8]
port 203 nsew signal output
rlabel metal2 s 27710 165957 27766 166757 6 io_oeb[9]
port 204 nsew signal output
rlabel metal2 s 2410 165957 2466 166757 6 io_out[0]
port 205 nsew signal output
rlabel metal2 s 31574 165957 31630 166757 6 io_out[10]
port 206 nsew signal output
rlabel metal2 s 34518 165957 34574 166757 6 io_out[11]
port 207 nsew signal output
rlabel metal2 s 37462 165957 37518 166757 6 io_out[12]
port 208 nsew signal output
rlabel metal2 s 40406 165957 40462 166757 6 io_out[13]
port 209 nsew signal output
rlabel metal2 s 43258 165957 43314 166757 6 io_out[14]
port 210 nsew signal output
rlabel metal2 s 46202 165957 46258 166757 6 io_out[15]
port 211 nsew signal output
rlabel metal2 s 49146 165957 49202 166757 6 io_out[16]
port 212 nsew signal output
rlabel metal2 s 52090 165957 52146 166757 6 io_out[17]
port 213 nsew signal output
rlabel metal2 s 54942 165957 54998 166757 6 io_out[18]
port 214 nsew signal output
rlabel metal2 s 57886 165957 57942 166757 6 io_out[19]
port 215 nsew signal output
rlabel metal2 s 5262 165957 5318 166757 6 io_out[1]
port 216 nsew signal output
rlabel metal2 s 60830 165957 60886 166757 6 io_out[20]
port 217 nsew signal output
rlabel metal2 s 63774 165957 63830 166757 6 io_out[21]
port 218 nsew signal output
rlabel metal2 s 66626 165957 66682 166757 6 io_out[22]
port 219 nsew signal output
rlabel metal2 s 69570 165957 69626 166757 6 io_out[23]
port 220 nsew signal output
rlabel metal2 s 72514 165957 72570 166757 6 io_out[24]
port 221 nsew signal output
rlabel metal2 s 75458 165957 75514 166757 6 io_out[25]
port 222 nsew signal output
rlabel metal2 s 78310 165957 78366 166757 6 io_out[26]
port 223 nsew signal output
rlabel metal2 s 81254 165957 81310 166757 6 io_out[27]
port 224 nsew signal output
rlabel metal2 s 84198 165957 84254 166757 6 io_out[28]
port 225 nsew signal output
rlabel metal2 s 87142 165957 87198 166757 6 io_out[29]
port 226 nsew signal output
rlabel metal2 s 8206 165957 8262 166757 6 io_out[2]
port 227 nsew signal output
rlabel metal2 s 89994 165957 90050 166757 6 io_out[30]
port 228 nsew signal output
rlabel metal2 s 92938 165957 92994 166757 6 io_out[31]
port 229 nsew signal output
rlabel metal2 s 95882 165957 95938 166757 6 io_out[32]
port 230 nsew signal output
rlabel metal2 s 98826 165957 98882 166757 6 io_out[33]
port 231 nsew signal output
rlabel metal2 s 101678 165957 101734 166757 6 io_out[34]
port 232 nsew signal output
rlabel metal2 s 104622 165957 104678 166757 6 io_out[35]
port 233 nsew signal output
rlabel metal2 s 107566 165957 107622 166757 6 io_out[36]
port 234 nsew signal output
rlabel metal2 s 110510 165957 110566 166757 6 io_out[37]
port 235 nsew signal output
rlabel metal2 s 11150 165957 11206 166757 6 io_out[3]
port 236 nsew signal output
rlabel metal2 s 14094 165957 14150 166757 6 io_out[4]
port 237 nsew signal output
rlabel metal2 s 16946 165957 17002 166757 6 io_out[5]
port 238 nsew signal output
rlabel metal2 s 19890 165957 19946 166757 6 io_out[6]
port 239 nsew signal output
rlabel metal2 s 22834 165957 22890 166757 6 io_out[7]
port 240 nsew signal output
rlabel metal2 s 25778 165957 25834 166757 6 io_out[8]
port 241 nsew signal output
rlabel metal2 s 28630 165957 28686 166757 6 io_out[9]
port 242 nsew signal output
rlabel metal2 s 100114 0 100170 800 6 irq[0]
port 243 nsew signal output
rlabel metal2 s 101034 0 101090 800 6 irq[1]
port 244 nsew signal output
rlabel metal2 s 102046 0 102102 800 6 irq[2]
port 245 nsew signal output
rlabel metal2 s 106738 0 106794 800 6 o_addr1[0]
port 246 nsew signal output
rlabel metal2 s 111430 0 111486 800 6 o_addr1[1]
port 247 nsew signal output
rlabel metal3 s 0 18232 800 18352 6 o_addr1[2]
port 248 nsew signal output
rlabel metal3 s 0 29520 800 29640 6 o_addr1[3]
port 249 nsew signal output
rlabel metal2 s 122654 0 122710 800 6 o_addr1[4]
port 250 nsew signal output
rlabel metal3 s 163813 54952 164613 55072 6 o_addr1[5]
port 251 nsew signal output
rlabel metal3 s 163813 60392 164613 60512 6 o_addr1[6]
port 252 nsew signal output
rlabel metal2 s 129278 0 129334 800 6 o_addr1[7]
port 253 nsew signal output
rlabel metal3 s 0 63520 800 63640 6 o_addr1[8]
port 254 nsew signal output
rlabel metal2 s 113362 165957 113418 166757 6 o_addr1_1[0]
port 255 nsew signal output
rlabel metal3 s 163813 14560 164613 14680 6 o_addr1_1[1]
port 256 nsew signal output
rlabel metal2 s 115386 165957 115442 166757 6 o_addr1_1[2]
port 257 nsew signal output
rlabel metal2 s 118238 165957 118294 166757 6 o_addr1_1[3]
port 258 nsew signal output
rlabel metal2 s 119250 165957 119306 166757 6 o_addr1_1[4]
port 259 nsew signal output
rlabel metal3 s 0 40808 800 40928 6 o_addr1_1[5]
port 260 nsew signal output
rlabel metal3 s 163813 57672 164613 57792 6 o_addr1_1[6]
port 261 nsew signal output
rlabel metal3 s 163813 68416 164613 68536 6 o_addr1_1[7]
port 262 nsew signal output
rlabel metal2 s 127990 165957 128046 166757 6 o_addr1_1[8]
port 263 nsew signal output
rlabel metal2 s 102966 0 103022 800 6 o_csb0
port 264 nsew signal output
rlabel metal2 s 111430 165957 111486 166757 6 o_csb0_1
port 265 nsew signal output
rlabel metal2 s 103886 0 103942 800 6 o_csb1
port 266 nsew signal output
rlabel metal3 s 163813 1232 164613 1352 6 o_csb1_1
port 267 nsew signal output
rlabel metal3 s 0 6944 800 7064 6 o_din0[0]
port 268 nsew signal output
rlabel metal2 s 131946 165957 132002 166757 6 o_din0[10]
port 269 nsew signal output
rlabel metal2 s 133878 165957 133934 166757 6 o_din0[11]
port 270 nsew signal output
rlabel metal3 s 0 83240 800 83360 6 o_din0[12]
port 271 nsew signal output
rlabel metal2 s 137742 165957 137798 166757 6 o_din0[13]
port 272 nsew signal output
rlabel metal2 s 139582 0 139638 800 6 o_din0[14]
port 273 nsew signal output
rlabel metal2 s 140594 0 140650 800 6 o_din0[15]
port 274 nsew signal output
rlabel metal3 s 163813 114112 164613 114232 6 o_din0[16]
port 275 nsew signal output
rlabel metal2 s 144366 0 144422 800 6 o_din0[17]
port 276 nsew signal output
rlabel metal2 s 143630 165957 143686 166757 6 o_din0[18]
port 277 nsew signal output
rlabel metal2 s 145562 165957 145618 166757 6 o_din0[19]
port 278 nsew signal output
rlabel metal2 s 113270 0 113326 800 6 o_din0[1]
port 279 nsew signal output
rlabel metal2 s 149426 165957 149482 166757 6 o_din0[20]
port 280 nsew signal output
rlabel metal2 s 151358 165957 151414 166757 6 o_din0[21]
port 281 nsew signal output
rlabel metal2 s 154302 165957 154358 166757 6 o_din0[22]
port 282 nsew signal output
rlabel metal2 s 151818 0 151874 800 6 o_din0[23]
port 283 nsew signal output
rlabel metal2 s 157246 165957 157302 166757 6 o_din0[24]
port 284 nsew signal output
rlabel metal3 s 0 139816 800 139936 6 o_din0[25]
port 285 nsew signal output
rlabel metal2 s 154670 0 154726 800 6 o_din0[26]
port 286 nsew signal output
rlabel metal2 s 156510 0 156566 800 6 o_din0[27]
port 287 nsew signal output
rlabel metal3 s 0 153960 800 154080 6 o_din0[28]
port 288 nsew signal output
rlabel metal2 s 160282 0 160338 800 6 o_din0[29]
port 289 nsew signal output
rlabel metal3 s 0 21088 800 21208 6 o_din0[2]
port 290 nsew signal output
rlabel metal3 s 0 156680 800 156800 6 o_din0[30]
port 291 nsew signal output
rlabel metal3 s 163813 165248 164613 165368 6 o_din0[31]
port 292 nsew signal output
rlabel metal3 s 0 32376 800 32496 6 o_din0[3]
port 293 nsew signal output
rlabel metal3 s 163813 46928 164613 47048 6 o_din0[4]
port 294 nsew signal output
rlabel metal2 s 121182 165957 121238 166757 6 o_din0[5]
port 295 nsew signal output
rlabel metal3 s 0 46520 800 46640 6 o_din0[6]
port 296 nsew signal output
rlabel metal3 s 0 54952 800 55072 6 o_din0[7]
port 297 nsew signal output
rlabel metal3 s 0 69096 800 69216 6 o_din0[8]
port 298 nsew signal output
rlabel metal3 s 0 71952 800 72072 6 o_din0[9]
port 299 nsew signal output
rlabel metal2 s 107658 0 107714 800 6 o_din0_1[0]
port 300 nsew signal output
rlabel metal3 s 163813 84600 164613 84720 6 o_din0_1[10]
port 301 nsew signal output
rlabel metal3 s 163813 95344 164613 95464 6 o_din0_1[11]
port 302 nsew signal output
rlabel metal3 s 0 80384 800 80504 6 o_din0_1[12]
port 303 nsew signal output
rlabel metal2 s 137742 0 137798 800 6 o_din0_1[13]
port 304 nsew signal output
rlabel metal2 s 138754 165957 138810 166757 6 o_din0_1[14]
port 305 nsew signal output
rlabel metal2 s 141606 165957 141662 166757 6 o_din0_1[15]
port 306 nsew signal output
rlabel metal2 s 141514 0 141570 800 6 o_din0_1[16]
port 307 nsew signal output
rlabel metal3 s 163813 116832 164613 116952 6 o_din0_1[17]
port 308 nsew signal output
rlabel metal3 s 0 111528 800 111648 6 o_din0_1[18]
port 309 nsew signal output
rlabel metal3 s 163813 122136 164613 122256 6 o_din0_1[19]
port 310 nsew signal output
rlabel metal2 s 112350 0 112406 800 6 o_din0_1[1]
port 311 nsew signal output
rlabel metal2 s 148506 165957 148562 166757 6 o_din0_1[20]
port 312 nsew signal output
rlabel metal2 s 150438 165957 150494 166757 6 o_din0_1[21]
port 313 nsew signal output
rlabel metal2 s 153290 165957 153346 166757 6 o_din0_1[22]
port 314 nsew signal output
rlabel metal2 s 150898 0 150954 800 6 o_din0_1[23]
port 315 nsew signal output
rlabel metal2 s 156234 165957 156290 166757 6 o_din0_1[24]
port 316 nsew signal output
rlabel metal3 s 163813 143760 164613 143880 6 o_din0_1[25]
port 317 nsew signal output
rlabel metal2 s 159178 165957 159234 166757 6 o_din0_1[26]
port 318 nsew signal output
rlabel metal3 s 0 145392 800 145512 6 o_din0_1[27]
port 319 nsew signal output
rlabel metal2 s 161110 165957 161166 166757 6 o_din0_1[28]
port 320 nsew signal output
rlabel metal2 s 159362 0 159418 800 6 o_din0_1[29]
port 321 nsew signal output
rlabel metal2 s 116306 165957 116362 166757 6 o_din0_1[2]
port 322 nsew signal output
rlabel metal2 s 162214 0 162270 800 6 o_din0_1[30]
port 323 nsew signal output
rlabel metal3 s 0 165248 800 165368 6 o_din0_1[31]
port 324 nsew signal output
rlabel metal2 s 119894 0 119950 800 6 o_din0_1[3]
port 325 nsew signal output
rlabel metal3 s 0 35232 800 35352 6 o_din0_1[4]
port 326 nsew signal output
rlabel metal2 s 125506 0 125562 800 6 o_din0_1[5]
port 327 nsew signal output
rlabel metal2 s 124126 165957 124182 166757 6 o_din0_1[6]
port 328 nsew signal output
rlabel metal2 s 127070 165957 127126 166757 6 o_din0_1[7]
port 329 nsew signal output
rlabel metal3 s 0 66240 800 66360 6 o_din0_1[8]
port 330 nsew signal output
rlabel metal3 s 163813 81880 164613 82000 6 o_din0_1[9]
port 331 nsew signal output
rlabel metal3 s 163813 6536 164613 6656 6 o_waddr0[0]
port 332 nsew signal output
rlabel metal3 s 0 12656 800 12776 6 o_waddr0[1]
port 333 nsew signal output
rlabel metal2 s 117042 0 117098 800 6 o_waddr0[2]
port 334 nsew signal output
rlabel metal3 s 163813 33464 164613 33584 6 o_waddr0[3]
port 335 nsew signal output
rlabel metal2 s 124586 0 124642 800 6 o_waddr0[4]
port 336 nsew signal output
rlabel metal2 s 127438 0 127494 800 6 o_waddr0[5]
port 337 nsew signal output
rlabel metal3 s 0 49376 800 49496 6 o_waddr0[6]
port 338 nsew signal output
rlabel metal3 s 0 57808 800 57928 6 o_waddr0[7]
port 339 nsew signal output
rlabel metal3 s 163813 76440 164613 76560 6 o_waddr0[8]
port 340 nsew signal output
rlabel metal2 s 108578 0 108634 800 6 o_waddr0_1[0]
port 341 nsew signal output
rlabel metal3 s 163813 17280 164613 17400 6 o_waddr0_1[1]
port 342 nsew signal output
rlabel metal3 s 163813 25304 164613 25424 6 o_waddr0_1[2]
port 343 nsew signal output
rlabel metal3 s 163813 30744 164613 30864 6 o_waddr0_1[3]
port 344 nsew signal output
rlabel metal2 s 123666 0 123722 800 6 o_waddr0_1[4]
port 345 nsew signal output
rlabel metal2 s 126426 0 126482 800 6 o_waddr0_1[5]
port 346 nsew signal output
rlabel metal3 s 163813 62976 164613 63096 6 o_waddr0_1[6]
port 347 nsew signal output
rlabel metal2 s 130198 0 130254 800 6 o_waddr0_1[7]
port 348 nsew signal output
rlabel metal3 s 163813 73720 164613 73840 6 o_waddr0_1[8]
port 349 nsew signal output
rlabel metal2 s 104806 0 104862 800 6 o_web0
port 350 nsew signal output
rlabel metal2 s 105726 0 105782 800 6 o_web0_1
port 351 nsew signal output
rlabel metal3 s 163813 9256 164613 9376 6 o_wmask0[0]
port 352 nsew signal output
rlabel metal2 s 115202 0 115258 800 6 o_wmask0[1]
port 353 nsew signal output
rlabel metal3 s 163813 28024 164613 28144 6 o_wmask0[2]
port 354 nsew signal output
rlabel metal3 s 163813 36184 164613 36304 6 o_wmask0[3]
port 355 nsew signal output
rlabel metal2 s 109498 0 109554 800 6 o_wmask0_1[0]
port 356 nsew signal output
rlabel metal2 s 114190 0 114246 800 6 o_wmask0_1[1]
port 357 nsew signal output
rlabel metal2 s 117318 165957 117374 166757 6 o_wmask0_1[2]
port 358 nsew signal output
rlabel metal2 s 120814 0 120870 800 6 o_wmask0_1[3]
port 359 nsew signal output
rlabel metal4 s 4208 2128 4528 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 34928 2128 35248 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 65648 2128 65968 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 96368 2128 96688 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 127088 2128 127408 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 157808 2128 158128 164336 6 vccd1
port 360 nsew power input
rlabel metal4 s 19568 2128 19888 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 50288 2128 50608 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 81008 2128 81328 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 111728 2128 112048 164336 6 vssd1
port 361 nsew ground input
rlabel metal4 s 142448 2128 142768 164336 6 vssd1
port 361 nsew ground input
rlabel metal2 s 478 0 534 800 6 wb_clk_i
port 362 nsew signal input
rlabel metal2 s 1398 0 1454 800 6 wb_rst_i
port 363 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 wbs_ack_o
port 364 nsew signal output
rlabel metal2 s 6090 0 6146 800 6 wbs_adr_i[0]
port 365 nsew signal input
rlabel metal2 s 38014 0 38070 800 6 wbs_adr_i[10]
port 366 nsew signal input
rlabel metal2 s 40866 0 40922 800 6 wbs_adr_i[11]
port 367 nsew signal input
rlabel metal2 s 43718 0 43774 800 6 wbs_adr_i[12]
port 368 nsew signal input
rlabel metal2 s 46478 0 46534 800 6 wbs_adr_i[13]
port 369 nsew signal input
rlabel metal2 s 49330 0 49386 800 6 wbs_adr_i[14]
port 370 nsew signal input
rlabel metal2 s 52182 0 52238 800 6 wbs_adr_i[15]
port 371 nsew signal input
rlabel metal2 s 54942 0 54998 800 6 wbs_adr_i[16]
port 372 nsew signal input
rlabel metal2 s 57794 0 57850 800 6 wbs_adr_i[17]
port 373 nsew signal input
rlabel metal2 s 60646 0 60702 800 6 wbs_adr_i[18]
port 374 nsew signal input
rlabel metal2 s 63406 0 63462 800 6 wbs_adr_i[19]
port 375 nsew signal input
rlabel metal2 s 9862 0 9918 800 6 wbs_adr_i[1]
port 376 nsew signal input
rlabel metal2 s 66258 0 66314 800 6 wbs_adr_i[20]
port 377 nsew signal input
rlabel metal2 s 69110 0 69166 800 6 wbs_adr_i[21]
port 378 nsew signal input
rlabel metal2 s 71870 0 71926 800 6 wbs_adr_i[22]
port 379 nsew signal input
rlabel metal2 s 74722 0 74778 800 6 wbs_adr_i[23]
port 380 nsew signal input
rlabel metal2 s 77574 0 77630 800 6 wbs_adr_i[24]
port 381 nsew signal input
rlabel metal2 s 80334 0 80390 800 6 wbs_adr_i[25]
port 382 nsew signal input
rlabel metal2 s 83186 0 83242 800 6 wbs_adr_i[26]
port 383 nsew signal input
rlabel metal2 s 86038 0 86094 800 6 wbs_adr_i[27]
port 384 nsew signal input
rlabel metal2 s 88798 0 88854 800 6 wbs_adr_i[28]
port 385 nsew signal input
rlabel metal2 s 91650 0 91706 800 6 wbs_adr_i[29]
port 386 nsew signal input
rlabel metal2 s 13634 0 13690 800 6 wbs_adr_i[2]
port 387 nsew signal input
rlabel metal2 s 94502 0 94558 800 6 wbs_adr_i[30]
port 388 nsew signal input
rlabel metal2 s 97262 0 97318 800 6 wbs_adr_i[31]
port 389 nsew signal input
rlabel metal2 s 17406 0 17462 800 6 wbs_adr_i[3]
port 390 nsew signal input
rlabel metal2 s 21086 0 21142 800 6 wbs_adr_i[4]
port 391 nsew signal input
rlabel metal2 s 23938 0 23994 800 6 wbs_adr_i[5]
port 392 nsew signal input
rlabel metal2 s 26790 0 26846 800 6 wbs_adr_i[6]
port 393 nsew signal input
rlabel metal2 s 29550 0 29606 800 6 wbs_adr_i[7]
port 394 nsew signal input
rlabel metal2 s 32402 0 32458 800 6 wbs_adr_i[8]
port 395 nsew signal input
rlabel metal2 s 35254 0 35310 800 6 wbs_adr_i[9]
port 396 nsew signal input
rlabel metal2 s 3238 0 3294 800 6 wbs_cyc_i
port 397 nsew signal input
rlabel metal2 s 7010 0 7066 800 6 wbs_dat_i[0]
port 398 nsew signal input
rlabel metal2 s 39026 0 39082 800 6 wbs_dat_i[10]
port 399 nsew signal input
rlabel metal2 s 41786 0 41842 800 6 wbs_dat_i[11]
port 400 nsew signal input
rlabel metal2 s 44638 0 44694 800 6 wbs_dat_i[12]
port 401 nsew signal input
rlabel metal2 s 47490 0 47546 800 6 wbs_dat_i[13]
port 402 nsew signal input
rlabel metal2 s 50250 0 50306 800 6 wbs_dat_i[14]
port 403 nsew signal input
rlabel metal2 s 53102 0 53158 800 6 wbs_dat_i[15]
port 404 nsew signal input
rlabel metal2 s 55954 0 56010 800 6 wbs_dat_i[16]
port 405 nsew signal input
rlabel metal2 s 58714 0 58770 800 6 wbs_dat_i[17]
port 406 nsew signal input
rlabel metal2 s 61566 0 61622 800 6 wbs_dat_i[18]
port 407 nsew signal input
rlabel metal2 s 64418 0 64474 800 6 wbs_dat_i[19]
port 408 nsew signal input
rlabel metal2 s 10782 0 10838 800 6 wbs_dat_i[1]
port 409 nsew signal input
rlabel metal2 s 67178 0 67234 800 6 wbs_dat_i[20]
port 410 nsew signal input
rlabel metal2 s 70030 0 70086 800 6 wbs_dat_i[21]
port 411 nsew signal input
rlabel metal2 s 72882 0 72938 800 6 wbs_dat_i[22]
port 412 nsew signal input
rlabel metal2 s 75642 0 75698 800 6 wbs_dat_i[23]
port 413 nsew signal input
rlabel metal2 s 78494 0 78550 800 6 wbs_dat_i[24]
port 414 nsew signal input
rlabel metal2 s 81346 0 81402 800 6 wbs_dat_i[25]
port 415 nsew signal input
rlabel metal2 s 84106 0 84162 800 6 wbs_dat_i[26]
port 416 nsew signal input
rlabel metal2 s 86958 0 87014 800 6 wbs_dat_i[27]
port 417 nsew signal input
rlabel metal2 s 89810 0 89866 800 6 wbs_dat_i[28]
port 418 nsew signal input
rlabel metal2 s 92570 0 92626 800 6 wbs_dat_i[29]
port 419 nsew signal input
rlabel metal2 s 14554 0 14610 800 6 wbs_dat_i[2]
port 420 nsew signal input
rlabel metal2 s 95422 0 95478 800 6 wbs_dat_i[30]
port 421 nsew signal input
rlabel metal2 s 98274 0 98330 800 6 wbs_dat_i[31]
port 422 nsew signal input
rlabel metal2 s 18326 0 18382 800 6 wbs_dat_i[3]
port 423 nsew signal input
rlabel metal2 s 22098 0 22154 800 6 wbs_dat_i[4]
port 424 nsew signal input
rlabel metal2 s 24858 0 24914 800 6 wbs_dat_i[5]
port 425 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 wbs_dat_i[6]
port 426 nsew signal input
rlabel metal2 s 30562 0 30618 800 6 wbs_dat_i[7]
port 427 nsew signal input
rlabel metal2 s 33322 0 33378 800 6 wbs_dat_i[8]
port 428 nsew signal input
rlabel metal2 s 36174 0 36230 800 6 wbs_dat_i[9]
port 429 nsew signal input
rlabel metal2 s 7930 0 7986 800 6 wbs_dat_o[0]
port 430 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 wbs_dat_o[10]
port 431 nsew signal output
rlabel metal2 s 42798 0 42854 800 6 wbs_dat_o[11]
port 432 nsew signal output
rlabel metal2 s 45558 0 45614 800 6 wbs_dat_o[12]
port 433 nsew signal output
rlabel metal2 s 48410 0 48466 800 6 wbs_dat_o[13]
port 434 nsew signal output
rlabel metal2 s 51262 0 51318 800 6 wbs_dat_o[14]
port 435 nsew signal output
rlabel metal2 s 54022 0 54078 800 6 wbs_dat_o[15]
port 436 nsew signal output
rlabel metal2 s 56874 0 56930 800 6 wbs_dat_o[16]
port 437 nsew signal output
rlabel metal2 s 59726 0 59782 800 6 wbs_dat_o[17]
port 438 nsew signal output
rlabel metal2 s 62486 0 62542 800 6 wbs_dat_o[18]
port 439 nsew signal output
rlabel metal2 s 65338 0 65394 800 6 wbs_dat_o[19]
port 440 nsew signal output
rlabel metal2 s 11702 0 11758 800 6 wbs_dat_o[1]
port 441 nsew signal output
rlabel metal2 s 68190 0 68246 800 6 wbs_dat_o[20]
port 442 nsew signal output
rlabel metal2 s 70950 0 71006 800 6 wbs_dat_o[21]
port 443 nsew signal output
rlabel metal2 s 73802 0 73858 800 6 wbs_dat_o[22]
port 444 nsew signal output
rlabel metal2 s 76654 0 76710 800 6 wbs_dat_o[23]
port 445 nsew signal output
rlabel metal2 s 79414 0 79470 800 6 wbs_dat_o[24]
port 446 nsew signal output
rlabel metal2 s 82266 0 82322 800 6 wbs_dat_o[25]
port 447 nsew signal output
rlabel metal2 s 85118 0 85174 800 6 wbs_dat_o[26]
port 448 nsew signal output
rlabel metal2 s 87878 0 87934 800 6 wbs_dat_o[27]
port 449 nsew signal output
rlabel metal2 s 90730 0 90786 800 6 wbs_dat_o[28]
port 450 nsew signal output
rlabel metal2 s 93582 0 93638 800 6 wbs_dat_o[29]
port 451 nsew signal output
rlabel metal2 s 15474 0 15530 800 6 wbs_dat_o[2]
port 452 nsew signal output
rlabel metal2 s 96342 0 96398 800 6 wbs_dat_o[30]
port 453 nsew signal output
rlabel metal2 s 99194 0 99250 800 6 wbs_dat_o[31]
port 454 nsew signal output
rlabel metal2 s 19246 0 19302 800 6 wbs_dat_o[3]
port 455 nsew signal output
rlabel metal2 s 23018 0 23074 800 6 wbs_dat_o[4]
port 456 nsew signal output
rlabel metal2 s 25870 0 25926 800 6 wbs_dat_o[5]
port 457 nsew signal output
rlabel metal2 s 28630 0 28686 800 6 wbs_dat_o[6]
port 458 nsew signal output
rlabel metal2 s 31482 0 31538 800 6 wbs_dat_o[7]
port 459 nsew signal output
rlabel metal2 s 34334 0 34390 800 6 wbs_dat_o[8]
port 460 nsew signal output
rlabel metal2 s 37094 0 37150 800 6 wbs_dat_o[9]
port 461 nsew signal output
rlabel metal2 s 8942 0 8998 800 6 wbs_sel_i[0]
port 462 nsew signal input
rlabel metal2 s 12622 0 12678 800 6 wbs_sel_i[1]
port 463 nsew signal input
rlabel metal2 s 16394 0 16450 800 6 wbs_sel_i[2]
port 464 nsew signal input
rlabel metal2 s 20166 0 20222 800 6 wbs_sel_i[3]
port 465 nsew signal input
rlabel metal2 s 4158 0 4214 800 6 wbs_stb_i
port 466 nsew signal input
rlabel metal2 s 5170 0 5226 800 6 wbs_we_i
port 467 nsew signal input
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 164613 166757
string LEFview TRUE
string GDS_FILE /project/openlane/user_proj/runs/user_proj/results/magic/user_proj.gds
string GDS_END 70415346
string GDS_START 110
<< end >>

