magic
tech sky130A
magscale 1 2
timestamp 1639150748
<< locali >>
rect 295257 700519 295291 700553
rect 295257 700485 295993 700519
rect 301513 700111 301547 700553
rect 301605 700111 301639 700689
rect 36001 697663 36035 699329
rect 65625 698343 65659 699329
rect 80161 698411 80195 699329
rect 95157 698479 95191 699329
rect 100033 698547 100067 699329
rect 109877 698683 109911 699329
rect 114569 698615 114603 699329
rect 148977 698751 149011 699329
rect 158821 698819 158855 699329
rect 163881 698887 163915 699329
rect 168849 699091 168883 699329
rect 173725 699023 173759 699329
rect 188445 699227 188479 699329
rect 379529 699295 379563 699465
rect 394157 699159 394191 699465
rect 408877 698955 408911 699465
rect 434729 697731 434763 697901
rect 434913 697527 434947 697765
rect 442365 697731 442399 697901
rect 453957 697799 453991 699465
rect 521853 697731 521887 699397
rect 442273 697663 442307 697697
rect 442273 697629 442457 697663
rect 551293 697595 551327 699397
rect 434763 697493 434947 697527
rect 7481 527 7515 697
rect 240517 595 240551 697
rect 281825 595 281859 765
rect 212123 561 212273 595
rect 224601 323 224635 493
rect 251189 391 251223 561
rect 283113 595 283147 697
rect 307677 663 307711 833
rect 280721 187 280755 561
rect 284585 323 284619 629
rect 297281 323 297315 561
rect 307953 527 307987 561
rect 307895 493 307987 527
rect 310253 255 310287 561
rect 311449 459 311483 561
rect 312645 391 312679 561
rect 315865 391 315899 629
rect 316049 527 316083 833
rect 338681 187 338715 561
rect 339877 459 339911 561
rect 340981 119 341015 561
rect 354597 527 354631 629
rect 369409 595 369443 697
rect 357817 119 357851 425
rect 367017 391 367051 561
rect 371801 595 371835 697
rect 392225 663 392259 833
rect 400321 663 400355 833
rect 405381 595 405415 1037
rect 380667 561 380817 595
rect 409245 595 409279 697
rect 360761 51 360795 221
rect 368213 51 368247 561
rect 371893 119 371927 493
rect 385969 255 386003 561
rect 413753 527 413787 1309
rect 397745 493 397837 527
rect 397745 391 397779 493
rect 416697 323 416731 697
rect 417157 595 417191 901
rect 417893 595 417927 1037
rect 418629 595 418663 765
rect 419917 595 419951 969
rect 426357 663 426391 1309
rect 427001 663 427035 969
rect 427921 663 427955 901
rect 399309 51 399343 289
rect 427277 255 427311 629
rect 428565 595 428599 697
rect 431877 663 431911 1105
rect 434453 663 434487 833
rect 438777 595 438811 1037
rect 439145 595 439179 765
rect 440157 595 440191 969
rect 441077 595 441111 969
rect 445033 663 445067 1105
rect 435557 51 435591 561
rect 449633 527 449667 1105
rect 452301 527 452335 1037
rect 452393 663 452427 765
rect 454325 731 454359 1037
rect 454417 663 454451 969
rect 455889 527 455923 901
rect 457085 663 457119 833
rect 458005 663 458039 969
rect 459201 663 459235 1037
rect 460305 663 460339 1241
rect 461961 663 461995 1105
rect 456993 51 457027 357
rect 457545 255 457579 561
rect 465549 459 465583 765
rect 466285 663 466319 901
rect 466377 663 466411 969
rect 468309 595 468343 1173
rect 471805 391 471839 969
rect 472817 663 472851 1105
rect 474565 663 474599 1241
rect 475761 595 475795 765
rect 475853 527 475887 765
rect 476773 459 476807 697
rect 479165 595 479199 1241
rect 461501 119 461535 357
rect 479533 255 479567 901
rect 480637 595 480671 901
rect 480729 391 480763 697
rect 480821 595 480855 969
rect 480913 119 480947 561
rect 481465 527 481499 833
rect 482937 119 482971 1173
rect 483765 527 483799 1037
rect 487445 663 487479 969
rect 487721 663 487755 1105
rect 489929 595 489963 765
rect 490481 595 490515 833
rect 492689 663 492723 901
rect 493333 663 493367 969
rect 494713 595 494747 1241
rect 498117 595 498151 833
rect 498945 595 498979 901
rect 499405 595 499439 1173
rect 500141 595 500175 1037
rect 502993 595 503027 1105
rect 486433 323 486467 561
rect 484961 119 484995 221
rect 493517 187 493551 561
rect 498209 119 498243 561
rect 503913 527 503947 1173
rect 504649 527 504683 1309
rect 505201 663 505235 765
rect 505753 663 505787 833
rect 507869 663 507903 1241
rect 505109 527 505143 629
rect 508605 255 508639 969
rect 508881 255 508915 697
rect 508973 323 509007 697
rect 509893 459 509927 629
rect 510353 459 510387 1105
rect 510997 459 511031 765
rect 512193 527 512227 969
rect 513757 527 513791 1173
rect 514769 391 514803 493
rect 514953 391 514987 901
rect 515413 391 515447 1037
rect 520749 663 520783 1309
rect 521853 663 521887 833
rect 524245 595 524279 1241
rect 524429 663 524463 833
rect 525073 527 525107 901
rect 526269 663 526303 765
rect 526637 595 526671 1105
rect 528845 595 528879 765
rect 529029 595 529063 969
rect 530685 731 530719 901
rect 538873 799 538907 901
rect 532985 595 533019 765
rect 540621 765 540839 799
rect 533077 663 533111 765
rect 533169 595 533203 629
rect 532985 561 533203 595
rect 540621 595 540655 765
rect 529489 323 529523 425
rect 540713 391 540747 697
rect 540805 595 540839 765
rect 540805 561 540897 595
rect 546233 527 546267 1241
rect 548901 527 548935 969
rect 550281 595 550315 765
rect 551201 595 551235 833
rect 553041 595 553075 1173
rect 555801 663 555835 1037
rect 558193 799 558227 969
rect 558745 663 558779 969
rect 529581 119 529615 289
rect 552673 119 552707 561
rect 553133 527 553167 561
rect 552983 493 553167 527
rect 553317 187 553351 357
rect 566933 51 566967 765
<< viali >>
rect 301605 700689 301639 700723
rect 295257 700553 295291 700587
rect 301513 700553 301547 700587
rect 295993 700485 296027 700519
rect 301513 700077 301547 700111
rect 301605 700077 301639 700111
rect 379529 699465 379563 699499
rect 36001 699329 36035 699363
rect 65625 699329 65659 699363
rect 80161 699329 80195 699363
rect 95157 699329 95191 699363
rect 100033 699329 100067 699363
rect 109877 699329 109911 699363
rect 109877 698649 109911 698683
rect 114569 699329 114603 699363
rect 148977 699329 149011 699363
rect 158821 699329 158855 699363
rect 163881 699329 163915 699363
rect 168849 699329 168883 699363
rect 168849 699057 168883 699091
rect 173725 699329 173759 699363
rect 188445 699329 188479 699363
rect 379529 699261 379563 699295
rect 394157 699465 394191 699499
rect 188445 699193 188479 699227
rect 394157 699125 394191 699159
rect 408877 699465 408911 699499
rect 173725 698989 173759 699023
rect 408877 698921 408911 698955
rect 453957 699465 453991 699499
rect 163881 698853 163915 698887
rect 158821 698785 158855 698819
rect 148977 698717 149011 698751
rect 114569 698581 114603 698615
rect 100033 698513 100067 698547
rect 95157 698445 95191 698479
rect 80161 698377 80195 698411
rect 65625 698309 65659 698343
rect 434729 697901 434763 697935
rect 442365 697901 442399 697935
rect 434729 697697 434763 697731
rect 434913 697765 434947 697799
rect 36001 697629 36035 697663
rect 453957 697765 453991 697799
rect 521853 699397 521887 699431
rect 442273 697697 442307 697731
rect 442365 697697 442399 697731
rect 521853 697697 521887 697731
rect 551293 699397 551327 699431
rect 442457 697629 442491 697663
rect 551293 697561 551327 697595
rect 434729 697493 434763 697527
rect 413753 1309 413787 1343
rect 405381 1037 405415 1071
rect 307677 833 307711 867
rect 281825 765 281859 799
rect 7481 697 7515 731
rect 240517 697 240551 731
rect 212089 561 212123 595
rect 212273 561 212307 595
rect 240517 561 240551 595
rect 251189 561 251223 595
rect 7481 493 7515 527
rect 224601 493 224635 527
rect 251189 357 251223 391
rect 280721 561 280755 595
rect 281825 561 281859 595
rect 283113 697 283147 731
rect 316049 833 316083 867
rect 283113 561 283147 595
rect 284585 629 284619 663
rect 307677 629 307711 663
rect 315865 629 315899 663
rect 224601 289 224635 323
rect 284585 289 284619 323
rect 297281 561 297315 595
rect 307953 561 307987 595
rect 307861 493 307895 527
rect 310253 561 310287 595
rect 297281 289 297315 323
rect 311449 561 311483 595
rect 311449 425 311483 459
rect 312645 561 312679 595
rect 312645 357 312679 391
rect 392225 833 392259 867
rect 369409 697 369443 731
rect 354597 629 354631 663
rect 316049 493 316083 527
rect 338681 561 338715 595
rect 315865 357 315899 391
rect 310253 221 310287 255
rect 280721 153 280755 187
rect 339877 561 339911 595
rect 339877 425 339911 459
rect 340981 561 341015 595
rect 338681 153 338715 187
rect 354597 493 354631 527
rect 367017 561 367051 595
rect 340981 85 341015 119
rect 357817 425 357851 459
rect 367017 357 367051 391
rect 368213 561 368247 595
rect 369409 561 369443 595
rect 371801 697 371835 731
rect 392225 629 392259 663
rect 400321 833 400355 867
rect 400321 629 400355 663
rect 371801 561 371835 595
rect 380633 561 380667 595
rect 380817 561 380851 595
rect 385969 561 386003 595
rect 405381 561 405415 595
rect 409245 697 409279 731
rect 409245 561 409279 595
rect 357817 85 357851 119
rect 360761 221 360795 255
rect 360761 17 360795 51
rect 371893 493 371927 527
rect 426357 1309 426391 1343
rect 417893 1037 417927 1071
rect 417157 901 417191 935
rect 397837 493 397871 527
rect 413753 493 413787 527
rect 416697 697 416731 731
rect 397745 357 397779 391
rect 417157 561 417191 595
rect 419917 969 419951 1003
rect 417893 561 417927 595
rect 418629 765 418663 799
rect 418629 561 418663 595
rect 504649 1309 504683 1343
rect 460305 1241 460339 1275
rect 431877 1105 431911 1139
rect 426357 629 426391 663
rect 427001 969 427035 1003
rect 427921 901 427955 935
rect 427001 629 427035 663
rect 427277 629 427311 663
rect 427921 629 427955 663
rect 428565 697 428599 731
rect 419917 561 419951 595
rect 385969 221 386003 255
rect 399309 289 399343 323
rect 416697 289 416731 323
rect 371893 85 371927 119
rect 368213 17 368247 51
rect 445033 1105 445067 1139
rect 438777 1037 438811 1071
rect 431877 629 431911 663
rect 434453 833 434487 867
rect 434453 629 434487 663
rect 440157 969 440191 1003
rect 428565 561 428599 595
rect 435557 561 435591 595
rect 438777 561 438811 595
rect 439145 765 439179 799
rect 439145 561 439179 595
rect 440157 561 440191 595
rect 441077 969 441111 1003
rect 445033 629 445067 663
rect 449633 1105 449667 1139
rect 441077 561 441111 595
rect 427277 221 427311 255
rect 399309 17 399343 51
rect 449633 493 449667 527
rect 452301 1037 452335 1071
rect 454325 1037 454359 1071
rect 452393 765 452427 799
rect 459201 1037 459235 1071
rect 454325 697 454359 731
rect 454417 969 454451 1003
rect 452393 629 452427 663
rect 458005 969 458039 1003
rect 454417 629 454451 663
rect 455889 901 455923 935
rect 452301 493 452335 527
rect 457085 833 457119 867
rect 457085 629 457119 663
rect 458005 629 458039 663
rect 459201 629 459235 663
rect 474565 1241 474599 1275
rect 468309 1173 468343 1207
rect 460305 629 460339 663
rect 461961 1105 461995 1139
rect 466377 969 466411 1003
rect 466285 901 466319 935
rect 461961 629 461995 663
rect 465549 765 465583 799
rect 455889 493 455923 527
rect 457545 561 457579 595
rect 435557 17 435591 51
rect 456993 357 457027 391
rect 466285 629 466319 663
rect 466377 629 466411 663
rect 472817 1105 472851 1139
rect 468309 561 468343 595
rect 471805 969 471839 1003
rect 465549 425 465583 459
rect 472817 629 472851 663
rect 479165 1241 479199 1275
rect 474565 629 474599 663
rect 475761 765 475795 799
rect 475761 561 475795 595
rect 475853 765 475887 799
rect 475853 493 475887 527
rect 476773 697 476807 731
rect 494713 1241 494747 1275
rect 482937 1173 482971 1207
rect 480821 969 480855 1003
rect 479165 561 479199 595
rect 479533 901 479567 935
rect 476773 425 476807 459
rect 457545 221 457579 255
rect 461501 357 461535 391
rect 471805 357 471839 391
rect 480637 901 480671 935
rect 480637 561 480671 595
rect 480729 697 480763 731
rect 481465 833 481499 867
rect 480821 561 480855 595
rect 480913 561 480947 595
rect 480729 357 480763 391
rect 479533 221 479567 255
rect 461501 85 461535 119
rect 481465 493 481499 527
rect 480913 85 480947 119
rect 487721 1105 487755 1139
rect 483765 1037 483799 1071
rect 487445 969 487479 1003
rect 487445 629 487479 663
rect 493333 969 493367 1003
rect 492689 901 492723 935
rect 490481 833 490515 867
rect 487721 629 487755 663
rect 489929 765 489963 799
rect 483765 493 483799 527
rect 486433 561 486467 595
rect 489929 561 489963 595
rect 492689 629 492723 663
rect 493333 629 493367 663
rect 499405 1173 499439 1207
rect 498945 901 498979 935
rect 490481 561 490515 595
rect 493517 561 493551 595
rect 494713 561 494747 595
rect 498117 833 498151 867
rect 498117 561 498151 595
rect 498209 561 498243 595
rect 498945 561 498979 595
rect 503913 1173 503947 1207
rect 502993 1105 503027 1139
rect 499405 561 499439 595
rect 500141 1037 500175 1071
rect 500141 561 500175 595
rect 502993 561 503027 595
rect 486433 289 486467 323
rect 482937 85 482971 119
rect 484961 221 484995 255
rect 493517 153 493551 187
rect 484961 85 484995 119
rect 503913 493 503947 527
rect 520749 1309 520783 1343
rect 507869 1241 507903 1275
rect 505753 833 505787 867
rect 505201 765 505235 799
rect 504649 493 504683 527
rect 505109 629 505143 663
rect 505201 629 505235 663
rect 505753 629 505787 663
rect 513757 1173 513791 1207
rect 510353 1105 510387 1139
rect 507869 629 507903 663
rect 508605 969 508639 1003
rect 505109 493 505143 527
rect 508605 221 508639 255
rect 508881 697 508915 731
rect 508973 697 509007 731
rect 509893 629 509927 663
rect 509893 425 509927 459
rect 512193 969 512227 1003
rect 510353 425 510387 459
rect 510997 765 511031 799
rect 512193 493 512227 527
rect 515413 1037 515447 1071
rect 514953 901 514987 935
rect 513757 493 513791 527
rect 514769 493 514803 527
rect 510997 425 511031 459
rect 514769 357 514803 391
rect 514953 357 514987 391
rect 524245 1241 524279 1275
rect 520749 629 520783 663
rect 521853 833 521887 867
rect 521853 629 521887 663
rect 546233 1241 546267 1275
rect 526637 1105 526671 1139
rect 525073 901 525107 935
rect 524429 833 524463 867
rect 524429 629 524463 663
rect 524245 561 524279 595
rect 526269 765 526303 799
rect 526269 629 526303 663
rect 529029 969 529063 1003
rect 526637 561 526671 595
rect 528845 765 528879 799
rect 528845 561 528879 595
rect 530685 901 530719 935
rect 538873 901 538907 935
rect 530685 697 530719 731
rect 532985 765 533019 799
rect 529029 561 529063 595
rect 533077 765 533111 799
rect 538873 765 538907 799
rect 533077 629 533111 663
rect 533169 629 533203 663
rect 540621 561 540655 595
rect 540713 697 540747 731
rect 525073 493 525107 527
rect 515413 357 515447 391
rect 529489 425 529523 459
rect 508973 289 509007 323
rect 540897 561 540931 595
rect 553041 1173 553075 1207
rect 546233 493 546267 527
rect 548901 969 548935 1003
rect 551201 833 551235 867
rect 550281 765 550315 799
rect 550281 561 550315 595
rect 555801 1037 555835 1071
rect 558193 969 558227 1003
rect 558193 765 558227 799
rect 558745 969 558779 1003
rect 555801 629 555835 663
rect 558745 629 558779 663
rect 566933 765 566967 799
rect 551201 561 551235 595
rect 552673 561 552707 595
rect 553041 561 553075 595
rect 553133 561 553167 595
rect 548901 493 548935 527
rect 540713 357 540747 391
rect 529489 289 529523 323
rect 529581 289 529615 323
rect 508881 221 508915 255
rect 498209 85 498243 119
rect 529581 85 529615 119
rect 552949 493 552983 527
rect 553317 357 553351 391
rect 553317 153 553351 187
rect 552673 85 552707 119
rect 456993 17 457027 51
rect 566933 17 566967 51
<< metal1 >>
rect 235442 703808 235448 703860
rect 235500 703848 235506 703860
rect 300854 703848 300860 703860
rect 235500 703820 300860 703848
rect 235500 703808 235506 703820
rect 300854 703808 300860 703820
rect 300912 703808 300918 703860
rect 271782 703740 271788 703792
rect 271840 703780 271846 703792
rect 364702 703780 364708 703792
rect 271840 703752 364708 703780
rect 271840 703740 271846 703752
rect 364702 703740 364708 703752
rect 364760 703740 364766 703792
rect 257246 703672 257252 703724
rect 257304 703712 257310 703724
rect 429470 703712 429476 703724
rect 257304 703684 429476 703712
rect 257304 703672 257310 703684
rect 429470 703672 429476 703684
rect 429528 703672 429534 703724
rect 242434 703604 242440 703656
rect 242492 703644 242498 703656
rect 430022 703644 430028 703656
rect 242492 703616 430028 703644
rect 242492 703604 242498 703616
rect 430022 703604 430028 703616
rect 430080 703604 430086 703656
rect 170490 703536 170496 703588
rect 170548 703576 170554 703588
rect 315482 703576 315488 703588
rect 170548 703548 315488 703576
rect 170548 703536 170554 703548
rect 315482 703536 315488 703548
rect 315540 703536 315546 703588
rect 227622 703468 227628 703520
rect 227680 703508 227686 703520
rect 464430 703508 464436 703520
rect 227680 703480 464436 703508
rect 227680 703468 227686 703480
rect 464430 703468 464436 703480
rect 464488 703468 464494 703520
rect 105446 703400 105452 703452
rect 105504 703440 105510 703452
rect 330294 703440 330300 703452
rect 105504 703412 330300 703440
rect 105504 703400 105510 703412
rect 330294 703400 330300 703412
rect 330352 703400 330358 703452
rect 40494 703332 40500 703384
rect 40552 703372 40558 703384
rect 345014 703372 345020 703384
rect 40552 703344 345020 703372
rect 40552 703332 40558 703344
rect 345014 703332 345020 703344
rect 345072 703332 345078 703384
rect 1486 703264 1492 703316
rect 1544 703304 1550 703316
rect 359734 703304 359740 703316
rect 1544 703276 359740 703304
rect 1544 703264 1550 703276
rect 359734 703264 359740 703276
rect 359792 703264 359798 703316
rect 212994 703196 213000 703248
rect 213052 703236 213058 703248
rect 576394 703236 576400 703248
rect 213052 703208 576400 703236
rect 213052 703196 213058 703208
rect 576394 703196 576400 703208
rect 576452 703196 576458 703248
rect 1578 703128 1584 703180
rect 1636 703168 1642 703180
rect 374454 703168 374460 703180
rect 1636 703140 374460 703168
rect 1636 703128 1642 703140
rect 374454 703128 374460 703140
rect 374512 703128 374518 703180
rect 198274 703060 198280 703112
rect 198332 703100 198338 703112
rect 575014 703100 575020 703112
rect 198332 703072 575020 703100
rect 198332 703060 198338 703072
rect 575014 703060 575020 703072
rect 575072 703060 575078 703112
rect 1670 702992 1676 703044
rect 1728 703032 1734 703044
rect 389174 703032 389180 703044
rect 1728 703004 389180 703032
rect 1728 702992 1734 703004
rect 389174 702992 389180 703004
rect 389232 702992 389238 703044
rect 183370 702924 183376 702976
rect 183428 702964 183434 702976
rect 573634 702964 573640 702976
rect 183428 702936 573640 702964
rect 183428 702924 183434 702936
rect 573634 702924 573640 702936
rect 573692 702924 573698 702976
rect 1762 702856 1768 702908
rect 1820 702896 1826 702908
rect 403894 702896 403900 702908
rect 1820 702868 403900 702896
rect 1820 702856 1826 702868
rect 403894 702856 403900 702868
rect 403952 702856 403958 702908
rect 139302 702788 139308 702840
rect 139360 702828 139366 702840
rect 578970 702828 578976 702840
rect 139360 702800 578976 702828
rect 139360 702788 139366 702800
rect 578970 702788 578976 702800
rect 579028 702788 579034 702840
rect 2590 702720 2596 702772
rect 2648 702760 2654 702772
rect 448146 702760 448152 702772
rect 2648 702732 448152 702760
rect 2648 702720 2654 702732
rect 448146 702720 448152 702732
rect 448204 702720 448210 702772
rect 2222 702652 2228 702704
rect 2280 702692 2286 702704
rect 477586 702692 477592 702704
rect 2280 702664 477592 702692
rect 2280 702652 2286 702664
rect 477586 702652 477592 702664
rect 477644 702652 477650 702704
rect 198 702584 204 702636
rect 256 702624 262 702636
rect 507118 702624 507124 702636
rect 256 702596 507124 702624
rect 256 702584 262 702596
rect 507118 702584 507124 702596
rect 507176 702584 507182 702636
rect 14 702516 20 702568
rect 72 702556 78 702568
rect 536834 702556 536840 702568
rect 72 702528 536840 702556
rect 72 702516 78 702528
rect 536834 702516 536840 702528
rect 536892 702516 536898 702568
rect 21450 702448 21456 702500
rect 21508 702488 21514 702500
rect 576118 702488 576124 702500
rect 21508 702460 576124 702488
rect 21508 702448 21514 702460
rect 576118 702448 576124 702460
rect 576176 702448 576182 702500
rect 85298 702380 85304 702432
rect 85356 702420 85362 702432
rect 569402 702420 569408 702432
rect 85356 702392 569408 702420
rect 85356 702380 85362 702392
rect 569402 702380 569408 702392
rect 569460 702380 569466 702432
rect 247402 702312 247408 702364
rect 247460 702352 247466 702364
rect 299382 702352 299388 702364
rect 247460 702324 299388 702352
rect 247460 702312 247466 702324
rect 299382 702312 299388 702324
rect 299440 702312 299446 702364
rect 217870 702244 217876 702296
rect 217928 702284 217934 702296
rect 313366 702284 313372 702296
rect 217928 702256 313372 702284
rect 217928 702244 217934 702256
rect 313366 702244 313372 702256
rect 313424 702244 313430 702296
rect 154022 702176 154028 702228
rect 154080 702216 154086 702228
rect 292574 702216 292580 702228
rect 154080 702188 292580 702216
rect 154080 702176 154086 702188
rect 292574 702176 292580 702188
rect 292632 702176 292638 702228
rect 299106 702176 299112 702228
rect 299164 702216 299170 702228
rect 320450 702216 320456 702228
rect 299164 702188 320456 702216
rect 299164 702176 299170 702188
rect 320450 702176 320456 702188
rect 320508 702176 320514 702228
rect 178586 702108 178592 702160
rect 178644 702148 178650 702160
rect 329190 702148 329196 702160
rect 178644 702120 329196 702148
rect 178644 702108 178650 702120
rect 329190 702108 329196 702120
rect 329248 702108 329254 702160
rect 329742 702108 329748 702160
rect 329800 702148 329806 702160
rect 349890 702148 349896 702160
rect 329800 702120 349896 702148
rect 329800 702108 329806 702120
rect 349890 702108 349896 702120
rect 349948 702108 349954 702160
rect 75454 702040 75460 702092
rect 75512 702080 75518 702092
rect 266446 702080 266452 702092
rect 75512 702052 266452 702080
rect 75512 702040 75518 702052
rect 266446 702040 266452 702052
rect 266504 702040 266510 702092
rect 304994 702040 305000 702092
rect 305052 702080 305058 702092
rect 438302 702080 438308 702092
rect 305052 702052 438308 702080
rect 305052 702040 305058 702052
rect 438302 702040 438308 702052
rect 438360 702040 438366 702092
rect 90174 701972 90180 702024
rect 90232 702012 90238 702024
rect 343634 702012 343640 702024
rect 90232 701984 343640 702012
rect 90232 701972 90238 701984
rect 343634 701972 343640 701984
rect 343692 701972 343698 702024
rect 349062 701972 349068 702024
rect 349120 702012 349126 702024
rect 467834 702012 467840 702024
rect 349120 701984 467840 702012
rect 349120 701972 349126 701984
rect 467834 701972 467840 701984
rect 467892 701972 467898 702024
rect 192938 701904 192944 701956
rect 192996 701944 193002 701956
rect 577590 701944 577596 701956
rect 192996 701916 577596 701944
rect 192996 701904 193002 701916
rect 577590 701904 577596 701916
rect 577648 701904 577654 701956
rect 4430 701836 4436 701888
rect 4488 701876 4494 701888
rect 414198 701876 414204 701888
rect 4488 701848 414204 701876
rect 4488 701836 4494 701848
rect 414198 701836 414204 701848
rect 414256 701836 414262 701888
rect 1946 701768 1952 701820
rect 2004 701808 2010 701820
rect 423674 701808 423680 701820
rect 2004 701780 423680 701808
rect 2004 701768 2010 701780
rect 423674 701768 423680 701780
rect 423732 701768 423738 701820
rect 144270 701700 144276 701752
rect 144328 701740 144334 701752
rect 572162 701740 572168 701752
rect 144328 701712 572168 701740
rect 144328 701700 144334 701712
rect 572162 701700 572168 701712
rect 572220 701700 572226 701752
rect 134426 701632 134432 701684
rect 134484 701672 134490 701684
rect 578878 701672 578884 701684
rect 134484 701644 578884 701672
rect 134484 701632 134490 701644
rect 578878 701632 578884 701644
rect 578936 701632 578942 701684
rect 129458 701564 129464 701616
rect 129516 701604 129522 701616
rect 573450 701604 573456 701616
rect 129516 701576 573456 701604
rect 129516 701564 129522 701576
rect 573450 701564 573456 701576
rect 573508 701564 573514 701616
rect 566 701496 572 701548
rect 624 701536 630 701548
rect 453022 701536 453028 701548
rect 624 701508 453028 701536
rect 624 701496 630 701508
rect 453022 701496 453028 701508
rect 453080 701496 453086 701548
rect 119706 701428 119712 701480
rect 119764 701468 119770 701480
rect 574830 701468 574836 701480
rect 119764 701440 574836 701468
rect 119764 701428 119770 701440
rect 574830 701428 574836 701440
rect 574888 701428 574894 701480
rect 658 701360 664 701412
rect 716 701400 722 701412
rect 458174 701400 458180 701412
rect 716 701372 458180 701400
rect 716 701360 722 701372
rect 458174 701360 458180 701372
rect 458232 701360 458238 701412
rect 2406 701292 2412 701344
rect 2464 701332 2470 701344
rect 472710 701332 472716 701344
rect 2464 701304 472716 701332
rect 2464 701292 2470 701304
rect 472710 701292 472716 701304
rect 472768 701292 472774 701344
rect 104802 701224 104808 701276
rect 104860 701264 104866 701276
rect 577498 701264 577504 701276
rect 104860 701236 577504 701264
rect 104860 701224 104866 701236
rect 577498 701224 577504 701236
rect 577556 701224 577562 701276
rect 474 701156 480 701208
rect 532 701196 538 701208
rect 482554 701196 482560 701208
rect 532 701168 482560 701196
rect 532 701156 538 701168
rect 482554 701156 482560 701168
rect 482612 701156 482618 701208
rect 4338 701088 4344 701140
rect 4396 701128 4402 701140
rect 487430 701128 487436 701140
rect 4396 701100 487436 701128
rect 4396 701088 4402 701100
rect 487430 701088 487436 701100
rect 487488 701088 487494 701140
rect 556890 701088 556896 701140
rect 556948 701128 556954 701140
rect 564434 701128 564440 701140
rect 556948 701100 564440 701128
rect 556948 701088 556954 701100
rect 564434 701088 564440 701100
rect 564492 701088 564498 701140
rect 281258 701020 281264 701072
rect 281316 701060 281322 701072
rect 305730 701060 305736 701072
rect 281316 701032 305736 701060
rect 281316 701020 281322 701032
rect 305730 701020 305736 701032
rect 305788 701020 305794 701072
rect 313274 701020 313280 701072
rect 313332 701060 313338 701072
rect 335354 701060 335360 701072
rect 313332 701032 335360 701060
rect 313332 701020 313338 701032
rect 335354 701020 335360 701032
rect 335412 701020 335418 701072
rect 424962 701020 424968 701072
rect 425020 701060 425026 701072
rect 443270 701060 443276 701072
rect 425020 701032 443276 701060
rect 425020 701020 425026 701032
rect 443270 701020 443276 701032
rect 443328 701020 443334 701072
rect 8110 700952 8116 701004
rect 8168 700992 8174 701004
rect 329742 700992 329748 701004
rect 8168 700964 329748 700992
rect 8168 700952 8174 700964
rect 329742 700952 329748 700964
rect 329800 700952 329806 701004
rect 464430 700952 464436 701004
rect 464488 700992 464494 701004
rect 559650 700992 559656 701004
rect 464488 700964 559656 700992
rect 464488 700952 464494 700964
rect 559650 700952 559656 700964
rect 559708 700952 559714 701004
rect 72970 700884 72976 700936
rect 73028 700924 73034 700936
rect 313274 700924 313280 700936
rect 73028 700896 313280 700924
rect 73028 700884 73034 700896
rect 313274 700884 313280 700896
rect 313332 700884 313338 700936
rect 252278 700816 252284 700868
rect 252336 700856 252342 700868
rect 478506 700856 478512 700868
rect 252336 700828 478512 700856
rect 252336 700816 252342 700828
rect 478506 700816 478512 700828
rect 478564 700816 478570 700868
rect 89162 700748 89168 700800
rect 89220 700788 89226 700800
rect 340046 700788 340052 700800
rect 89220 700760 340052 700788
rect 89220 700748 89226 700760
rect 340046 700748 340052 700760
rect 340104 700748 340110 700800
rect 343634 700748 343640 700800
rect 343692 700788 343698 700800
rect 580534 700788 580540 700800
rect 343692 700760 580540 700788
rect 343692 700748 343698 700760
rect 580534 700748 580540 700760
rect 580592 700748 580598 700800
rect 137830 700680 137836 700732
rect 137888 700720 137894 700732
rect 299106 700720 299112 700732
rect 137888 700692 299112 700720
rect 137888 700680 137894 700692
rect 299106 700680 299112 700692
rect 299164 700680 299170 700732
rect 299382 700680 299388 700732
rect 299440 700720 299446 700732
rect 301593 700723 301651 700729
rect 301593 700720 301605 700723
rect 299440 700692 301605 700720
rect 299440 700680 299446 700692
rect 301593 700689 301605 700692
rect 301639 700689 301651 700723
rect 301593 700683 301651 700689
rect 329190 700680 329196 700732
rect 329248 700720 329254 700732
rect 580718 700720 580724 700732
rect 329248 700692 580724 700720
rect 329248 700680 329254 700692
rect 580718 700680 580724 700692
rect 580776 700680 580782 700732
rect 154114 700612 154120 700664
rect 154172 700652 154178 700664
rect 325326 700652 325332 700664
rect 154172 700624 325332 700652
rect 154172 700612 154178 700624
rect 325326 700612 325332 700624
rect 325384 700612 325390 700664
rect 326062 700612 326068 700664
rect 326120 700652 326126 700664
rect 580442 700652 580448 700664
rect 326120 700624 580448 700652
rect 326120 700612 326126 700624
rect 580442 700612 580448 700624
rect 580500 700612 580506 700664
rect 3602 700544 3608 700596
rect 3660 700584 3666 700596
rect 260834 700584 260840 700596
rect 3660 700556 260840 700584
rect 3660 700544 3666 700556
rect 260834 700544 260840 700556
rect 260892 700544 260898 700596
rect 267642 700544 267648 700596
rect 267700 700584 267706 700596
rect 291378 700584 291384 700596
rect 267700 700556 291384 700584
rect 267700 700544 267706 700556
rect 291378 700544 291384 700556
rect 291436 700544 291442 700596
rect 292574 700544 292580 700596
rect 292632 700584 292638 700596
rect 295245 700587 295303 700593
rect 295245 700584 295257 700587
rect 292632 700556 295257 700584
rect 292632 700544 292638 700556
rect 295245 700553 295257 700556
rect 295291 700553 295303 700587
rect 295245 700547 295303 700553
rect 295334 700544 295340 700596
rect 295392 700584 295398 700596
rect 300118 700584 300124 700596
rect 295392 700556 300124 700584
rect 295392 700544 295398 700556
rect 300118 700544 300124 700556
rect 300176 700544 300182 700596
rect 301501 700587 301559 700593
rect 301501 700553 301513 700587
rect 301547 700584 301559 700587
rect 310606 700584 310612 700596
rect 301547 700556 310612 700584
rect 301547 700553 301559 700556
rect 301501 700547 301559 700553
rect 310606 700544 310612 700556
rect 310664 700544 310670 700596
rect 313366 700544 313372 700596
rect 313424 700584 313430 700596
rect 580074 700584 580080 700596
rect 313424 700556 580080 700584
rect 313424 700544 313430 700556
rect 580074 700544 580080 700556
rect 580132 700544 580138 700596
rect 3694 700476 3700 700528
rect 3752 700516 3758 700528
rect 266354 700516 266360 700528
rect 3752 700488 266360 700516
rect 3752 700476 3758 700488
rect 266354 700476 266360 700488
rect 266412 700476 266418 700528
rect 283834 700476 283840 700528
rect 283892 700516 283898 700528
rect 295886 700516 295892 700528
rect 283892 700488 295892 700516
rect 283892 700476 283898 700488
rect 295886 700476 295892 700488
rect 295944 700476 295950 700528
rect 295981 700519 296039 700525
rect 295981 700485 295993 700519
rect 296027 700516 296039 700519
rect 580626 700516 580632 700528
rect 296027 700488 580632 700516
rect 296027 700485 296039 700488
rect 295981 700479 296039 700485
rect 580626 700476 580632 700488
rect 580684 700476 580690 700528
rect 232682 700408 232688 700460
rect 232740 700448 232746 700460
rect 527174 700448 527180 700460
rect 232740 700420 527180 700448
rect 232740 700408 232746 700420
rect 527174 700408 527180 700420
rect 527232 700408 527238 700460
rect 237098 700340 237104 700392
rect 237156 700380 237162 700392
rect 543458 700380 543464 700392
rect 237156 700352 543464 700380
rect 237156 700340 237162 700352
rect 543458 700340 543464 700352
rect 543516 700340 543522 700392
rect 24302 700272 24308 700324
rect 24360 700312 24366 700324
rect 354950 700312 354956 700324
rect 24360 700284 354956 700312
rect 24360 700272 24366 700284
rect 354950 700272 354956 700284
rect 355008 700272 355014 700324
rect 430022 700272 430028 700324
rect 430080 700312 430086 700324
rect 494790 700312 494796 700324
rect 430080 700284 494796 700312
rect 430080 700272 430086 700284
rect 494790 700272 494796 700284
rect 494848 700272 494854 700324
rect 266998 700204 267004 700256
rect 267056 700244 267062 700256
rect 413646 700244 413652 700256
rect 267056 700216 413652 700244
rect 267056 700204 267062 700216
rect 413646 700204 413652 700216
rect 413704 700204 413710 700256
rect 261800 700136 261806 700188
rect 261858 700176 261864 700188
rect 397454 700176 397460 700188
rect 261858 700148 397460 700176
rect 261858 700136 261864 700148
rect 397454 700136 397460 700148
rect 397512 700136 397518 700188
rect 202782 700068 202788 700120
rect 202840 700068 202846 700120
rect 218974 700068 218980 700120
rect 219032 700108 219038 700120
rect 301501 700111 301559 700117
rect 301501 700108 301513 700111
rect 219032 700080 301513 700108
rect 219032 700068 219038 700080
rect 301501 700077 301513 700080
rect 301547 700077 301559 700111
rect 301501 700071 301559 700077
rect 301593 700111 301651 700117
rect 301593 700077 301605 700111
rect 301639 700108 301651 700111
rect 462314 700108 462320 700120
rect 301639 700080 462320 700108
rect 301639 700077 301651 700080
rect 301593 700071 301651 700077
rect 462314 700068 462320 700080
rect 462372 700068 462378 700120
rect 202800 700040 202828 700068
rect 281258 700040 281264 700052
rect 202800 700012 281264 700040
rect 281258 700000 281264 700012
rect 281316 700000 281322 700052
rect 281350 700000 281356 700052
rect 281408 700040 281414 700052
rect 348786 700040 348792 700052
rect 281408 700012 348792 700040
rect 281408 700000 281414 700012
rect 348786 700000 348792 700012
rect 348844 700000 348850 700052
rect 276842 699932 276848 699984
rect 276900 699972 276906 699984
rect 332502 699972 332508 699984
rect 276900 699944 332508 699972
rect 276900 699932 276906 699944
rect 332502 699932 332508 699944
rect 332560 699932 332566 699984
rect 222838 699864 222844 699916
rect 222896 699904 222902 699916
rect 577682 699904 577688 699916
rect 222896 699876 577688 699904
rect 222896 699864 222902 699876
rect 577682 699864 577688 699876
rect 577740 699864 577746 699916
rect 4246 699796 4252 699848
rect 4304 699836 4310 699848
rect 364610 699836 364616 699848
rect 4304 699808 364616 699836
rect 4304 699796 4310 699808
rect 364610 699796 364616 699808
rect 364668 699796 364674 699848
rect 208118 699728 208124 699780
rect 208176 699768 208182 699780
rect 570874 699768 570880 699780
rect 208176 699740 570880 699768
rect 208176 699728 208182 699740
rect 570874 699728 570880 699740
rect 570932 699728 570938 699780
rect 2958 699660 2964 699712
rect 3016 699700 3022 699712
rect 369762 699700 369768 699712
rect 3016 699672 369768 699700
rect 3016 699660 3022 699672
rect 369762 699660 369768 699672
rect 369820 699660 369826 699712
rect 3326 699592 3332 699644
rect 3384 699632 3390 699644
rect 304994 699632 305000 699644
rect 3384 699604 305000 699632
rect 3384 699592 3390 699604
rect 304994 699592 305000 699604
rect 305052 699592 305058 699644
rect 266446 699524 266452 699576
rect 266504 699564 266510 699576
rect 580350 699564 580356 699576
rect 266504 699536 580356 699564
rect 266504 699524 266510 699536
rect 580350 699524 580356 699536
rect 580408 699524 580414 699576
rect 3970 699456 3976 699508
rect 4028 699496 4034 699508
rect 349062 699496 349068 699508
rect 4028 699468 349068 699496
rect 4028 699456 4034 699468
rect 349062 699456 349068 699468
rect 349120 699456 349126 699508
rect 379514 699496 379520 699508
rect 379475 699468 379520 699496
rect 379514 699456 379520 699468
rect 379572 699456 379578 699508
rect 394142 699496 394148 699508
rect 394103 699468 394148 699496
rect 394142 699456 394148 699468
rect 394200 699456 394206 699508
rect 408862 699496 408868 699508
rect 408823 699468 408868 699496
rect 408862 699456 408868 699468
rect 408920 699456 408926 699508
rect 453942 699496 453948 699508
rect 453903 699468 453948 699496
rect 453942 699456 453948 699468
rect 454000 699456 454006 699508
rect 3234 699388 3240 699440
rect 3292 699428 3298 699440
rect 424962 699428 424968 699440
rect 3292 699400 424968 699428
rect 3292 699388 3298 699400
rect 424962 699388 424968 699400
rect 425020 699388 425026 699440
rect 521838 699428 521844 699440
rect 521799 699400 521844 699428
rect 521838 699388 521844 699400
rect 521896 699388 521902 699440
rect 551278 699428 551284 699440
rect 551239 699400 551284 699428
rect 551278 699388 551284 699400
rect 551336 699388 551342 699440
rect 35986 699360 35992 699372
rect 35947 699332 35992 699360
rect 35986 699320 35992 699332
rect 36044 699320 36050 699372
rect 65610 699360 65616 699372
rect 65571 699332 65616 699360
rect 65610 699320 65616 699332
rect 65668 699320 65674 699372
rect 80146 699360 80152 699372
rect 80107 699332 80152 699360
rect 80146 699320 80152 699332
rect 80204 699320 80210 699372
rect 95142 699360 95148 699372
rect 95103 699332 95148 699360
rect 95142 699320 95148 699332
rect 95200 699320 95206 699372
rect 100018 699360 100024 699372
rect 99979 699332 100024 699360
rect 100018 699320 100024 699332
rect 100076 699320 100082 699372
rect 109862 699360 109868 699372
rect 109823 699332 109868 699360
rect 109862 699320 109868 699332
rect 109920 699320 109926 699372
rect 114554 699360 114560 699372
rect 114515 699332 114560 699360
rect 114554 699320 114560 699332
rect 114612 699320 114618 699372
rect 148962 699360 148968 699372
rect 148923 699332 148968 699360
rect 148962 699320 148968 699332
rect 149020 699320 149026 699372
rect 158806 699360 158812 699372
rect 158767 699332 158812 699360
rect 158806 699320 158812 699332
rect 158864 699320 158870 699372
rect 163866 699360 163872 699372
rect 163827 699332 163872 699360
rect 163866 699320 163872 699332
rect 163924 699320 163930 699372
rect 168834 699360 168840 699372
rect 168795 699332 168840 699360
rect 168834 699320 168840 699332
rect 168892 699320 168898 699372
rect 173710 699360 173716 699372
rect 173671 699332 173716 699360
rect 173710 699320 173716 699332
rect 173768 699320 173774 699372
rect 188430 699360 188436 699372
rect 188391 699332 188436 699360
rect 188430 699320 188436 699332
rect 188488 699320 188494 699372
rect 202966 699320 202972 699372
rect 203024 699360 203030 699372
rect 572254 699360 572260 699372
rect 203024 699332 572260 699360
rect 203024 699320 203030 699332
rect 572254 699320 572260 699332
rect 572312 699320 572318 699372
rect 934 699252 940 699304
rect 992 699292 998 699304
rect 379517 699295 379575 699301
rect 379517 699292 379529 699295
rect 992 699264 379529 699292
rect 992 699252 998 699264
rect 379517 699261 379529 699264
rect 379563 699261 379575 699295
rect 379517 699255 379575 699261
rect 188433 699227 188491 699233
rect 188433 699193 188445 699227
rect 188479 699224 188491 699227
rect 569586 699224 569592 699236
rect 188479 699196 569592 699224
rect 188479 699193 188491 699196
rect 188433 699187 188491 699193
rect 569586 699184 569592 699196
rect 569644 699184 569650 699236
rect 842 699116 848 699168
rect 900 699156 906 699168
rect 394145 699159 394203 699165
rect 394145 699156 394157 699159
rect 900 699128 394157 699156
rect 900 699116 906 699128
rect 394145 699125 394157 699128
rect 394191 699125 394203 699159
rect 394145 699119 394203 699125
rect 168837 699091 168895 699097
rect 168837 699057 168849 699091
rect 168883 699088 168895 699091
rect 565354 699088 565360 699100
rect 168883 699060 565360 699088
rect 168883 699057 168895 699060
rect 168837 699051 168895 699057
rect 565354 699048 565360 699060
rect 565412 699048 565418 699100
rect 173713 699023 173771 699029
rect 173713 698989 173725 699023
rect 173759 699020 173771 699023
rect 573542 699020 573548 699032
rect 173759 698992 573548 699020
rect 173759 698989 173771 698992
rect 173713 698983 173771 698989
rect 573542 698980 573548 698992
rect 573600 698980 573606 699032
rect 750 698912 756 698964
rect 808 698952 814 698964
rect 408865 698955 408923 698961
rect 408865 698952 408877 698955
rect 808 698924 408877 698952
rect 808 698912 814 698924
rect 408865 698921 408877 698924
rect 408911 698921 408923 698955
rect 408865 698915 408923 698921
rect 163869 698887 163927 698893
rect 163869 698853 163881 698887
rect 163915 698884 163927 698887
rect 576302 698884 576308 698896
rect 163915 698856 576308 698884
rect 163915 698853 163927 698856
rect 163869 698847 163927 698853
rect 576302 698844 576308 698856
rect 576360 698844 576366 698896
rect 158809 698819 158867 698825
rect 158809 698785 158821 698819
rect 158855 698816 158867 698819
rect 570782 698816 570788 698828
rect 158855 698788 570788 698816
rect 158855 698785 158867 698788
rect 158809 698779 158867 698785
rect 570782 698776 570788 698788
rect 570840 698776 570846 698828
rect 148965 698751 149023 698757
rect 148965 698717 148977 698751
rect 149011 698748 149023 698751
rect 576210 698748 576216 698760
rect 149011 698720 576216 698748
rect 149011 698717 149023 698720
rect 148965 698711 149023 698717
rect 576210 698708 576216 698720
rect 576268 698708 576274 698760
rect 109865 698683 109923 698689
rect 109865 698649 109877 698683
rect 109911 698680 109923 698683
rect 569494 698680 569500 698692
rect 109911 698652 569500 698680
rect 109911 698649 109923 698652
rect 109865 698643 109923 698649
rect 569494 698640 569500 698652
rect 569552 698640 569558 698692
rect 114557 698615 114615 698621
rect 114557 698581 114569 698615
rect 114603 698612 114615 698615
rect 574922 698612 574928 698624
rect 114603 698584 574928 698612
rect 114603 698581 114615 698584
rect 114557 698575 114615 698581
rect 574922 698572 574928 698584
rect 574980 698572 574986 698624
rect 100021 698547 100079 698553
rect 100021 698513 100033 698547
rect 100067 698544 100079 698547
rect 570690 698544 570696 698556
rect 100067 698516 570696 698544
rect 100067 698513 100079 698516
rect 100021 698507 100079 698513
rect 570690 698504 570696 698516
rect 570748 698504 570754 698556
rect 95145 698479 95203 698485
rect 95145 698445 95157 698479
rect 95191 698476 95203 698479
rect 565262 698476 565268 698488
rect 95191 698448 565268 698476
rect 95191 698445 95203 698448
rect 95145 698439 95203 698445
rect 565262 698436 565268 698448
rect 565320 698436 565326 698488
rect 80149 698411 80207 698417
rect 80149 698377 80161 698411
rect 80195 698408 80207 698411
rect 566734 698408 566740 698420
rect 80195 698380 566740 698408
rect 80195 698377 80207 698380
rect 80149 698371 80207 698377
rect 566734 698368 566740 698380
rect 566792 698368 566798 698420
rect 65613 698343 65671 698349
rect 65613 698309 65625 698343
rect 65659 698340 65671 698343
rect 566550 698340 566556 698352
rect 65659 698312 566556 698340
rect 65659 698309 65671 698312
rect 65613 698303 65671 698309
rect 566550 698300 566556 698312
rect 566608 698300 566614 698352
rect 434717 697935 434775 697941
rect 434717 697901 434729 697935
rect 434763 697932 434775 697935
rect 442353 697935 442411 697941
rect 442353 697932 442365 697935
rect 434763 697904 442365 697932
rect 434763 697901 434775 697904
rect 434717 697895 434775 697901
rect 442353 697901 442365 697904
rect 442399 697901 442411 697935
rect 442353 697895 442411 697901
rect 434901 697799 434959 697805
rect 434901 697765 434913 697799
rect 434947 697796 434959 697799
rect 453945 697799 454003 697805
rect 453945 697796 453957 697799
rect 434947 697768 453957 697796
rect 434947 697765 434959 697768
rect 434901 697759 434959 697765
rect 453945 697765 453957 697768
rect 453991 697765 454003 697799
rect 453945 697759 454003 697765
rect 106 697688 112 697740
rect 164 697728 170 697740
rect 434717 697731 434775 697737
rect 434717 697728 434729 697731
rect 164 697700 434729 697728
rect 164 697688 170 697700
rect 434717 697697 434729 697700
rect 434763 697697 434775 697731
rect 442261 697731 442319 697737
rect 442261 697728 442273 697731
rect 434717 697691 434775 697697
rect 434824 697700 442273 697728
rect 35989 697663 36047 697669
rect 35989 697629 36001 697663
rect 36035 697660 36047 697663
rect 434824 697660 434852 697700
rect 442261 697697 442273 697700
rect 442307 697697 442319 697731
rect 442261 697691 442319 697697
rect 442353 697731 442411 697737
rect 442353 697697 442365 697731
rect 442399 697728 442411 697731
rect 521841 697731 521899 697737
rect 521841 697728 521853 697731
rect 442399 697700 521853 697728
rect 442399 697697 442411 697700
rect 442353 697691 442411 697697
rect 521841 697697 521853 697700
rect 521887 697697 521899 697731
rect 521841 697691 521899 697697
rect 36035 697632 434852 697660
rect 442445 697663 442503 697669
rect 36035 697629 36047 697632
rect 35989 697623 36047 697629
rect 442445 697629 442457 697663
rect 442491 697660 442503 697663
rect 574738 697660 574744 697672
rect 442491 697632 574744 697660
rect 442491 697629 442503 697632
rect 442445 697623 442503 697629
rect 574738 697620 574744 697632
rect 574796 697620 574802 697672
rect 2038 697552 2044 697604
rect 2096 697592 2102 697604
rect 551281 697595 551339 697601
rect 551281 697592 551293 697595
rect 2096 697564 439544 697592
rect 2096 697552 2102 697564
rect 3418 697484 3424 697536
rect 3476 697524 3482 697536
rect 434717 697527 434775 697533
rect 434717 697524 434729 697527
rect 3476 697496 434729 697524
rect 3476 697484 3482 697496
rect 434717 697493 434729 697496
rect 434763 697493 434775 697527
rect 439516 697524 439544 697564
rect 444346 697564 551293 697592
rect 444346 697524 444374 697564
rect 551281 697561 551293 697564
rect 551327 697561 551339 697595
rect 551281 697555 551339 697561
rect 439516 697496 444374 697524
rect 434717 697487 434775 697493
rect 577682 684428 577688 684480
rect 577740 684468 577746 684480
rect 580810 684468 580816 684480
rect 577740 684440 580816 684468
rect 577740 684428 577746 684440
rect 580810 684428 580816 684440
rect 580868 684428 580874 684480
rect 576394 671984 576400 672036
rect 576452 672024 576458 672036
rect 579614 672024 579620 672036
rect 576452 671996 579620 672024
rect 576452 671984 576458 671996
rect 579614 671984 579620 671996
rect 579672 671984 579678 672036
rect 572254 644376 572260 644428
rect 572312 644416 572318 644428
rect 580166 644416 580172 644428
rect 572312 644388 580172 644416
rect 572312 644376 572318 644388
rect 580166 644376 580172 644388
rect 580224 644376 580230 644428
rect 570874 632000 570880 632052
rect 570932 632040 570938 632052
rect 580166 632040 580172 632052
rect 570932 632012 580172 632040
rect 570932 632000 570938 632012
rect 580166 632000 580172 632012
rect 580224 632000 580230 632052
rect 575014 618196 575020 618248
rect 575072 618236 575078 618248
rect 580166 618236 580172 618248
rect 575072 618208 580172 618236
rect 575072 618196 575078 618208
rect 580166 618196 580172 618208
rect 580224 618196 580230 618248
rect 569586 591948 569592 592000
rect 569644 591988 569650 592000
rect 580166 591988 580172 592000
rect 569644 591960 580172 591988
rect 569644 591948 569650 591960
rect 580166 591948 580172 591960
rect 580224 591948 580230 592000
rect 577590 578144 577596 578196
rect 577648 578184 577654 578196
rect 580810 578184 580816 578196
rect 577648 578156 580816 578184
rect 577648 578144 577654 578156
rect 580810 578144 580816 578156
rect 580868 578144 580874 578196
rect 573634 564340 573640 564392
rect 573692 564380 573698 564392
rect 580166 564380 580172 564392
rect 573692 564352 580172 564380
rect 573692 564340 573698 564352
rect 580166 564340 580172 564352
rect 580224 564340 580230 564392
rect 573542 538160 573548 538212
rect 573600 538200 573606 538212
rect 580166 538200 580172 538212
rect 573600 538172 580172 538200
rect 573600 538160 573606 538172
rect 580166 538160 580172 538172
rect 580224 538160 580230 538212
rect 2774 514836 2780 514888
rect 2832 514876 2838 514888
rect 4430 514876 4436 514888
rect 2832 514848 4436 514876
rect 2832 514836 2838 514848
rect 4430 514836 4436 514848
rect 4488 514836 4494 514888
rect 565354 511912 565360 511964
rect 565412 511952 565418 511964
rect 580166 511952 580172 511964
rect 565412 511924 580172 511952
rect 565412 511912 565418 511924
rect 580166 511912 580172 511924
rect 580224 511912 580230 511964
rect 570782 485732 570788 485784
rect 570840 485772 570846 485784
rect 579614 485772 579620 485784
rect 570840 485744 579620 485772
rect 570840 485732 570846 485744
rect 579614 485732 579620 485744
rect 579672 485732 579678 485784
rect 576302 471928 576308 471980
rect 576360 471968 576366 471980
rect 579798 471968 579804 471980
rect 576360 471940 579804 471968
rect 576360 471928 576366 471940
rect 579798 471928 579804 471940
rect 579856 471928 579862 471980
rect 572162 431876 572168 431928
rect 572220 431916 572226 431928
rect 579706 431916 579712 431928
rect 572220 431888 579712 431916
rect 572220 431876 572226 431888
rect 579706 431876 579712 431888
rect 579764 431876 579770 431928
rect 576210 419432 576216 419484
rect 576268 419472 576274 419484
rect 580166 419472 580172 419484
rect 576268 419444 580172 419472
rect 576268 419432 576274 419444
rect 580166 419432 580172 419444
rect 580224 419432 580230 419484
rect 573450 379448 573456 379500
rect 573508 379488 573514 379500
rect 579614 379488 579620 379500
rect 573508 379460 579620 379488
rect 573508 379448 573514 379460
rect 579614 379448 579620 379460
rect 579672 379448 579678 379500
rect 572070 353200 572076 353252
rect 572128 353240 572134 353252
rect 580166 353240 580172 353252
rect 572128 353212 580172 353240
rect 572128 353200 572134 353212
rect 580166 353200 580172 353212
rect 580224 353200 580230 353252
rect 574922 325592 574928 325644
rect 574980 325632 574986 325644
rect 580166 325632 580172 325644
rect 574980 325604 580172 325632
rect 574980 325592 574986 325604
rect 580166 325592 580172 325604
rect 580224 325592 580230 325644
rect 574830 313216 574836 313268
rect 574888 313256 574894 313268
rect 580166 313256 580172 313268
rect 574888 313228 580172 313256
rect 574888 313216 574894 313228
rect 580166 313216 580172 313228
rect 580224 313216 580230 313268
rect 569494 299412 569500 299464
rect 569552 299452 569558 299464
rect 580166 299452 580172 299464
rect 569552 299424 580172 299452
rect 569552 299412 569558 299424
rect 580166 299412 580172 299424
rect 580224 299412 580230 299464
rect 570690 273164 570696 273216
rect 570748 273204 570754 273216
rect 579614 273204 579620 273216
rect 570748 273176 579620 273204
rect 570748 273164 570754 273176
rect 579614 273164 579620 273176
rect 579672 273164 579678 273216
rect 577498 259360 577504 259412
rect 577556 259400 577562 259412
rect 580626 259400 580632 259412
rect 577556 259372 580632 259400
rect 577556 259360 577562 259372
rect 580626 259360 580632 259372
rect 580684 259360 580690 259412
rect 565262 245556 565268 245608
rect 565320 245596 565326 245608
rect 580166 245596 580172 245608
rect 565320 245568 580172 245596
rect 565320 245556 565326 245568
rect 580166 245556 580172 245568
rect 580224 245556 580230 245608
rect 569402 233180 569408 233232
rect 569460 233220 569466 233232
rect 579982 233220 579988 233232
rect 569460 233192 579988 233220
rect 569460 233180 569466 233192
rect 579982 233180 579988 233192
rect 580040 233180 580046 233232
rect 566734 206932 566740 206984
rect 566792 206972 566798 206984
rect 580166 206972 580172 206984
rect 566792 206944 580172 206972
rect 566792 206932 566798 206944
rect 580166 206932 580172 206944
rect 580224 206932 580230 206984
rect 566550 166948 566556 167000
rect 566608 166988 566614 167000
rect 580166 166988 580172 167000
rect 566608 166960 580172 166988
rect 566608 166948 566614 166960
rect 580166 166948 580172 166960
rect 580224 166948 580230 167000
rect 569310 153144 569316 153196
rect 569368 153184 569374 153196
rect 579798 153184 579804 153196
rect 569368 153156 579804 153184
rect 569368 153144 569374 153156
rect 579798 153144 579804 153156
rect 579856 153144 579862 153196
rect 573358 139340 573364 139392
rect 573416 139380 573422 139392
rect 580166 139380 580172 139392
rect 573416 139352 580172 139380
rect 573416 139340 573422 139352
rect 580166 139340 580172 139352
rect 580224 139340 580230 139392
rect 565170 126896 565176 126948
rect 565228 126936 565234 126948
rect 580166 126936 580172 126948
rect 565228 126908 580172 126936
rect 565228 126896 565234 126908
rect 580166 126896 580172 126908
rect 580224 126896 580230 126948
rect 566642 113092 566648 113144
rect 566700 113132 566706 113144
rect 580166 113132 580172 113144
rect 566700 113104 580172 113132
rect 566700 113092 566706 113104
rect 580166 113092 580172 113104
rect 580224 113092 580230 113144
rect 571978 100648 571984 100700
rect 572036 100688 572042 100700
rect 580166 100688 580172 100700
rect 572036 100660 580172 100688
rect 572036 100648 572042 100660
rect 580166 100648 580172 100660
rect 580224 100648 580230 100700
rect 574738 86912 574744 86964
rect 574796 86952 574802 86964
rect 580166 86952 580172 86964
rect 574796 86924 580172 86952
rect 574796 86912 574802 86924
rect 580166 86912 580172 86924
rect 580224 86912 580230 86964
rect 565078 73108 565084 73160
rect 565136 73148 565142 73160
rect 579982 73148 579988 73160
rect 565136 73120 579988 73148
rect 565136 73108 565142 73120
rect 579982 73108 579988 73120
rect 580040 73108 580046 73160
rect 570598 60664 570604 60716
rect 570656 60704 570662 60716
rect 580166 60704 580172 60716
rect 570656 60676 580172 60704
rect 570656 60664 570662 60676
rect 580166 60664 580172 60676
rect 580224 60664 580230 60716
rect 576118 46860 576124 46912
rect 576176 46900 576182 46912
rect 580166 46900 580172 46912
rect 576176 46872 580172 46900
rect 576176 46860 576182 46872
rect 580166 46860 580172 46872
rect 580224 46860 580230 46912
rect 566458 33056 566464 33108
rect 566516 33096 566522 33108
rect 580166 33096 580172 33108
rect 566516 33068 580172 33096
rect 566516 33056 566522 33068
rect 580166 33056 580172 33068
rect 580224 33056 580230 33108
rect 569218 20612 569224 20664
rect 569276 20652 569282 20664
rect 580166 20652 580172 20664
rect 569276 20624 580172 20652
rect 569276 20612 569282 20624
rect 580166 20612 580172 20624
rect 580224 20612 580230 20664
rect 569126 3068 569132 3120
rect 569184 3108 569190 3120
rect 577406 3108 577412 3120
rect 569184 3080 577412 3108
rect 569184 3068 569190 3080
rect 577406 3068 577412 3080
rect 577464 3068 577470 3120
rect 563698 3000 563704 3052
rect 563756 3040 563762 3052
rect 583386 3040 583392 3052
rect 563756 3012 583392 3040
rect 563756 3000 563762 3012
rect 583386 3000 583392 3012
rect 583444 3000 583450 3052
rect 563514 2932 563520 2984
rect 563572 2972 563578 2984
rect 573910 2972 573916 2984
rect 563572 2944 573916 2972
rect 563572 2932 563578 2944
rect 573910 2932 573916 2944
rect 573968 2932 573974 2984
rect 563790 2864 563796 2916
rect 563848 2904 563854 2916
rect 563848 2876 567194 2904
rect 563848 2864 563854 2876
rect 567166 2836 567194 2876
rect 575474 2864 575480 2916
rect 575532 2904 575538 2916
rect 582190 2904 582196 2916
rect 575532 2876 582196 2904
rect 575532 2864 575538 2876
rect 582190 2864 582196 2876
rect 582248 2864 582254 2916
rect 576302 2836 576308 2848
rect 567166 2808 576308 2836
rect 576302 2796 576308 2808
rect 576360 2796 576366 2848
rect 2958 2048 2964 2100
rect 3016 2088 3022 2100
rect 564434 2088 564440 2100
rect 3016 2060 564440 2088
rect 3016 2048 3022 2060
rect 564434 2048 564440 2060
rect 564492 2048 564498 2100
rect 565814 1368 565820 1420
rect 565872 1408 565878 1420
rect 569034 1408 569040 1420
rect 565872 1380 569040 1408
rect 565872 1368 565878 1380
rect 569034 1368 569040 1380
rect 569092 1368 569098 1420
rect 413741 1343 413799 1349
rect 413741 1309 413753 1343
rect 413787 1340 413799 1343
rect 426345 1343 426403 1349
rect 426345 1340 426357 1343
rect 413787 1312 426357 1340
rect 413787 1309 413799 1312
rect 413741 1303 413799 1309
rect 426345 1309 426357 1312
rect 426391 1309 426403 1343
rect 426345 1303 426403 1309
rect 504637 1343 504695 1349
rect 504637 1309 504649 1343
rect 504683 1340 504695 1343
rect 520737 1343 520795 1349
rect 520737 1340 520749 1343
rect 504683 1312 520749 1340
rect 504683 1309 504695 1312
rect 504637 1303 504695 1309
rect 520737 1309 520749 1312
rect 520783 1309 520795 1343
rect 520737 1303 520795 1309
rect 460293 1275 460351 1281
rect 460293 1241 460305 1275
rect 460339 1272 460351 1275
rect 474553 1275 474611 1281
rect 474553 1272 474565 1275
rect 460339 1244 474565 1272
rect 460339 1241 460351 1244
rect 460293 1235 460351 1241
rect 474553 1241 474565 1244
rect 474599 1241 474611 1275
rect 474553 1235 474611 1241
rect 479153 1275 479211 1281
rect 479153 1241 479165 1275
rect 479199 1272 479211 1275
rect 494701 1275 494759 1281
rect 494701 1272 494713 1275
rect 479199 1244 494713 1272
rect 479199 1241 479211 1244
rect 479153 1235 479211 1241
rect 494701 1241 494713 1244
rect 494747 1241 494759 1275
rect 494701 1235 494759 1241
rect 507857 1275 507915 1281
rect 507857 1241 507869 1275
rect 507903 1272 507915 1275
rect 524233 1275 524291 1281
rect 524233 1272 524245 1275
rect 507903 1244 524245 1272
rect 507903 1241 507915 1244
rect 507857 1235 507915 1241
rect 524233 1241 524245 1244
rect 524279 1241 524291 1275
rect 524233 1235 524291 1241
rect 546221 1275 546279 1281
rect 546221 1241 546233 1275
rect 546267 1272 546279 1275
rect 564434 1272 564440 1284
rect 546267 1244 564440 1272
rect 546267 1241 546279 1244
rect 546221 1235 546279 1241
rect 564434 1232 564440 1244
rect 564492 1232 564498 1284
rect 468297 1207 468355 1213
rect 468297 1173 468309 1207
rect 468343 1204 468355 1207
rect 482925 1207 482983 1213
rect 482925 1204 482937 1207
rect 468343 1176 482937 1204
rect 468343 1173 468355 1176
rect 468297 1167 468355 1173
rect 482925 1173 482937 1176
rect 482971 1173 482983 1207
rect 499393 1207 499451 1213
rect 499393 1204 499405 1207
rect 482925 1167 482983 1173
rect 490576 1176 499405 1204
rect 431865 1139 431923 1145
rect 431865 1105 431877 1139
rect 431911 1136 431923 1139
rect 445021 1139 445079 1145
rect 445021 1136 445033 1139
rect 431911 1108 445033 1136
rect 431911 1105 431923 1108
rect 431865 1099 431923 1105
rect 445021 1105 445033 1108
rect 445067 1105 445079 1139
rect 445021 1099 445079 1105
rect 449621 1139 449679 1145
rect 449621 1105 449633 1139
rect 449667 1136 449679 1139
rect 461949 1139 462007 1145
rect 461949 1136 461961 1139
rect 449667 1108 461961 1136
rect 449667 1105 449679 1108
rect 449621 1099 449679 1105
rect 461949 1105 461961 1108
rect 461995 1105 462007 1139
rect 461949 1099 462007 1105
rect 472805 1139 472863 1145
rect 472805 1105 472817 1139
rect 472851 1136 472863 1139
rect 487709 1139 487767 1145
rect 487709 1136 487721 1139
rect 472851 1108 487721 1136
rect 472851 1105 472863 1108
rect 472805 1099 472863 1105
rect 487709 1105 487721 1108
rect 487755 1105 487767 1139
rect 487709 1099 487767 1105
rect 405369 1071 405427 1077
rect 405369 1037 405381 1071
rect 405415 1068 405427 1071
rect 417881 1071 417939 1077
rect 417881 1068 417893 1071
rect 405415 1040 417893 1068
rect 405415 1037 405427 1040
rect 405369 1031 405427 1037
rect 417881 1037 417893 1040
rect 417927 1037 417939 1071
rect 417881 1031 417939 1037
rect 438765 1071 438823 1077
rect 438765 1037 438777 1071
rect 438811 1068 438823 1071
rect 452289 1071 452347 1077
rect 452289 1068 452301 1071
rect 438811 1040 452301 1068
rect 438811 1037 438823 1040
rect 438765 1031 438823 1037
rect 452289 1037 452301 1040
rect 452335 1037 452347 1071
rect 452289 1031 452347 1037
rect 454313 1071 454371 1077
rect 454313 1037 454325 1071
rect 454359 1068 454371 1071
rect 459189 1071 459247 1077
rect 459189 1068 459201 1071
rect 454359 1040 459201 1068
rect 454359 1037 454371 1040
rect 454313 1031 454371 1037
rect 459189 1037 459201 1040
rect 459235 1037 459247 1071
rect 459189 1031 459247 1037
rect 483753 1071 483811 1077
rect 483753 1037 483765 1071
rect 483799 1068 483811 1071
rect 490576 1068 490604 1176
rect 499393 1173 499405 1176
rect 499439 1173 499451 1207
rect 499393 1167 499451 1173
rect 503901 1207 503959 1213
rect 503901 1173 503913 1207
rect 503947 1204 503959 1207
rect 513745 1207 513803 1213
rect 513745 1204 513757 1207
rect 503947 1176 513757 1204
rect 503947 1173 503959 1176
rect 503901 1167 503959 1173
rect 513745 1173 513757 1176
rect 513791 1173 513803 1207
rect 513745 1167 513803 1173
rect 553029 1207 553087 1213
rect 553029 1173 553041 1207
rect 553075 1204 553087 1207
rect 571518 1204 571524 1216
rect 553075 1176 571524 1204
rect 553075 1173 553087 1176
rect 553029 1167 553087 1173
rect 571518 1164 571524 1176
rect 571576 1164 571582 1216
rect 502981 1139 503039 1145
rect 502981 1136 502993 1139
rect 483799 1040 490604 1068
rect 490668 1108 502993 1136
rect 483799 1037 483811 1040
rect 483753 1031 483811 1037
rect 419905 1003 419963 1009
rect 419905 1000 419917 1003
rect 408466 972 419917 1000
rect 307665 867 307723 873
rect 307665 833 307677 867
rect 307711 864 307723 867
rect 316037 867 316095 873
rect 316037 864 316049 867
rect 307711 836 316049 864
rect 307711 833 307723 836
rect 307665 827 307723 833
rect 316037 833 316049 836
rect 316083 833 316095 867
rect 316037 827 316095 833
rect 392213 867 392271 873
rect 392213 833 392225 867
rect 392259 864 392271 867
rect 400309 867 400367 873
rect 400309 864 400321 867
rect 392259 836 400321 864
rect 392259 833 392271 836
rect 392213 827 392271 833
rect 400309 833 400321 836
rect 400355 833 400367 867
rect 400309 827 400367 833
rect 281813 799 281871 805
rect 281813 765 281825 799
rect 281859 796 281871 799
rect 281859 768 288388 796
rect 281859 765 281871 768
rect 281813 759 281871 765
rect 7469 731 7527 737
rect 7469 697 7481 731
rect 7515 728 7527 731
rect 240505 731 240563 737
rect 240505 728 240517 731
rect 7515 700 11560 728
rect 7515 697 7527 700
rect 7469 691 7527 697
rect 11532 672 11560 700
rect 237346 700 240517 728
rect 1670 620 1676 672
rect 1728 660 1734 672
rect 5350 660 5356 672
rect 1728 632 5356 660
rect 1728 620 1734 632
rect 5350 620 5356 632
rect 5408 620 5414 672
rect 6454 620 6460 672
rect 6512 660 6518 672
rect 10042 660 10048 672
rect 6512 632 10048 660
rect 6512 620 6518 632
rect 10042 620 10048 632
rect 10100 620 10106 672
rect 10152 632 11468 660
rect 566 552 572 604
rect 624 592 630 604
rect 4338 592 4344 604
rect 624 564 4344 592
rect 624 552 630 564
rect 4338 552 4344 564
rect 4396 552 4402 604
rect 5258 552 5264 604
rect 5316 592 5322 604
rect 8846 592 8852 604
rect 5316 564 8852 592
rect 5316 552 5322 564
rect 8846 552 8852 564
rect 8904 552 8910 604
rect 7466 524 7472 536
rect 7427 496 7472 524
rect 7466 484 7472 496
rect 7524 484 7530 536
rect 8570 484 8576 536
rect 8628 524 8634 536
rect 10152 524 10180 632
rect 11146 552 11152 604
rect 11204 552 11210 604
rect 11440 592 11468 632
rect 11514 620 11520 672
rect 11572 620 11578 672
rect 12618 660 12624 672
rect 11716 632 12624 660
rect 11716 592 11744 632
rect 12618 620 12624 632
rect 12676 620 12682 672
rect 13354 620 13360 672
rect 13412 660 13418 672
rect 16666 660 16672 672
rect 13412 632 16672 660
rect 13412 620 13418 632
rect 16666 620 16672 632
rect 16724 620 16730 672
rect 20622 620 20628 672
rect 20680 660 20686 672
rect 23474 660 23480 672
rect 20680 632 23480 660
rect 20680 620 20686 632
rect 23474 620 23480 632
rect 23532 620 23538 672
rect 25774 660 25780 672
rect 23584 632 25780 660
rect 11440 564 11744 592
rect 12342 552 12348 604
rect 12400 592 12406 604
rect 15562 592 15568 604
rect 12400 564 15568 592
rect 12400 552 12406 564
rect 15562 552 15568 564
rect 15620 552 15626 604
rect 19426 552 19432 604
rect 19484 592 19490 604
rect 22370 592 22376 604
rect 19484 564 22376 592
rect 19484 552 19490 564
rect 22370 552 22376 564
rect 22428 552 22434 604
rect 23014 552 23020 604
rect 23072 592 23078 604
rect 23584 592 23612 632
rect 25774 620 25780 632
rect 25832 620 25838 672
rect 28810 620 28816 672
rect 28868 660 28874 672
rect 31662 660 31668 672
rect 28868 632 31668 660
rect 28868 620 28874 632
rect 31662 620 31668 632
rect 31720 620 31726 672
rect 34790 620 34796 672
rect 34848 660 34854 672
rect 37274 660 37280 672
rect 34848 632 37280 660
rect 34848 620 34854 632
rect 37274 620 37280 632
rect 37332 620 37338 672
rect 38378 620 38384 672
rect 38436 660 38442 672
rect 38436 632 39804 660
rect 38436 620 38442 632
rect 24854 592 24860 604
rect 23072 564 23612 592
rect 23072 552 23078 564
rect 24826 552 24860 592
rect 24912 552 24918 604
rect 25314 552 25320 604
rect 25372 592 25378 604
rect 28074 592 28080 604
rect 25372 564 28080 592
rect 25372 552 25378 564
rect 28074 552 28080 564
rect 28132 552 28138 604
rect 28718 552 28724 604
rect 28776 592 28782 604
rect 29178 592 29184 604
rect 28776 564 29184 592
rect 28776 552 28782 564
rect 29178 552 29184 564
rect 29236 552 29242 604
rect 30098 552 30104 604
rect 30156 592 30162 604
rect 32582 592 32588 604
rect 30156 564 32588 592
rect 30156 552 30162 564
rect 32582 552 32588 564
rect 32640 552 32646 604
rect 37182 552 37188 604
rect 37240 552 37246 604
rect 39574 552 39580 604
rect 39632 552 39638 604
rect 39776 592 39804 632
rect 40678 620 40684 672
rect 40736 660 40742 672
rect 42794 660 42800 672
rect 40736 632 42800 660
rect 40736 620 40742 632
rect 42794 620 42800 632
rect 42852 620 42858 672
rect 46658 620 46664 672
rect 46716 660 46722 672
rect 48498 660 48504 672
rect 46716 632 48504 660
rect 46716 620 46722 632
rect 48498 620 48504 632
rect 48556 620 48562 672
rect 48958 620 48964 672
rect 49016 660 49022 672
rect 50798 660 50804 672
rect 49016 632 50804 660
rect 49016 620 49022 632
rect 50798 620 50804 632
rect 50856 620 50862 672
rect 63218 620 63224 672
rect 63276 660 63282 672
rect 63276 632 63494 660
rect 63276 620 63282 632
rect 40770 592 40776 604
rect 39776 564 40776 592
rect 40770 552 40776 564
rect 40828 552 40834 604
rect 41874 552 41880 604
rect 41932 592 41938 604
rect 43990 592 43996 604
rect 41932 564 43996 592
rect 41932 552 41938 564
rect 43990 552 43996 564
rect 44048 552 44054 604
rect 47854 552 47860 604
rect 47912 592 47918 604
rect 49602 592 49608 604
rect 47912 564 49608 592
rect 47912 552 47918 564
rect 49602 552 49608 564
rect 49660 552 49666 604
rect 50154 552 50160 604
rect 50212 552 50218 604
rect 51350 552 51356 604
rect 51408 592 51414 604
rect 53006 592 53012 604
rect 51408 564 53012 592
rect 51408 552 51414 564
rect 53006 552 53012 564
rect 53064 552 53070 604
rect 54938 552 54944 604
rect 54996 592 55002 604
rect 56410 592 56416 604
rect 54996 564 56416 592
rect 54996 552 55002 564
rect 56410 552 56416 564
rect 56468 552 56474 604
rect 62022 552 62028 604
rect 62080 592 62086 604
rect 63310 592 63316 604
rect 62080 564 63316 592
rect 62080 552 62086 564
rect 63310 552 63316 564
rect 63368 552 63374 604
rect 63466 592 63494 632
rect 64322 620 64328 672
rect 64380 660 64386 672
rect 65610 660 65616 672
rect 64380 632 65616 660
rect 64380 620 64386 632
rect 65610 620 65616 632
rect 65668 620 65674 672
rect 66714 620 66720 672
rect 66772 660 66778 672
rect 68002 660 68008 672
rect 66772 632 68008 660
rect 66772 620 66778 632
rect 68002 620 68008 632
rect 68060 620 68066 672
rect 69106 620 69112 672
rect 69164 660 69170 672
rect 70578 660 70584 672
rect 69164 632 70584 660
rect 69164 620 69170 632
rect 70578 620 70584 632
rect 70636 620 70642 672
rect 133230 620 133236 672
rect 133288 660 133294 672
rect 134150 660 134156 672
rect 133288 632 134156 660
rect 133288 620 133294 632
rect 134150 620 134156 632
rect 134208 620 134214 672
rect 136174 620 136180 672
rect 136232 660 136238 672
rect 137646 660 137652 672
rect 136232 632 137652 660
rect 136232 620 136238 632
rect 137646 620 137652 632
rect 137704 620 137710 672
rect 138750 620 138756 672
rect 138808 660 138814 672
rect 140038 660 140044 672
rect 138808 632 140044 660
rect 138808 620 138814 632
rect 140038 620 140044 632
rect 140096 620 140102 672
rect 151354 620 151360 672
rect 151412 660 151418 672
rect 153010 660 153016 672
rect 151412 632 153016 660
rect 151412 620 151418 632
rect 153010 620 153016 632
rect 153068 620 153074 672
rect 153654 620 153660 672
rect 153712 660 153718 672
rect 155402 660 155408 672
rect 153712 632 155408 660
rect 153712 620 153718 632
rect 155402 620 155408 632
rect 155460 620 155466 672
rect 162762 620 162768 672
rect 162820 660 162826 672
rect 164878 660 164884 672
rect 162820 632 164884 660
rect 162820 620 162826 632
rect 164878 620 164884 632
rect 164936 620 164942 672
rect 166074 660 166080 672
rect 165908 632 166080 660
rect 64414 592 64420 604
rect 63466 564 64420 592
rect 64414 552 64420 564
rect 64472 552 64478 604
rect 65518 552 65524 604
rect 65576 592 65582 604
rect 66806 592 66812 604
rect 65576 564 66812 592
rect 65576 552 65582 564
rect 66806 552 66812 564
rect 66864 552 66870 604
rect 70302 552 70308 604
rect 70360 592 70366 604
rect 71222 592 71228 604
rect 70360 564 71228 592
rect 70360 552 70366 564
rect 71222 552 71228 564
rect 71280 552 71286 604
rect 76190 552 76196 604
rect 76248 592 76254 604
rect 76926 592 76932 604
rect 76248 564 76932 592
rect 76248 552 76254 564
rect 76926 552 76932 564
rect 76984 552 76990 604
rect 77386 552 77392 604
rect 77444 592 77450 604
rect 78030 592 78036 604
rect 77444 564 78036 592
rect 77444 552 77450 564
rect 78030 552 78036 564
rect 78088 552 78094 604
rect 78582 552 78588 604
rect 78640 592 78646 604
rect 79134 592 79140 604
rect 78640 564 79140 592
rect 78640 552 78646 564
rect 79134 552 79140 564
rect 79192 552 79198 604
rect 79686 552 79692 604
rect 79744 592 79750 604
rect 80330 592 80336 604
rect 79744 564 80336 592
rect 79744 552 79750 564
rect 80330 552 80336 564
rect 80388 552 80394 604
rect 80882 552 80888 604
rect 80940 592 80946 604
rect 81434 592 81440 604
rect 80940 564 81440 592
rect 80940 552 80946 564
rect 81434 552 81440 564
rect 81492 552 81498 604
rect 82078 552 82084 604
rect 82136 592 82142 604
rect 82722 592 82728 604
rect 82136 564 82728 592
rect 82136 552 82142 564
rect 82722 552 82728 564
rect 82780 552 82786 604
rect 121822 552 121828 604
rect 121880 592 121886 604
rect 122282 592 122288 604
rect 121880 564 122288 592
rect 121880 552 121886 564
rect 122282 552 122288 564
rect 122340 552 122346 604
rect 124122 552 124128 604
rect 124180 592 124186 604
rect 124674 592 124680 604
rect 124180 564 124680 592
rect 124180 552 124186 564
rect 124674 552 124680 564
rect 124732 552 124738 604
rect 125226 552 125232 604
rect 125284 592 125290 604
rect 125870 592 125876 604
rect 125284 564 125876 592
rect 125284 552 125290 564
rect 125870 552 125876 564
rect 125928 552 125934 604
rect 126422 552 126428 604
rect 126480 592 126486 604
rect 126974 592 126980 604
rect 126480 564 126980 592
rect 126480 552 126486 564
rect 126974 552 126980 564
rect 127032 552 127038 604
rect 127526 552 127532 604
rect 127584 592 127590 604
rect 128170 592 128176 604
rect 127584 564 128176 592
rect 127584 552 127590 564
rect 128170 552 128176 564
rect 128228 552 128234 604
rect 128630 552 128636 604
rect 128688 592 128694 604
rect 129366 592 129372 604
rect 128688 564 129372 592
rect 128688 552 128694 564
rect 129366 552 129372 564
rect 129424 552 129430 604
rect 133874 552 133880 604
rect 133932 592 133938 604
rect 135254 592 135260 604
rect 133932 564 135260 592
rect 133932 552 133938 564
rect 135254 552 135260 564
rect 135312 552 135318 604
rect 136450 552 136456 604
rect 136508 552 136514 604
rect 137554 552 137560 604
rect 137612 592 137618 604
rect 138842 592 138848 604
rect 137612 564 138848 592
rect 137612 552 137618 564
rect 138842 552 138848 564
rect 138900 552 138906 604
rect 139946 552 139952 604
rect 140004 592 140010 604
rect 141234 592 141240 604
rect 140004 564 141240 592
rect 140004 552 140010 564
rect 141234 552 141240 564
rect 141292 552 141298 604
rect 144546 552 144552 604
rect 144604 592 144610 604
rect 145926 592 145932 604
rect 144604 564 145932 592
rect 144604 552 144610 564
rect 145926 552 145932 564
rect 145984 552 145990 604
rect 146846 552 146852 604
rect 146904 592 146910 604
rect 148318 592 148324 604
rect 146904 564 148324 592
rect 146904 552 146910 564
rect 148318 552 148324 564
rect 148376 552 148382 604
rect 152550 552 152556 604
rect 152608 592 152614 604
rect 154206 592 154212 604
rect 152608 564 154212 592
rect 152608 552 152614 564
rect 154206 552 154212 564
rect 154264 552 154270 604
rect 154758 552 154764 604
rect 154816 592 154822 604
rect 156598 592 156604 604
rect 154816 564 156604 592
rect 154816 552 154822 564
rect 156598 552 156604 564
rect 156656 552 156662 604
rect 157058 552 157064 604
rect 157116 592 157122 604
rect 158898 592 158904 604
rect 157116 564 158904 592
rect 157116 552 157122 564
rect 158898 552 158904 564
rect 158956 552 158962 604
rect 161566 552 161572 604
rect 161624 592 161630 604
rect 163682 592 163688 604
rect 161624 564 163688 592
rect 161624 552 161630 564
rect 163682 552 163688 564
rect 163740 552 163746 604
rect 8628 496 10180 524
rect 11164 524 11192 552
rect 14458 524 14464 536
rect 11164 496 14464 524
rect 8628 484 8634 496
rect 14458 484 14464 496
rect 14516 484 14522 536
rect 18506 484 18512 536
rect 18564 524 18570 536
rect 21266 524 21272 536
rect 18564 496 21272 524
rect 18564 484 18570 496
rect 21266 484 21272 496
rect 21324 484 21330 536
rect 22002 484 22008 536
rect 22060 524 22066 536
rect 24826 524 24854 552
rect 22060 496 24854 524
rect 22060 484 22066 496
rect 3234 416 3240 468
rect 3292 456 3298 468
rect 6638 456 6644 468
rect 3292 428 6644 456
rect 3292 416 3298 428
rect 6638 416 6644 428
rect 6696 416 6702 468
rect 24854 416 24860 468
rect 24912 456 24918 468
rect 26878 456 26884 468
rect 24912 428 26884 456
rect 24912 416 24918 428
rect 26878 416 26884 428
rect 26936 416 26942 468
rect 37200 456 37228 552
rect 39592 456 39620 552
rect 50172 524 50200 552
rect 51902 524 51908 536
rect 50172 496 51908 524
rect 51902 484 51908 496
rect 51960 484 51966 536
rect 67726 484 67732 536
rect 67784 524 67790 536
rect 69382 524 69388 536
rect 67784 496 69388 524
rect 67784 484 67790 496
rect 69382 484 69388 496
rect 69440 484 69446 536
rect 134978 484 134984 536
rect 135036 524 135042 536
rect 136468 524 136496 552
rect 135036 496 136496 524
rect 135036 484 135042 496
rect 141050 484 141056 536
rect 141108 524 141114 536
rect 142062 524 142068 536
rect 141108 496 142068 524
rect 141108 484 141114 496
rect 142062 484 142068 496
rect 142120 484 142126 536
rect 158162 484 158168 536
rect 158220 524 158226 536
rect 159726 524 159732 536
rect 158220 496 159732 524
rect 158220 484 158226 496
rect 159726 484 159732 496
rect 159784 484 159790 536
rect 42150 456 42156 468
rect 37200 428 38654 456
rect 39592 428 42156 456
rect 14550 348 14556 400
rect 14608 388 14614 400
rect 17862 388 17868 400
rect 14608 360 17868 388
rect 14608 348 14614 360
rect 17862 348 17868 360
rect 17920 348 17926 400
rect 38626 388 38654 428
rect 42150 416 42156 428
rect 42208 416 42214 468
rect 163406 416 163412 468
rect 163464 456 163470 468
rect 165908 456 165936 632
rect 166074 620 166080 632
rect 166132 620 166138 672
rect 167086 620 167092 672
rect 167144 660 167150 672
rect 169570 660 169576 672
rect 167144 632 169576 660
rect 167144 620 167150 632
rect 169570 620 169576 632
rect 169628 620 169634 672
rect 180886 620 180892 672
rect 180944 660 180950 672
rect 183738 660 183744 672
rect 180944 632 183744 660
rect 180944 620 180950 632
rect 183738 620 183744 632
rect 183796 620 183802 672
rect 186130 660 186136 672
rect 184216 632 186136 660
rect 165982 552 165988 604
rect 166040 592 166046 604
rect 168374 592 168380 604
rect 166040 564 168380 592
rect 166040 552 166046 564
rect 168374 552 168380 564
rect 168432 552 168438 604
rect 170674 552 170680 604
rect 170732 592 170738 604
rect 173158 592 173164 604
rect 170732 564 173164 592
rect 170732 552 170738 564
rect 173158 552 173164 564
rect 173216 552 173222 604
rect 179782 552 179788 604
rect 179840 592 179846 604
rect 182542 592 182548 604
rect 179840 564 182548 592
rect 179840 552 179846 564
rect 182542 552 182548 564
rect 182600 552 182606 604
rect 183186 552 183192 604
rect 183244 592 183250 604
rect 184216 592 184244 632
rect 186130 620 186136 632
rect 186188 620 186194 672
rect 191098 620 191104 672
rect 191156 660 191162 672
rect 194410 660 194416 672
rect 191156 632 194416 660
rect 191156 620 191162 632
rect 194410 620 194416 632
rect 194468 620 194474 672
rect 211614 620 211620 672
rect 211672 660 211678 672
rect 215662 660 215668 672
rect 211672 632 215668 660
rect 211672 620 211678 632
rect 215662 620 215668 632
rect 215720 620 215726 672
rect 219526 620 219532 672
rect 219584 660 219590 672
rect 219584 632 223988 660
rect 219584 620 219590 632
rect 223960 604 223988 632
rect 226150 620 226156 672
rect 226208 660 226214 672
rect 231026 660 231032 672
rect 226208 632 231032 660
rect 226208 620 226214 632
rect 231026 620 231032 632
rect 231084 620 231090 672
rect 234614 660 234620 672
rect 231780 632 234620 660
rect 183244 564 184244 592
rect 183244 552 183250 564
rect 189994 552 190000 604
rect 190052 592 190058 604
rect 193214 592 193220 604
rect 190052 564 193220 592
rect 190052 552 190058 564
rect 193214 552 193220 564
rect 193272 552 193278 604
rect 196802 552 196808 604
rect 196860 552 196866 604
rect 199102 592 199108 604
rect 198706 564 199108 592
rect 187694 484 187700 536
rect 187752 524 187758 536
rect 191006 524 191012 536
rect 187752 496 191012 524
rect 187752 484 187758 496
rect 191006 484 191012 496
rect 191064 484 191070 536
rect 192938 484 192944 536
rect 192996 524 193002 536
rect 196820 524 196848 552
rect 192996 496 196848 524
rect 192996 484 193002 496
rect 163464 428 165936 456
rect 163464 416 163470 428
rect 39850 388 39856 400
rect 38626 360 39856 388
rect 39850 348 39856 360
rect 39908 348 39914 400
rect 42886 348 42892 400
rect 42944 388 42950 400
rect 45094 388 45100 400
rect 42944 360 45100 388
rect 42944 348 42950 360
rect 45094 348 45100 360
rect 45152 348 45158 400
rect 71314 348 71320 400
rect 71372 388 71378 400
rect 72326 388 72332 400
rect 71372 360 72332 388
rect 71372 348 71378 360
rect 72326 348 72332 360
rect 72384 348 72390 400
rect 72418 348 72424 400
rect 72476 388 72482 400
rect 73522 388 73528 400
rect 72476 360 73528 388
rect 72476 348 72482 360
rect 73522 348 73528 360
rect 73580 348 73586 400
rect 73614 348 73620 400
rect 73672 388 73678 400
rect 74626 388 74632 400
rect 73672 360 74632 388
rect 73672 348 73678 360
rect 74626 348 74632 360
rect 74684 348 74690 400
rect 130930 348 130936 400
rect 130988 388 130994 400
rect 131942 388 131948 400
rect 130988 360 131948 388
rect 130988 348 130994 360
rect 131942 348 131948 360
rect 132000 348 132006 400
rect 132034 348 132040 400
rect 132092 388 132098 400
rect 133138 388 133144 400
rect 132092 360 133144 388
rect 132092 348 132098 360
rect 133138 348 133144 360
rect 133196 348 133202 400
rect 160462 348 160468 400
rect 160520 388 160526 400
rect 162670 388 162676 400
rect 160520 360 162676 388
rect 160520 348 160526 360
rect 162670 348 162676 360
rect 162728 348 162734 400
rect 195238 348 195244 400
rect 195296 388 195302 400
rect 198706 388 198734 564
rect 199102 552 199108 564
rect 199160 552 199166 604
rect 203610 552 203616 604
rect 203668 592 203674 604
rect 204162 592 204168 604
rect 203668 564 204168 592
rect 203668 552 203674 564
rect 204162 552 204168 564
rect 204220 552 204226 604
rect 205726 552 205732 604
rect 205784 592 205790 604
rect 209774 592 209780 604
rect 205784 564 209780 592
rect 205784 552 205790 564
rect 209774 552 209780 564
rect 209832 552 209838 604
rect 210418 552 210424 604
rect 210476 592 210482 604
rect 212077 595 212135 601
rect 212077 592 212089 595
rect 210476 564 212089 592
rect 210476 552 210482 564
rect 212077 561 212089 564
rect 212123 561 212135 595
rect 212077 555 212135 561
rect 212166 552 212172 604
rect 212224 552 212230 604
rect 212261 595 212319 601
rect 212261 561 212273 595
rect 212307 592 212319 595
rect 214466 592 214472 604
rect 212307 564 214472 592
rect 212307 561 212319 564
rect 212261 555 212319 561
rect 214466 552 214472 564
rect 214524 552 214530 604
rect 218422 552 218428 604
rect 218480 592 218486 604
rect 222746 592 222752 604
rect 218480 564 222752 592
rect 218480 552 218486 564
rect 222746 552 222752 564
rect 222804 552 222810 604
rect 223942 552 223948 604
rect 224000 552 224006 604
rect 225046 552 225052 604
rect 225104 592 225110 604
rect 229830 592 229836 604
rect 225104 564 227714 592
rect 225104 552 225110 564
rect 208394 484 208400 536
rect 208452 524 208458 536
rect 212184 524 212212 552
rect 208452 496 212212 524
rect 224589 527 224647 533
rect 208452 484 208458 496
rect 224589 493 224601 527
rect 224635 524 224647 527
rect 225322 524 225328 536
rect 224635 496 225328 524
rect 224635 493 224647 496
rect 224589 487 224647 493
rect 225322 484 225328 496
rect 225380 484 225386 536
rect 226518 484 226524 536
rect 226576 484 226582 536
rect 227686 524 227714 564
rect 229066 564 229836 592
rect 229066 524 229094 564
rect 229830 552 229836 564
rect 229888 552 229894 604
rect 227686 496 229094 524
rect 229646 484 229652 536
rect 229704 524 229710 536
rect 231780 524 231808 632
rect 234614 620 234620 632
rect 234672 620 234678 672
rect 235442 620 235448 672
rect 235500 660 235506 672
rect 237346 660 237374 700
rect 240505 697 240517 700
rect 240551 697 240563 731
rect 283101 731 283159 737
rect 283101 728 283113 731
rect 240505 691 240563 697
rect 275986 700 283113 728
rect 235500 632 237374 660
rect 235500 620 235506 632
rect 237742 620 237748 672
rect 237800 660 237806 672
rect 242894 660 242900 672
rect 237800 632 242900 660
rect 237800 620 237806 632
rect 242894 620 242900 632
rect 242952 620 242958 672
rect 247954 620 247960 672
rect 248012 660 248018 672
rect 253474 660 253480 672
rect 248012 632 253480 660
rect 248012 620 248018 632
rect 253474 620 253480 632
rect 253532 620 253538 672
rect 255774 620 255780 672
rect 255832 660 255838 672
rect 261754 660 261760 672
rect 255832 632 261760 660
rect 255832 620 255838 632
rect 261754 620 261760 632
rect 261812 620 261818 672
rect 262674 620 262680 672
rect 262732 660 262738 672
rect 268838 660 268844 672
rect 262732 632 268844 660
rect 262732 620 262738 632
rect 268838 620 268844 632
rect 268896 620 268902 672
rect 275830 620 275836 672
rect 275888 660 275894 672
rect 275986 660 276014 700
rect 283101 697 283113 700
rect 283147 697 283159 731
rect 283101 691 283159 697
rect 275888 632 276014 660
rect 275888 620 275894 632
rect 277486 620 277492 672
rect 277544 660 277550 672
rect 284294 660 284300 672
rect 277544 632 284300 660
rect 277544 620 277550 632
rect 284294 620 284300 632
rect 284352 620 284358 672
rect 284573 663 284631 669
rect 284573 629 284585 663
rect 284619 660 284631 663
rect 286594 660 286600 672
rect 284619 632 286600 660
rect 284619 629 284631 632
rect 284573 623 284631 629
rect 286594 620 286600 632
rect 286652 620 286658 672
rect 288360 660 288388 768
rect 321526 768 324314 796
rect 292546 700 298508 728
rect 288986 660 288992 672
rect 288360 632 288992 660
rect 288986 620 288992 632
rect 289044 620 289050 672
rect 291102 620 291108 672
rect 291160 660 291166 672
rect 292546 660 292574 700
rect 298480 672 298508 700
rect 304966 700 309088 728
rect 291160 632 292574 660
rect 291160 620 291166 632
rect 293402 620 293408 672
rect 293460 660 293466 672
rect 293460 632 298416 660
rect 293460 620 293466 632
rect 231854 552 231860 604
rect 231912 592 231918 604
rect 237006 592 237012 604
rect 231912 564 237012 592
rect 231912 552 231918 564
rect 237006 552 237012 564
rect 237064 552 237070 604
rect 238110 552 238116 604
rect 238168 552 238174 604
rect 239306 592 239312 604
rect 238404 564 239312 592
rect 229704 496 231808 524
rect 229704 484 229710 496
rect 233142 484 233148 536
rect 233200 524 233206 536
rect 238128 524 238156 552
rect 233200 496 238156 524
rect 233200 484 233206 496
rect 212534 416 212540 468
rect 212592 456 212598 468
rect 216582 456 216588 468
rect 212592 428 216588 456
rect 212592 416 212598 428
rect 216582 416 216588 428
rect 216640 416 216646 468
rect 221826 416 221832 468
rect 221884 456 221890 468
rect 226536 456 226564 484
rect 221884 428 226564 456
rect 221884 416 221890 428
rect 234338 416 234344 468
rect 234396 456 234402 468
rect 238404 456 238432 564
rect 239306 552 239312 564
rect 239364 552 239370 604
rect 240502 592 240508 604
rect 240463 564 240508 592
rect 240502 552 240508 564
rect 240560 552 240566 604
rect 249978 552 249984 604
rect 250036 552 250042 604
rect 251174 592 251180 604
rect 251135 564 251180 592
rect 251174 552 251180 564
rect 251232 552 251238 604
rect 252278 552 252284 604
rect 252336 592 252342 604
rect 252336 564 252554 592
rect 252336 552 252342 564
rect 244550 484 244556 536
rect 244608 524 244614 536
rect 249996 524 250024 552
rect 244608 496 250024 524
rect 252526 524 252554 564
rect 254578 552 254584 604
rect 254636 592 254642 604
rect 260650 592 260656 604
rect 254636 564 260656 592
rect 254636 552 254642 564
rect 260650 552 260656 564
rect 260708 552 260714 604
rect 266538 592 266544 604
rect 261496 564 266544 592
rect 258074 524 258080 536
rect 252526 496 258080 524
rect 244608 484 244614 496
rect 258074 484 258080 496
rect 258132 484 258138 536
rect 260466 484 260472 536
rect 260524 524 260530 536
rect 261496 524 261524 564
rect 266538 552 266544 564
rect 266596 552 266602 604
rect 267734 552 267740 604
rect 267792 552 267798 604
rect 270034 592 270040 604
rect 268212 564 270040 592
rect 260524 496 261524 524
rect 260524 484 260530 496
rect 261570 484 261576 536
rect 261628 524 261634 536
rect 267752 524 267780 552
rect 261628 496 267780 524
rect 261628 484 261634 496
rect 234396 428 238432 456
rect 234396 416 234402 428
rect 239950 416 239956 468
rect 240008 456 240014 468
rect 244918 456 244924 468
rect 240008 428 244924 456
rect 240008 416 240014 428
rect 244918 416 244924 428
rect 244976 416 244982 468
rect 246758 416 246764 468
rect 246816 456 246822 468
rect 252554 456 252560 468
rect 246816 428 252560 456
rect 246816 416 246822 428
rect 252554 416 252560 428
rect 252612 416 252618 468
rect 259086 416 259092 468
rect 259144 416 259150 468
rect 263686 416 263692 468
rect 263744 456 263750 468
rect 268212 456 268240 564
rect 270034 552 270040 564
rect 270092 552 270098 604
rect 271782 552 271788 604
rect 271840 592 271846 604
rect 271840 564 278544 592
rect 271840 552 271846 564
rect 278516 536 278544 564
rect 279510 552 279516 604
rect 279568 552 279574 604
rect 280706 592 280712 604
rect 280667 564 280712 592
rect 280706 552 280712 564
rect 280764 552 280770 604
rect 281810 592 281816 604
rect 281771 564 281816 592
rect 281810 552 281816 564
rect 281868 552 281874 604
rect 283098 592 283104 604
rect 283059 564 283104 592
rect 283098 552 283104 564
rect 283156 552 283162 604
rect 288802 552 288808 604
rect 288860 592 288866 604
rect 296070 592 296076 604
rect 288860 564 296076 592
rect 288860 552 288866 564
rect 296070 552 296076 564
rect 296128 552 296134 604
rect 297266 592 297272 604
rect 297227 564 297272 592
rect 297266 552 297272 564
rect 297324 552 297330 604
rect 298388 592 298416 632
rect 298462 620 298468 672
rect 298520 620 298526 672
rect 300762 660 300768 672
rect 299584 632 300768 660
rect 299584 592 299612 632
rect 300762 620 300768 632
rect 300820 620 300826 672
rect 301314 620 301320 672
rect 301372 660 301378 672
rect 304966 660 304994 700
rect 309060 672 309088 700
rect 307662 660 307668 672
rect 301372 632 304994 660
rect 307623 632 307668 660
rect 301372 620 301378 632
rect 307662 620 307668 632
rect 307720 620 307726 672
rect 309042 620 309048 672
rect 309100 620 309106 672
rect 311342 620 311348 672
rect 311400 660 311406 672
rect 315853 663 315911 669
rect 315853 660 315865 663
rect 311400 632 315865 660
rect 311400 620 311406 632
rect 315853 629 315865 632
rect 315899 629 315911 663
rect 315853 623 315911 629
rect 315942 620 315948 672
rect 316000 660 316006 672
rect 316000 632 318288 660
rect 316000 620 316006 632
rect 298388 564 299612 592
rect 299658 552 299664 604
rect 299716 552 299722 604
rect 301958 592 301964 604
rect 299768 564 301964 592
rect 268378 484 268384 536
rect 268436 524 268442 536
rect 274542 524 274548 536
rect 268436 496 274548 524
rect 268436 484 268442 496
rect 274542 484 274548 496
rect 274600 484 274606 536
rect 278498 484 278504 536
rect 278556 484 278562 536
rect 263744 428 268240 456
rect 263744 416 263750 428
rect 270678 416 270684 468
rect 270736 456 270742 468
rect 276750 456 276756 468
rect 270736 428 276756 456
rect 270736 416 270742 428
rect 276750 416 276756 428
rect 276808 416 276814 468
rect 195296 360 198734 388
rect 195296 348 195302 360
rect 217226 348 217232 400
rect 217284 388 217290 400
rect 221734 388 221740 400
rect 217284 360 221740 388
rect 217284 348 217290 360
rect 221734 348 221740 360
rect 221792 348 221798 400
rect 222470 348 222476 400
rect 222528 388 222534 400
rect 227254 388 227260 400
rect 222528 360 227260 388
rect 222528 348 222534 360
rect 227254 348 227260 360
rect 227312 348 227318 400
rect 245654 348 245660 400
rect 245712 388 245718 400
rect 251177 391 251235 397
rect 251177 388 251189 391
rect 245712 360 251189 388
rect 245712 348 245718 360
rect 251177 357 251189 360
rect 251223 357 251235 391
rect 251177 351 251235 357
rect 253106 348 253112 400
rect 253164 388 253170 400
rect 259104 388 259132 416
rect 253164 360 259132 388
rect 253164 348 253170 360
rect 259270 348 259276 400
rect 259328 388 259334 400
rect 264974 388 264980 400
rect 259328 360 264980 388
rect 259328 348 259334 360
rect 264974 348 264980 360
rect 265032 348 265038 400
rect 272886 348 272892 400
rect 272944 388 272950 400
rect 279528 388 279556 552
rect 292206 484 292212 536
rect 292264 524 292270 536
rect 299676 524 299704 552
rect 292264 496 299704 524
rect 292264 484 292270 496
rect 280430 416 280436 468
rect 280488 456 280494 468
rect 285674 456 285680 468
rect 280488 428 285680 456
rect 280488 416 280494 428
rect 285674 416 285680 428
rect 285732 416 285738 468
rect 287606 416 287612 468
rect 287664 456 287670 468
rect 293862 456 293868 468
rect 287664 428 293868 456
rect 287664 416 287670 428
rect 293862 416 293868 428
rect 293920 416 293926 468
rect 272944 360 279556 388
rect 272944 348 272950 360
rect 294506 348 294512 400
rect 294564 388 294570 400
rect 299768 388 299796 564
rect 301958 552 301964 564
rect 302016 552 302022 604
rect 307941 595 307999 601
rect 307941 561 307953 595
rect 307987 592 307999 595
rect 308030 592 308036 604
rect 307987 564 308036 592
rect 307987 561 307999 564
rect 307941 555 307999 561
rect 308030 552 308036 564
rect 308088 552 308094 604
rect 310238 592 310244 604
rect 310199 564 310244 592
rect 310238 552 310244 564
rect 310296 552 310302 604
rect 311434 592 311440 604
rect 311395 564 311440 592
rect 311434 552 311440 564
rect 311492 552 311498 604
rect 312630 592 312636 604
rect 312591 564 312636 592
rect 312630 552 312636 564
rect 312688 552 312694 604
rect 317322 592 317328 604
rect 314626 564 317328 592
rect 300210 484 300216 536
rect 300268 524 300274 536
rect 307849 527 307907 533
rect 307849 524 307861 527
rect 300268 496 307861 524
rect 300268 484 300274 496
rect 307849 493 307861 496
rect 307895 493 307907 527
rect 307849 487 307907 493
rect 308766 484 308772 536
rect 308824 524 308830 536
rect 314626 524 314654 564
rect 317322 552 317328 564
rect 317380 552 317386 604
rect 318260 592 318288 632
rect 318334 620 318340 672
rect 318392 660 318398 672
rect 321526 660 321554 768
rect 318392 632 321554 660
rect 324286 660 324314 768
rect 383120 768 394280 796
rect 369397 731 369455 737
rect 369397 728 369409 731
rect 359292 700 369409 728
rect 359292 672 359320 700
rect 369397 697 369409 700
rect 369443 697 369455 731
rect 371789 731 371847 737
rect 371789 728 371801 731
rect 369397 691 369455 697
rect 371528 700 371801 728
rect 326798 660 326804 672
rect 324286 632 326804 660
rect 318392 620 318398 632
rect 326798 620 326804 632
rect 326856 620 326862 672
rect 327442 620 327448 672
rect 327500 660 327506 672
rect 327500 632 336504 660
rect 327500 620 327506 632
rect 324406 592 324412 604
rect 318260 564 324412 592
rect 324406 552 324412 564
rect 324464 552 324470 604
rect 325602 552 325608 604
rect 325660 552 325666 604
rect 326338 552 326344 604
rect 326396 592 326402 604
rect 335262 592 335268 604
rect 326396 564 335268 592
rect 326396 552 326402 564
rect 335262 552 335268 564
rect 335320 552 335326 604
rect 316034 524 316040 536
rect 308824 496 314654 524
rect 315995 496 316040 524
rect 308824 484 308830 496
rect 316034 484 316040 496
rect 316092 484 316098 536
rect 317138 484 317144 536
rect 317196 524 317202 536
rect 325620 524 325648 552
rect 336476 536 336504 632
rect 339770 620 339776 672
rect 339828 660 339834 672
rect 339828 632 342254 660
rect 339828 620 339834 632
rect 336642 552 336648 604
rect 336700 592 336706 604
rect 337470 592 337476 604
rect 336700 564 337476 592
rect 336700 552 336706 564
rect 337470 552 337476 564
rect 337528 552 337534 604
rect 338666 592 338672 604
rect 338627 564 338672 592
rect 338666 552 338672 564
rect 338724 552 338730 604
rect 339862 592 339868 604
rect 339823 564 339868 592
rect 339862 552 339868 564
rect 339920 552 339926 604
rect 340966 592 340972 604
rect 340927 564 340972 592
rect 340966 552 340972 564
rect 341024 552 341030 604
rect 342226 592 342254 632
rect 343174 620 343180 672
rect 343232 660 343238 672
rect 352834 660 352840 672
rect 343232 632 352840 660
rect 343232 620 343238 632
rect 352834 620 352840 632
rect 352892 620 352898 672
rect 354585 663 354643 669
rect 354585 629 354597 663
rect 354631 660 354643 663
rect 354631 632 358814 660
rect 354631 629 354643 632
rect 354585 623 354643 629
rect 349246 592 349252 604
rect 342226 564 349252 592
rect 349246 552 349252 564
rect 349304 552 349310 604
rect 357526 592 357532 604
rect 350506 564 357532 592
rect 317196 496 325648 524
rect 317196 484 317202 496
rect 336458 484 336464 536
rect 336516 484 336522 536
rect 337194 484 337200 536
rect 337252 524 337258 536
rect 346762 524 346768 536
rect 337252 496 346768 524
rect 337252 484 337258 496
rect 346762 484 346768 496
rect 346820 484 346826 536
rect 347682 484 347688 536
rect 347740 524 347746 536
rect 350506 524 350534 564
rect 357526 552 357532 564
rect 357584 552 357590 604
rect 358786 592 358814 632
rect 359274 620 359280 672
rect 359332 620 359338 672
rect 360378 620 360384 672
rect 360436 660 360442 672
rect 363782 660 363788 672
rect 360436 632 363788 660
rect 360436 620 360442 632
rect 363782 620 363788 632
rect 363840 620 363846 672
rect 366082 620 366088 672
rect 366140 660 366146 672
rect 371528 660 371556 700
rect 371789 697 371801 700
rect 371835 697 371847 731
rect 371789 691 371847 697
rect 372586 700 380848 728
rect 366140 632 371556 660
rect 366140 620 366146 632
rect 371602 620 371608 672
rect 371660 660 371666 672
rect 372586 660 372614 700
rect 371660 632 372614 660
rect 371660 620 371666 632
rect 373902 620 373908 672
rect 373960 660 373966 672
rect 380820 660 380848 700
rect 383120 672 383148 768
rect 394252 672 394280 768
rect 404326 768 407160 796
rect 404326 728 404354 768
rect 396046 700 404354 728
rect 382366 660 382372 672
rect 373960 632 380756 660
rect 380820 632 382372 660
rect 373960 620 373966 632
rect 361942 592 361948 604
rect 358786 564 361948 592
rect 361942 552 361948 564
rect 362000 552 362006 604
rect 367002 592 367008 604
rect 366963 564 367008 592
rect 367002 552 367008 564
rect 367060 552 367066 604
rect 368198 592 368204 604
rect 368159 564 368204 592
rect 368198 552 368204 564
rect 368256 552 368262 604
rect 369394 592 369400 604
rect 369355 564 369400 592
rect 369394 552 369400 564
rect 369452 552 369458 604
rect 371694 552 371700 604
rect 371752 552 371758 604
rect 371789 595 371847 601
rect 371789 561 371801 595
rect 371835 592 371847 595
rect 376478 592 376484 604
rect 371835 564 376484 592
rect 371835 561 371847 564
rect 371789 555 371847 561
rect 376478 552 376484 564
rect 376536 552 376542 604
rect 379514 552 379520 604
rect 379572 592 379578 604
rect 380621 595 380679 601
rect 380621 592 380633 595
rect 379572 564 380633 592
rect 379572 552 379578 564
rect 380621 561 380633 564
rect 380667 561 380679 595
rect 380621 555 380679 561
rect 347740 496 350534 524
rect 347740 484 347746 496
rect 352466 484 352472 536
rect 352524 524 352530 536
rect 354585 527 354643 533
rect 354585 524 354597 527
rect 352524 496 354597 524
rect 352524 484 352530 496
rect 354585 493 354597 496
rect 354631 493 354643 527
rect 354585 487 354643 493
rect 354674 484 354680 536
rect 354732 524 354738 536
rect 354732 496 358814 524
rect 354732 484 354738 496
rect 303614 416 303620 468
rect 303672 456 303678 468
rect 311437 459 311495 465
rect 311437 456 311449 459
rect 303672 428 311449 456
rect 303672 416 303678 428
rect 311437 425 311449 428
rect 311483 425 311495 459
rect 311437 419 311495 425
rect 312446 416 312452 468
rect 312504 456 312510 468
rect 320726 456 320732 468
rect 312504 428 320732 456
rect 312504 416 312510 428
rect 320726 416 320732 428
rect 320784 416 320790 468
rect 321830 456 321836 468
rect 320928 428 321836 456
rect 294564 360 299796 388
rect 294564 348 294570 360
rect 304718 348 304724 400
rect 304776 388 304782 400
rect 312633 391 312691 397
rect 312633 388 312645 391
rect 304776 360 312645 388
rect 304776 348 304782 360
rect 312633 357 312645 360
rect 312679 357 312691 391
rect 314838 388 314844 400
rect 312633 351 312691 357
rect 313246 360 314844 388
rect 220170 280 220176 332
rect 220228 320 220234 332
rect 224589 323 224647 329
rect 224589 320 224601 323
rect 220228 292 224601 320
rect 220228 280 220234 292
rect 224589 289 224601 292
rect 224635 289 224647 323
rect 224589 283 224647 289
rect 243354 280 243360 332
rect 243412 320 243418 332
rect 248966 320 248972 332
rect 243412 292 248972 320
rect 243412 280 243418 292
rect 248966 280 248972 292
rect 249024 280 249030 332
rect 249702 280 249708 332
rect 249760 320 249766 332
rect 255222 320 255228 332
rect 249760 292 255228 320
rect 249760 280 249766 292
rect 255222 280 255228 292
rect 255280 280 255286 332
rect 256878 280 256884 332
rect 256936 320 256942 332
rect 262766 320 262772 332
rect 256936 292 262772 320
rect 256936 280 256942 292
rect 262766 280 262772 292
rect 262824 280 262830 332
rect 279234 280 279240 332
rect 279292 320 279298 332
rect 284573 323 284631 329
rect 284573 320 284585 323
rect 279292 292 284585 320
rect 279292 280 279298 292
rect 284573 289 284585 292
rect 284619 289 284631 323
rect 284573 283 284631 289
rect 289814 280 289820 332
rect 289872 320 289878 332
rect 297269 323 297327 329
rect 297269 320 297281 323
rect 289872 292 297281 320
rect 289872 280 289878 292
rect 297269 289 297281 292
rect 297315 289 297327 323
rect 297269 283 297327 289
rect 297910 280 297916 332
rect 297968 320 297974 332
rect 305730 320 305736 332
rect 297968 292 305736 320
rect 297968 280 297974 292
rect 305730 280 305736 292
rect 305788 280 305794 332
rect 307018 280 307024 332
rect 307076 320 307082 332
rect 313246 320 313274 360
rect 314838 348 314844 360
rect 314896 348 314902 400
rect 315853 391 315911 397
rect 315853 357 315865 391
rect 315899 388 315911 391
rect 318886 388 318892 400
rect 315899 360 318892 388
rect 315899 357 315911 360
rect 315853 351 315911 357
rect 318886 348 318892 360
rect 318944 348 318950 400
rect 307076 292 313274 320
rect 307076 280 307082 292
rect 313642 280 313648 332
rect 313700 320 313706 332
rect 320928 320 320956 428
rect 321830 416 321836 428
rect 321888 416 321894 468
rect 325142 416 325148 468
rect 325200 456 325206 468
rect 325200 428 329834 456
rect 325200 416 325206 428
rect 327810 388 327816 400
rect 321526 360 327816 388
rect 321526 320 321554 360
rect 327810 348 327816 360
rect 327868 348 327874 400
rect 329806 388 329834 428
rect 330846 416 330852 468
rect 330904 456 330910 468
rect 339865 459 339923 465
rect 339865 456 339877 459
rect 330904 428 339877 456
rect 330904 416 330910 428
rect 339865 425 339877 428
rect 339911 425 339923 459
rect 339865 419 339923 425
rect 340598 416 340604 468
rect 340656 456 340662 468
rect 348418 456 348424 468
rect 340656 428 348424 456
rect 340656 416 340662 428
rect 348418 416 348424 428
rect 348476 416 348482 468
rect 353570 416 353576 468
rect 353628 456 353634 468
rect 357805 459 357863 465
rect 357805 456 357817 459
rect 353628 428 357817 456
rect 353628 416 353634 428
rect 357805 425 357817 428
rect 357851 425 357863 459
rect 358786 456 358814 496
rect 361482 484 361488 536
rect 361540 524 361546 536
rect 361540 496 369854 524
rect 361540 484 361546 496
rect 364794 456 364800 468
rect 358786 428 364800 456
rect 357805 419 357863 425
rect 364794 416 364800 428
rect 364852 416 364858 468
rect 369826 456 369854 496
rect 371712 456 371740 552
rect 371881 527 371939 533
rect 371881 493 371893 527
rect 371927 524 371939 527
rect 374362 524 374368 536
rect 371927 496 374368 524
rect 371927 493 371939 496
rect 371881 487 371939 493
rect 374362 484 374368 496
rect 374420 484 374426 536
rect 377398 484 377404 536
rect 377456 524 377462 536
rect 380728 524 380756 632
rect 382366 620 382372 632
rect 382424 620 382430 672
rect 383102 620 383108 672
rect 383160 620 383166 672
rect 390278 660 390284 672
rect 383626 632 390284 660
rect 380805 595 380863 601
rect 380805 561 380817 595
rect 380851 592 380863 595
rect 383626 592 383654 632
rect 390278 620 390284 632
rect 390336 620 390342 672
rect 392210 660 392216 672
rect 392171 632 392216 660
rect 392210 620 392216 632
rect 392268 620 392274 672
rect 394234 620 394240 672
rect 394292 620 394298 672
rect 395614 620 395620 672
rect 395672 660 395678 672
rect 396046 660 396074 700
rect 400309 663 400367 669
rect 395672 632 396074 660
rect 397426 632 400260 660
rect 395672 620 395678 632
rect 385954 592 385960 604
rect 380851 564 383654 592
rect 385915 564 385960 592
rect 380851 561 380863 564
rect 380805 555 380863 561
rect 385954 552 385960 564
rect 386012 552 386018 604
rect 388254 592 388260 604
rect 387766 564 388260 592
rect 381998 524 382004 536
rect 377456 496 380664 524
rect 380728 496 382004 524
rect 377456 484 377462 496
rect 369826 428 371740 456
rect 372706 416 372712 468
rect 372764 456 372770 468
rect 379606 456 379612 468
rect 372764 428 379612 456
rect 372764 416 372770 428
rect 379606 416 379612 428
rect 379664 416 379670 468
rect 380636 456 380664 496
rect 381998 484 382004 496
rect 382056 484 382062 536
rect 387766 456 387794 564
rect 388254 552 388260 564
rect 388312 552 388318 604
rect 393314 552 393320 604
rect 393372 592 393378 604
rect 397426 592 397454 632
rect 400122 592 400128 604
rect 393372 564 397454 592
rect 397748 564 400128 592
rect 393372 552 393378 564
rect 388806 484 388812 536
rect 388864 524 388870 536
rect 397748 524 397776 564
rect 400122 552 400128 564
rect 400180 552 400186 604
rect 400232 592 400260 632
rect 400309 629 400321 663
rect 400355 660 400367 663
rect 403066 660 403072 672
rect 400355 632 403072 660
rect 400355 629 400367 632
rect 400309 623 400367 629
rect 403066 620 403072 632
rect 403124 620 403130 672
rect 403434 620 403440 672
rect 403492 660 403498 672
rect 407132 660 407160 768
rect 408466 728 408494 972
rect 419905 969 419917 972
rect 419951 969 419963 1003
rect 419905 963 419963 969
rect 426989 1003 427047 1009
rect 426989 969 427001 1003
rect 427035 1000 427047 1003
rect 440145 1003 440203 1009
rect 440145 1000 440157 1003
rect 427035 972 440157 1000
rect 427035 969 427047 972
rect 426989 963 427047 969
rect 440145 969 440157 972
rect 440191 969 440203 1003
rect 440145 963 440203 969
rect 441065 1003 441123 1009
rect 441065 969 441077 1003
rect 441111 1000 441123 1003
rect 454405 1003 454463 1009
rect 454405 1000 454417 1003
rect 441111 972 454417 1000
rect 441111 969 441123 972
rect 441065 963 441123 969
rect 454405 969 454417 972
rect 454451 969 454463 1003
rect 454405 963 454463 969
rect 457993 1003 458051 1009
rect 457993 969 458005 1003
rect 458039 1000 458051 1003
rect 466365 1003 466423 1009
rect 466365 1000 466377 1003
rect 458039 972 466377 1000
rect 458039 969 458051 972
rect 457993 963 458051 969
rect 466365 969 466377 972
rect 466411 969 466423 1003
rect 466365 963 466423 969
rect 471793 1003 471851 1009
rect 471793 969 471805 1003
rect 471839 1000 471851 1003
rect 480809 1003 480867 1009
rect 480809 1000 480821 1003
rect 471839 972 480821 1000
rect 471839 969 471851 972
rect 471793 963 471851 969
rect 480809 969 480821 972
rect 480855 969 480867 1003
rect 480809 963 480867 969
rect 487433 1003 487491 1009
rect 487433 969 487445 1003
rect 487479 1000 487491 1003
rect 490668 1000 490696 1108
rect 502981 1105 502993 1108
rect 503027 1105 503039 1139
rect 502981 1099 503039 1105
rect 510341 1139 510399 1145
rect 510341 1105 510353 1139
rect 510387 1136 510399 1139
rect 526625 1139 526683 1145
rect 526625 1136 526637 1139
rect 510387 1108 526637 1136
rect 510387 1105 510399 1108
rect 510341 1099 510399 1105
rect 526625 1105 526637 1108
rect 526671 1105 526683 1139
rect 526625 1099 526683 1105
rect 500129 1071 500187 1077
rect 500129 1037 500141 1071
rect 500175 1068 500187 1071
rect 515401 1071 515459 1077
rect 515401 1068 515413 1071
rect 500175 1040 515413 1068
rect 500175 1037 500187 1040
rect 500129 1031 500187 1037
rect 515401 1037 515413 1040
rect 515447 1037 515459 1071
rect 515401 1031 515459 1037
rect 555789 1071 555847 1077
rect 555789 1037 555801 1071
rect 555835 1068 555847 1071
rect 563514 1068 563520 1080
rect 555835 1040 563520 1068
rect 555835 1037 555847 1040
rect 555789 1031 555847 1037
rect 563514 1028 563520 1040
rect 563572 1028 563578 1080
rect 487479 972 490696 1000
rect 493321 1003 493379 1009
rect 487479 969 487491 972
rect 487433 963 487491 969
rect 493321 969 493333 1003
rect 493367 1000 493379 1003
rect 508593 1003 508651 1009
rect 508593 1000 508605 1003
rect 493367 972 508605 1000
rect 493367 969 493379 972
rect 493321 963 493379 969
rect 508593 969 508605 972
rect 508639 969 508651 1003
rect 508593 963 508651 969
rect 512181 1003 512239 1009
rect 512181 969 512193 1003
rect 512227 1000 512239 1003
rect 529017 1003 529075 1009
rect 529017 1000 529029 1003
rect 512227 972 529029 1000
rect 512227 969 512239 972
rect 512181 963 512239 969
rect 529017 969 529029 972
rect 529063 969 529075 1003
rect 529017 963 529075 969
rect 548889 1003 548947 1009
rect 548889 969 548901 1003
rect 548935 1000 548947 1003
rect 558181 1003 558239 1009
rect 558181 1000 558193 1003
rect 548935 972 558193 1000
rect 548935 969 548947 972
rect 548889 963 548947 969
rect 558181 969 558193 972
rect 558227 969 558239 1003
rect 558181 963 558239 969
rect 558733 1003 558791 1009
rect 558733 969 558745 1003
rect 558779 1000 558791 1003
rect 569126 1000 569132 1012
rect 558779 972 569132 1000
rect 558779 969 558791 972
rect 558733 963 558791 969
rect 569126 960 569132 972
rect 569184 960 569190 1012
rect 417145 935 417203 941
rect 417145 901 417157 935
rect 417191 932 417203 935
rect 427909 935 427967 941
rect 427909 932 427921 935
rect 417191 904 427921 932
rect 417191 901 417203 904
rect 417145 895 417203 901
rect 427909 901 427921 904
rect 427955 901 427967 935
rect 455877 935 455935 941
rect 455877 932 455889 935
rect 427909 895 427967 901
rect 443196 904 455889 932
rect 434441 867 434499 873
rect 434441 864 434453 867
rect 411226 836 421144 864
rect 408144 700 408494 728
rect 409233 731 409291 737
rect 408144 672 408172 700
rect 409233 697 409245 731
rect 409279 728 409291 731
rect 411226 728 411254 836
rect 418617 799 418675 805
rect 418617 796 418629 799
rect 409279 700 411254 728
rect 416608 768 418629 796
rect 409279 697 409291 700
rect 409233 691 409291 697
rect 407206 660 407212 672
rect 403492 632 407068 660
rect 407132 632 407212 660
rect 403492 620 403498 632
rect 404814 592 404820 604
rect 400232 564 404820 592
rect 404814 552 404820 564
rect 404872 552 404878 604
rect 405366 592 405372 604
rect 405327 564 405372 592
rect 405366 552 405372 564
rect 405424 552 405430 604
rect 407040 592 407068 632
rect 407206 620 407212 632
rect 407264 620 407270 672
rect 408126 620 408132 672
rect 408184 620 408190 672
rect 415486 660 415492 672
rect 408466 632 415492 660
rect 408466 592 408494 632
rect 415486 620 415492 632
rect 415544 620 415550 672
rect 409230 592 409236 604
rect 407040 564 408494 592
rect 409191 564 409236 592
rect 409230 552 409236 564
rect 409288 552 409294 604
rect 412634 552 412640 604
rect 412692 592 412698 604
rect 416608 592 416636 768
rect 418617 765 418629 768
rect 418663 765 418675 799
rect 418617 759 418675 765
rect 416685 731 416743 737
rect 416685 697 416697 731
rect 416731 728 416743 731
rect 416731 700 420914 728
rect 416731 697 416743 700
rect 416685 691 416743 697
rect 420886 660 420914 700
rect 421116 672 421144 836
rect 425026 836 434453 864
rect 421006 660 421012 672
rect 420886 632 421012 660
rect 421006 620 421012 632
rect 421064 620 421070 672
rect 421098 620 421104 672
rect 421156 620 421162 672
rect 421742 620 421748 672
rect 421800 660 421806 672
rect 425026 660 425054 836
rect 434441 833 434453 836
rect 434487 833 434499 867
rect 434441 827 434499 833
rect 439133 799 439191 805
rect 439133 796 439145 799
rect 428016 768 439145 796
rect 428016 728 428044 768
rect 439133 765 439145 768
rect 439179 765 439191 799
rect 439133 759 439191 765
rect 428553 731 428611 737
rect 428553 728 428565 731
rect 426084 700 428044 728
rect 428108 700 428565 728
rect 426084 672 426112 700
rect 421800 632 425054 660
rect 421800 620 421806 632
rect 426066 620 426072 672
rect 426124 620 426130 672
rect 426342 620 426348 672
rect 426400 660 426406 672
rect 426986 660 426992 672
rect 426400 632 426445 660
rect 426947 632 426992 660
rect 426400 620 426406 632
rect 426986 620 426992 632
rect 427044 620 427050 672
rect 427262 660 427268 672
rect 427223 632 427268 660
rect 427262 620 427268 632
rect 427320 620 427326 672
rect 427906 660 427912 672
rect 427867 632 427912 660
rect 427906 620 427912 632
rect 427964 620 427970 672
rect 417142 592 417148 604
rect 412692 564 416636 592
rect 417103 564 417148 592
rect 412692 552 412698 564
rect 417142 552 417148 564
rect 417200 552 417206 604
rect 417878 592 417884 604
rect 417839 564 417884 592
rect 417878 552 417884 564
rect 417936 552 417942 604
rect 418614 592 418620 604
rect 418575 564 418620 592
rect 418614 552 418620 564
rect 418672 552 418678 604
rect 419902 592 419908 604
rect 419863 564 419908 592
rect 419902 552 419908 564
rect 419960 552 419966 604
rect 420546 552 420552 604
rect 420604 592 420610 604
rect 428108 592 428136 700
rect 428553 697 428565 700
rect 428599 697 428611 731
rect 428553 691 428611 697
rect 430546 700 441568 728
rect 428366 620 428372 672
rect 428424 660 428430 672
rect 430546 660 430574 700
rect 441540 672 441568 700
rect 431862 660 431868 672
rect 428424 632 430574 660
rect 431823 632 431868 660
rect 428424 620 428430 632
rect 431862 620 431868 632
rect 431920 620 431926 672
rect 434438 660 434444 672
rect 434399 632 434444 660
rect 434438 620 434444 632
rect 434496 620 434502 672
rect 434548 632 441476 660
rect 420604 564 428136 592
rect 420604 552 420610 564
rect 428458 552 428464 604
rect 428516 552 428522 604
rect 428553 595 428611 601
rect 428553 561 428565 595
rect 428599 592 428611 595
rect 433242 592 433248 604
rect 428599 564 433248 592
rect 428599 561 428611 564
rect 428553 555 428611 561
rect 433242 552 433248 564
rect 433300 552 433306 604
rect 388864 496 397776 524
rect 397825 527 397883 533
rect 388864 484 388870 496
rect 397825 493 397837 527
rect 397871 524 397883 527
rect 407482 524 407488 536
rect 397871 496 407488 524
rect 397871 493 397883 496
rect 397825 487 397883 493
rect 407482 484 407488 496
rect 407540 484 407546 536
rect 413738 524 413744 536
rect 413699 496 413744 524
rect 413738 484 413744 496
rect 413796 484 413802 536
rect 422754 524 422760 536
rect 415366 496 422760 524
rect 380636 428 387794 456
rect 393958 416 393964 468
rect 394016 456 394022 468
rect 394016 428 397868 456
rect 394016 416 394022 428
rect 333606 388 333612 400
rect 329806 360 333612 388
rect 333606 348 333612 360
rect 333664 348 333670 400
rect 336550 348 336556 400
rect 336608 388 336614 400
rect 344738 388 344744 400
rect 336608 360 344744 388
rect 336608 348 336614 360
rect 344738 348 344744 360
rect 344796 348 344802 400
rect 345566 348 345572 400
rect 345624 388 345630 400
rect 355042 388 355048 400
rect 345624 360 355048 388
rect 345624 348 345630 360
rect 355042 348 355048 360
rect 355100 348 355106 400
rect 356974 348 356980 400
rect 357032 388 357038 400
rect 367005 391 367063 397
rect 367005 388 367017 391
rect 357032 360 367017 388
rect 357032 348 357038 360
rect 367005 357 367017 360
rect 367051 357 367063 391
rect 367005 351 367063 357
rect 370406 348 370412 400
rect 370464 388 370470 400
rect 379054 388 379060 400
rect 370464 360 379060 388
rect 370464 348 370470 360
rect 379054 348 379060 360
rect 379112 348 379118 400
rect 381906 348 381912 400
rect 381964 388 381970 400
rect 393222 388 393228 400
rect 381964 360 393228 388
rect 381964 348 381970 360
rect 393222 348 393228 360
rect 393280 348 393286 400
rect 397454 348 397460 400
rect 397512 388 397518 400
rect 397733 391 397791 397
rect 397733 388 397745 391
rect 397512 360 397745 388
rect 397512 348 397518 360
rect 397733 357 397745 360
rect 397779 357 397791 391
rect 397840 388 397868 428
rect 401134 416 401140 468
rect 401192 456 401198 468
rect 412910 456 412916 468
rect 401192 428 412916 456
rect 401192 416 401198 428
rect 412910 416 412916 428
rect 412968 416 412974 468
rect 405826 388 405832 400
rect 397840 360 405832 388
rect 397733 351 397791 357
rect 405826 348 405832 360
rect 405884 348 405890 400
rect 410334 348 410340 400
rect 410392 388 410398 400
rect 415366 388 415394 496
rect 422754 484 422760 496
rect 422812 484 422818 536
rect 416130 416 416136 468
rect 416188 456 416194 468
rect 428476 456 428504 552
rect 429470 484 429476 536
rect 429528 524 429534 536
rect 434548 524 434576 632
rect 435542 592 435548 604
rect 435503 564 435548 592
rect 435542 552 435548 564
rect 435600 552 435606 604
rect 438762 592 438768 604
rect 438723 564 438768 592
rect 438762 552 438768 564
rect 438820 552 438826 604
rect 439130 592 439136 604
rect 439091 564 439136 592
rect 439130 552 439136 564
rect 439188 552 439194 604
rect 440145 595 440203 601
rect 440145 561 440157 595
rect 440191 592 440203 595
rect 440326 592 440332 604
rect 440191 564 440332 592
rect 440191 561 440203 564
rect 440145 555 440203 561
rect 440326 552 440332 564
rect 440384 552 440390 604
rect 441062 592 441068 604
rect 441023 564 441068 592
rect 441062 552 441068 564
rect 441120 552 441126 604
rect 441448 592 441476 632
rect 441522 620 441528 672
rect 441580 620 441586 672
rect 442166 620 442172 672
rect 442224 660 442230 672
rect 443196 660 443224 904
rect 455877 901 455889 904
rect 455923 901 455935 935
rect 466273 935 466331 941
rect 466273 932 466285 935
rect 455877 895 455935 901
rect 465368 904 466285 932
rect 457073 867 457131 873
rect 457073 864 457085 867
rect 445726 836 457085 864
rect 445726 728 445754 836
rect 457073 833 457085 836
rect 457119 833 457131 867
rect 465368 864 465396 904
rect 466273 901 466285 904
rect 466319 901 466331 935
rect 479521 935 479579 941
rect 479521 932 479533 935
rect 466273 895 466331 901
rect 466426 904 479533 932
rect 466426 864 466454 904
rect 479521 901 479533 904
rect 479567 901 479579 935
rect 479521 895 479579 901
rect 480625 935 480683 941
rect 480625 901 480637 935
rect 480671 932 480683 935
rect 492677 935 492735 941
rect 492677 932 492689 935
rect 480671 904 492689 932
rect 480671 901 480683 904
rect 480625 895 480683 901
rect 492677 901 492689 904
rect 492723 901 492735 935
rect 492677 895 492735 901
rect 498933 935 498991 941
rect 498933 901 498945 935
rect 498979 932 498991 935
rect 514941 935 514999 941
rect 514941 932 514953 935
rect 498979 904 514953 932
rect 498979 901 498991 904
rect 498933 895 498991 901
rect 514941 901 514953 904
rect 514987 901 514999 935
rect 514941 895 514999 901
rect 525061 935 525119 941
rect 525061 901 525073 935
rect 525107 932 525119 935
rect 530673 935 530731 941
rect 530673 932 530685 935
rect 525107 904 530685 932
rect 525107 901 525119 904
rect 525061 895 525119 901
rect 530673 901 530685 904
rect 530719 901 530731 935
rect 530673 895 530731 901
rect 538861 935 538919 941
rect 538861 901 538873 935
rect 538907 932 538919 935
rect 538907 904 542354 932
rect 538907 901 538919 904
rect 538861 895 538919 901
rect 457073 827 457131 833
rect 460906 836 465396 864
rect 465460 836 466454 864
rect 481453 867 481511 873
rect 452381 799 452439 805
rect 452381 765 452393 799
rect 452427 796 452439 799
rect 460906 796 460934 836
rect 465460 796 465488 836
rect 481453 833 481465 867
rect 481499 864 481511 867
rect 490469 867 490527 873
rect 490469 864 490481 867
rect 481499 836 490481 864
rect 481499 833 481511 836
rect 481453 827 481511 833
rect 490469 833 490481 836
rect 490515 833 490527 867
rect 498105 867 498163 873
rect 498105 864 498117 867
rect 490469 827 490527 833
rect 490576 836 498117 864
rect 452427 768 460934 796
rect 464724 768 465488 796
rect 465537 799 465595 805
rect 452427 765 452439 768
rect 452381 759 452439 765
rect 454313 731 454371 737
rect 454313 728 454325 731
rect 443288 700 445754 728
rect 449866 700 454325 728
rect 443288 672 443316 700
rect 442224 632 443224 660
rect 442224 620 442230 632
rect 443270 620 443276 672
rect 443328 620 443334 672
rect 445018 660 445024 672
rect 444979 632 445024 660
rect 445018 620 445024 632
rect 445076 620 445082 672
rect 445570 620 445576 672
rect 445628 660 445634 672
rect 449866 660 449894 700
rect 454313 697 454325 700
rect 454359 697 454371 731
rect 454313 691 454371 697
rect 454604 700 458220 728
rect 452378 660 452384 672
rect 445628 632 449894 660
rect 452339 632 452384 660
rect 445628 620 445634 632
rect 452378 620 452384 632
rect 452436 620 452442 672
rect 454405 663 454463 669
rect 454405 629 454417 663
rect 454451 660 454463 663
rect 454494 660 454500 672
rect 454451 632 454500 660
rect 454451 629 454463 632
rect 454405 623 454463 629
rect 454494 620 454500 632
rect 454552 620 454558 672
rect 442626 592 442632 604
rect 441448 564 442632 592
rect 442626 552 442632 564
rect 442684 552 442690 604
rect 444466 552 444472 604
rect 444524 592 444530 604
rect 454604 592 454632 700
rect 458192 672 458220 700
rect 464724 672 464752 768
rect 465537 765 465549 799
rect 465583 796 465595 799
rect 475749 799 475807 805
rect 475749 796 475761 799
rect 465583 768 475761 796
rect 465583 765 465595 768
rect 465537 759 465595 765
rect 475749 765 475761 768
rect 475795 765 475807 799
rect 475749 759 475807 765
rect 475841 799 475899 805
rect 475841 765 475853 799
rect 475887 796 475899 799
rect 489917 799 489975 805
rect 489917 796 489929 799
rect 475887 768 489929 796
rect 475887 765 475899 768
rect 475841 759 475899 765
rect 489917 765 489929 768
rect 489963 765 489975 799
rect 489917 759 489975 765
rect 476761 731 476819 737
rect 476761 697 476773 731
rect 476807 728 476819 731
rect 480717 731 480775 737
rect 480717 728 480729 731
rect 476807 700 480729 728
rect 476807 697 476819 700
rect 476761 691 476819 697
rect 480717 697 480729 700
rect 480763 697 480775 731
rect 480717 691 480775 697
rect 487126 700 488534 728
rect 457070 620 457076 672
rect 457128 660 457134 672
rect 457990 660 457996 672
rect 457128 632 457173 660
rect 457951 632 457996 660
rect 457128 620 457134 632
rect 457990 620 457996 632
rect 458048 620 458054 672
rect 458174 620 458180 672
rect 458232 620 458238 672
rect 459186 660 459192 672
rect 459147 632 459192 660
rect 459186 620 459192 632
rect 459244 620 459250 672
rect 460290 660 460296 672
rect 460251 632 460296 660
rect 460290 620 460296 632
rect 460348 620 460354 672
rect 461946 660 461952 672
rect 461907 632 461952 660
rect 461946 620 461952 632
rect 462004 620 462010 672
rect 464706 620 464712 672
rect 464764 620 464770 672
rect 466270 660 466276 672
rect 466231 632 466276 660
rect 466270 620 466276 632
rect 466328 620 466334 672
rect 466365 663 466423 669
rect 466365 629 466377 663
rect 466411 660 466423 663
rect 472250 660 472256 672
rect 466411 632 472256 660
rect 466411 629 466423 632
rect 466365 623 466423 629
rect 472250 620 472256 632
rect 472308 620 472314 672
rect 472802 660 472808 672
rect 472763 632 472808 660
rect 472802 620 472808 632
rect 472860 620 472866 672
rect 474550 660 474556 672
rect 474511 632 474556 660
rect 474550 620 474556 632
rect 474608 620 474614 672
rect 484026 660 484032 672
rect 474706 632 484032 660
rect 444524 564 454632 592
rect 444524 552 444530 564
rect 455598 552 455604 604
rect 455656 592 455662 604
rect 457533 595 457591 601
rect 457533 592 457545 595
rect 455656 564 457545 592
rect 455656 552 455662 564
rect 457533 561 457545 564
rect 457579 561 457591 595
rect 461486 592 461492 604
rect 457533 555 457591 561
rect 459526 564 461492 592
rect 429528 496 434576 524
rect 429528 484 429534 496
rect 435358 484 435364 536
rect 435416 524 435422 536
rect 448238 524 448244 536
rect 435416 496 448244 524
rect 435416 484 435422 496
rect 448238 484 448244 496
rect 448296 484 448302 536
rect 449618 524 449624 536
rect 449579 496 449624 524
rect 449618 484 449624 496
rect 449676 484 449682 536
rect 452286 524 452292 536
rect 452247 496 452292 524
rect 452286 484 452292 496
rect 452344 484 452350 536
rect 455874 524 455880 536
rect 455835 496 455880 524
rect 455874 484 455880 496
rect 455932 484 455938 536
rect 459526 524 459554 564
rect 461486 552 461492 564
rect 461544 552 461550 604
rect 461762 552 461768 604
rect 461820 592 461826 604
rect 467466 592 467472 604
rect 461820 564 467472 592
rect 461820 552 461826 564
rect 467466 552 467472 564
rect 467524 552 467530 604
rect 468294 592 468300 604
rect 468255 564 468300 592
rect 468294 552 468300 564
rect 468352 552 468358 604
rect 468478 524 468484 536
rect 456168 496 459554 524
rect 461320 496 468484 524
rect 416188 428 428504 456
rect 416188 416 416194 428
rect 430390 416 430396 468
rect 430448 456 430454 468
rect 443638 456 443644 468
rect 430448 428 443644 456
rect 430448 416 430454 428
rect 443638 416 443644 428
rect 443696 416 443702 468
rect 446674 416 446680 468
rect 446732 456 446738 468
rect 456058 456 456064 468
rect 446732 428 456064 456
rect 446732 416 446738 428
rect 456058 416 456064 428
rect 456116 416 456122 468
rect 410392 360 415394 388
rect 410392 348 410398 360
rect 418338 348 418344 400
rect 418396 388 418402 400
rect 430666 388 430672 400
rect 418396 360 430672 388
rect 418396 348 418402 360
rect 430666 348 430672 360
rect 430724 348 430730 400
rect 433058 348 433064 400
rect 433116 388 433122 400
rect 446030 388 446036 400
rect 433116 360 446036 388
rect 433116 348 433122 360
rect 446030 348 446036 360
rect 446088 348 446094 400
rect 447870 348 447876 400
rect 447928 388 447934 400
rect 456168 388 456196 496
rect 447928 360 456196 388
rect 456981 391 457039 397
rect 447928 348 447934 360
rect 456981 357 456993 391
rect 457027 388 457039 391
rect 461320 388 461348 496
rect 468478 484 468484 496
rect 468536 484 468542 536
rect 469214 484 469220 536
rect 469272 524 469278 536
rect 474706 524 474734 632
rect 484026 620 484032 632
rect 484084 620 484090 672
rect 485130 620 485136 672
rect 485188 660 485194 672
rect 487126 660 487154 700
rect 487430 660 487436 672
rect 485188 632 487154 660
rect 487391 632 487436 660
rect 485188 620 485194 632
rect 487430 620 487436 632
rect 487488 620 487494 672
rect 487706 620 487712 672
rect 487764 660 487770 672
rect 488506 660 488534 700
rect 490576 660 490604 836
rect 498105 833 498117 836
rect 498151 833 498163 867
rect 498105 827 498163 833
rect 505741 867 505799 873
rect 505741 833 505753 867
rect 505787 864 505799 867
rect 521841 867 521899 873
rect 521841 864 521853 867
rect 505787 836 521853 864
rect 505787 833 505799 836
rect 505741 827 505799 833
rect 521841 833 521853 836
rect 521887 833 521899 867
rect 521841 827 521899 833
rect 524417 867 524475 873
rect 524417 833 524429 867
rect 524463 864 524475 867
rect 524463 836 540836 864
rect 524463 833 524475 836
rect 524417 827 524475 833
rect 505189 799 505247 805
rect 505189 796 505201 799
rect 492876 768 505201 796
rect 492674 660 492680 672
rect 487764 632 487809 660
rect 488506 632 490604 660
rect 492635 632 492680 660
rect 487764 620 487770 632
rect 492674 620 492680 632
rect 492732 620 492738 672
rect 475746 592 475752 604
rect 475707 564 475752 592
rect 475746 552 475752 564
rect 475804 552 475810 604
rect 479150 592 479156 604
rect 479111 564 479156 592
rect 479150 552 479156 564
rect 479208 552 479214 604
rect 480622 592 480628 604
rect 480583 564 480628 592
rect 480622 552 480628 564
rect 480680 552 480686 604
rect 480806 592 480812 604
rect 480767 564 480812 592
rect 480806 552 480812 564
rect 480864 552 480870 604
rect 480901 595 480959 601
rect 480901 561 480913 595
rect 480947 592 480959 595
rect 485222 592 485228 604
rect 480947 564 485228 592
rect 480947 561 480959 564
rect 480901 555 480959 561
rect 485222 552 485228 564
rect 485280 552 485286 604
rect 486418 592 486424 604
rect 486379 564 486424 592
rect 486418 552 486424 564
rect 486476 552 486482 604
rect 489914 592 489920 604
rect 489875 564 489920 592
rect 489914 552 489920 564
rect 489972 552 489978 604
rect 490469 595 490527 601
rect 490469 561 490481 595
rect 490515 592 490527 595
rect 492582 592 492588 604
rect 490515 564 492588 592
rect 490515 561 490527 564
rect 490469 555 490527 561
rect 492582 552 492588 564
rect 492640 552 492646 604
rect 469272 496 474734 524
rect 469272 484 469278 496
rect 475102 484 475108 536
rect 475160 524 475166 536
rect 475841 527 475899 533
rect 475841 524 475853 527
rect 475160 496 475853 524
rect 475160 484 475166 496
rect 475841 493 475853 496
rect 475887 493 475899 527
rect 475841 487 475899 493
rect 476206 484 476212 536
rect 476264 524 476270 536
rect 481450 524 481456 536
rect 476264 496 478874 524
rect 481411 496 481456 524
rect 476264 484 476270 496
rect 461394 416 461400 468
rect 461452 456 461458 468
rect 465537 459 465595 465
rect 465537 456 465549 459
rect 461452 428 465549 456
rect 461452 416 461458 428
rect 465537 425 465549 428
rect 465583 425 465595 459
rect 465537 419 465595 425
rect 465994 416 466000 468
rect 466052 456 466058 468
rect 476761 459 476819 465
rect 476761 456 476773 459
rect 466052 428 476773 456
rect 466052 416 466058 428
rect 476761 425 476773 428
rect 476807 425 476819 459
rect 478846 456 478874 496
rect 481450 484 481456 496
rect 481508 484 481514 536
rect 483750 524 483756 536
rect 483711 496 483756 524
rect 483750 484 483756 496
rect 483808 484 483814 536
rect 489730 484 489736 536
rect 489788 524 489794 536
rect 492876 524 492904 768
rect 505189 765 505201 768
rect 505235 765 505247 799
rect 505189 759 505247 765
rect 510985 799 511043 805
rect 510985 765 510997 799
rect 511031 796 511043 799
rect 526257 799 526315 805
rect 511031 768 523356 796
rect 511031 765 511043 768
rect 510985 759 511043 765
rect 508869 731 508927 737
rect 508869 728 508881 731
rect 495406 700 508881 728
rect 493318 660 493324 672
rect 493279 632 493324 660
rect 493318 620 493324 632
rect 493376 620 493382 672
rect 494422 620 494428 672
rect 494480 660 494486 672
rect 495406 660 495434 700
rect 508869 697 508881 700
rect 508915 697 508927 731
rect 508869 691 508927 697
rect 508961 731 509019 737
rect 508961 697 508973 731
rect 509007 728 509019 731
rect 509007 700 522988 728
rect 509007 697 509019 700
rect 508961 691 509019 697
rect 505097 663 505155 669
rect 505097 660 505109 663
rect 494480 632 495434 660
rect 495544 632 505109 660
rect 494480 620 494486 632
rect 493502 592 493508 604
rect 493463 564 493508 592
rect 493502 552 493508 564
rect 493560 552 493566 604
rect 494698 592 494704 604
rect 494659 564 494704 592
rect 494698 552 494704 564
rect 494756 552 494762 604
rect 489788 496 492904 524
rect 489788 484 489794 496
rect 478846 428 488534 456
rect 476761 419 476819 425
rect 457027 360 461348 388
rect 461489 391 461547 397
rect 457027 357 457039 360
rect 456981 351 457039 357
rect 461489 357 461501 391
rect 461535 388 461547 391
rect 464982 388 464988 400
rect 461535 360 464988 388
rect 461535 357 461547 360
rect 461489 351 461547 357
rect 464982 348 464988 360
rect 465040 348 465046 400
rect 467190 348 467196 400
rect 467248 388 467254 400
rect 471793 391 471851 397
rect 471793 388 471805 391
rect 467248 360 471805 388
rect 467248 348 467254 360
rect 471793 357 471805 360
rect 471839 357 471851 391
rect 480714 388 480720 400
rect 480675 360 480720 388
rect 471793 351 471851 357
rect 480714 348 480720 360
rect 480772 348 480778 400
rect 488506 388 488534 428
rect 492122 416 492128 468
rect 492180 456 492186 468
rect 495544 456 495572 632
rect 505097 629 505109 632
rect 505143 629 505155 663
rect 505097 623 505155 629
rect 505186 620 505192 672
rect 505244 660 505250 672
rect 505738 660 505744 672
rect 505244 632 505289 660
rect 505699 632 505744 660
rect 505244 620 505250 632
rect 505738 620 505744 632
rect 505796 620 505802 672
rect 507854 620 507860 672
rect 507912 660 507918 672
rect 509881 663 509939 669
rect 507912 632 507957 660
rect 507912 620 507918 632
rect 509881 629 509893 663
rect 509927 660 509939 663
rect 517146 660 517152 672
rect 509927 632 517152 660
rect 509927 629 509939 632
rect 509881 623 509939 629
rect 517146 620 517152 632
rect 517204 620 517210 672
rect 518986 620 518992 672
rect 519044 660 519050 672
rect 520734 660 520740 672
rect 519044 632 519400 660
rect 520695 632 520740 660
rect 519044 620 519050 632
rect 498102 592 498108 604
rect 498063 564 498108 592
rect 498102 552 498108 564
rect 498160 552 498166 604
rect 498194 552 498200 604
rect 498252 592 498258 604
rect 498930 592 498936 604
rect 498252 564 498297 592
rect 498891 564 498936 592
rect 498252 552 498258 564
rect 498930 552 498936 564
rect 498988 552 498994 604
rect 499390 592 499396 604
rect 499351 564 499396 592
rect 499390 552 499396 564
rect 499448 552 499454 604
rect 500126 592 500132 604
rect 500087 564 500132 592
rect 500126 552 500132 564
rect 500184 552 500190 604
rect 502978 592 502984 604
rect 502939 564 502984 592
rect 502978 552 502984 564
rect 503036 552 503042 604
rect 503530 552 503536 604
rect 503588 592 503594 604
rect 519262 592 519268 604
rect 503588 564 519268 592
rect 503588 552 503594 564
rect 519262 552 519268 564
rect 519320 552 519326 604
rect 519372 592 519400 632
rect 520734 620 520740 632
rect 520792 620 520798 672
rect 521838 660 521844 672
rect 521799 632 521844 660
rect 521838 620 521844 632
rect 521896 620 521902 672
rect 522960 660 522988 700
rect 523328 672 523356 768
rect 526257 765 526269 799
rect 526303 796 526315 799
rect 528833 799 528891 805
rect 526303 768 527174 796
rect 526303 765 526315 768
rect 526257 759 526315 765
rect 523420 700 526852 728
rect 523034 660 523040 672
rect 522960 632 523040 660
rect 523034 620 523040 632
rect 523092 620 523098 672
rect 523310 620 523316 672
rect 523368 620 523374 672
rect 523420 592 523448 700
rect 523954 620 523960 672
rect 524012 660 524018 672
rect 524417 663 524475 669
rect 524417 660 524429 663
rect 524012 632 524429 660
rect 524012 620 524018 632
rect 524417 629 524429 632
rect 524463 629 524475 663
rect 526254 660 526260 672
rect 526215 632 526260 660
rect 524417 623 524475 629
rect 526254 620 526260 632
rect 526312 620 526318 672
rect 524230 592 524236 604
rect 519372 564 523448 592
rect 524191 564 524236 592
rect 524230 552 524236 564
rect 524288 552 524294 604
rect 526622 592 526628 604
rect 526583 564 526628 592
rect 526622 552 526628 564
rect 526680 552 526686 604
rect 526824 592 526852 700
rect 527146 660 527174 768
rect 528833 765 528845 799
rect 528879 796 528891 799
rect 532973 799 533031 805
rect 532973 796 532985 799
rect 528879 768 532985 796
rect 528879 765 528891 768
rect 528833 759 528891 765
rect 532973 765 532985 768
rect 533019 765 533031 799
rect 532973 759 533031 765
rect 533065 799 533123 805
rect 533065 765 533077 799
rect 533111 796 533123 799
rect 538861 799 538919 805
rect 538861 796 538873 799
rect 533111 768 538873 796
rect 533111 765 533123 768
rect 533065 759 533123 765
rect 538861 765 538873 768
rect 538907 765 538919 799
rect 538861 759 538919 765
rect 530673 731 530731 737
rect 530673 697 530685 731
rect 530719 728 530731 731
rect 540701 731 540759 737
rect 540701 728 540713 731
rect 530719 700 540713 728
rect 530719 697 530731 700
rect 530673 691 530731 697
rect 540701 697 540713 700
rect 540747 697 540759 731
rect 540701 691 540759 697
rect 533062 660 533068 672
rect 527146 632 531360 660
rect 533023 632 533068 660
rect 528833 595 528891 601
rect 528833 592 528845 595
rect 526824 564 528845 592
rect 528833 561 528845 564
rect 528879 561 528891 595
rect 529014 592 529020 604
rect 528975 564 529020 592
rect 528833 555 528891 561
rect 529014 552 529020 564
rect 529072 552 529078 604
rect 530118 592 530124 604
rect 529124 564 530124 592
rect 497826 484 497832 536
rect 497884 524 497890 536
rect 503901 527 503959 533
rect 503901 524 503913 527
rect 497884 496 503913 524
rect 497884 484 497890 496
rect 503901 493 503913 496
rect 503947 493 503959 527
rect 504634 524 504640 536
rect 504595 496 504640 524
rect 503901 487 503959 493
rect 504634 484 504640 496
rect 504692 484 504698 536
rect 505097 527 505155 533
rect 505097 493 505109 527
rect 505143 524 505155 527
rect 507302 524 507308 536
rect 505143 496 507308 524
rect 505143 493 505155 496
rect 505097 487 505155 493
rect 507302 484 507308 496
rect 507360 484 507366 536
rect 509234 484 509240 536
rect 509292 524 509298 536
rect 512178 524 512184 536
rect 509292 496 512040 524
rect 512139 496 512184 524
rect 509292 484 509298 496
rect 492180 428 495572 456
rect 492180 416 492186 428
rect 501230 416 501236 468
rect 501288 456 501294 468
rect 509881 459 509939 465
rect 509881 456 509893 459
rect 501288 428 509893 456
rect 501288 416 501294 428
rect 509881 425 509893 428
rect 509927 425 509939 459
rect 510338 456 510344 468
rect 510299 428 510344 456
rect 509881 419 509939 425
rect 510338 416 510344 428
rect 510396 416 510402 468
rect 510982 456 510988 468
rect 510943 428 510988 456
rect 510982 416 510988 428
rect 511040 416 511046 468
rect 512012 456 512040 496
rect 512178 484 512184 496
rect 512236 484 512242 536
rect 513742 524 513748 536
rect 513703 496 513748 524
rect 513742 484 513748 496
rect 513800 484 513806 536
rect 514757 527 514815 533
rect 514757 493 514769 527
rect 514803 524 514815 527
rect 525058 524 525064 536
rect 514803 496 524414 524
rect 525019 496 525064 524
rect 514803 493 514815 496
rect 514757 487 514815 493
rect 523218 456 523224 468
rect 512012 428 523224 456
rect 523218 416 523224 428
rect 523276 416 523282 468
rect 524386 456 524414 496
rect 525058 484 525064 496
rect 525116 484 525122 536
rect 529124 456 529152 564
rect 530118 552 530124 564
rect 530176 552 530182 604
rect 531332 524 531360 632
rect 533062 620 533068 632
rect 533120 620 533126 672
rect 533157 663 533215 669
rect 533157 629 533169 663
rect 533203 660 533215 663
rect 535822 660 535828 672
rect 533203 632 535828 660
rect 533203 629 533215 632
rect 533157 623 533215 629
rect 535822 620 535828 632
rect 535880 620 535886 672
rect 540808 604 540836 836
rect 542326 796 542354 904
rect 551189 867 551247 873
rect 551189 833 551201 867
rect 551235 864 551247 867
rect 565814 864 565820 876
rect 551235 836 565820 864
rect 551235 833 551247 836
rect 551189 827 551247 833
rect 565814 824 565820 836
rect 565872 824 565878 876
rect 550269 799 550327 805
rect 550269 796 550281 799
rect 542326 768 550281 796
rect 550269 765 550281 768
rect 550315 765 550327 799
rect 558181 799 558239 805
rect 550269 759 550327 765
rect 553366 768 553808 796
rect 540974 620 540980 672
rect 541032 660 541038 672
rect 553366 660 553394 768
rect 553780 672 553808 768
rect 558181 765 558193 799
rect 558227 796 558239 799
rect 566826 796 566832 808
rect 558227 768 566832 796
rect 558227 765 558239 768
rect 558181 759 558239 765
rect 566826 756 566832 768
rect 566884 756 566890 808
rect 566921 799 566979 805
rect 566921 765 566933 799
rect 566967 796 566979 799
rect 570322 796 570328 808
rect 566967 768 570328 796
rect 566967 765 566979 768
rect 566921 759 566979 765
rect 570322 756 570328 768
rect 570380 756 570386 808
rect 575106 728 575112 740
rect 556908 700 575112 728
rect 556908 672 556936 700
rect 575106 688 575112 700
rect 575164 688 575170 740
rect 541032 632 553394 660
rect 541032 620 541038 632
rect 553762 620 553768 672
rect 553820 620 553826 672
rect 555786 660 555792 672
rect 555747 632 555792 660
rect 555786 620 555792 632
rect 555844 620 555850 672
rect 556890 620 556896 672
rect 556948 620 556954 672
rect 558730 660 558736 672
rect 558691 632 558736 660
rect 558730 620 558736 632
rect 558788 620 558794 672
rect 562594 620 562600 672
rect 562652 660 562658 672
rect 575474 660 575480 672
rect 562652 632 575480 660
rect 562652 620 562658 632
rect 575474 620 575480 632
rect 575532 620 575538 672
rect 531866 552 531872 604
rect 531924 592 531930 604
rect 540609 595 540667 601
rect 540609 592 540621 595
rect 531924 564 540621 592
rect 531924 552 531930 564
rect 540609 561 540621 564
rect 540655 561 540667 595
rect 540609 555 540667 561
rect 540790 552 540796 604
rect 540848 552 540854 604
rect 540885 595 540943 601
rect 540885 561 540897 595
rect 540931 592 540943 595
rect 549070 592 549076 604
rect 540931 564 549076 592
rect 540931 561 540943 564
rect 540885 555 540943 561
rect 549070 552 549076 564
rect 549128 552 549134 604
rect 550266 592 550272 604
rect 550227 564 550272 592
rect 550266 552 550272 564
rect 550324 552 550330 604
rect 551186 592 551192 604
rect 551147 564 551192 592
rect 551186 552 551192 564
rect 551244 552 551250 604
rect 552658 592 552664 604
rect 552619 564 552664 592
rect 552658 552 552664 564
rect 552716 552 552722 604
rect 553026 592 553032 604
rect 552987 564 553032 592
rect 553026 552 553032 564
rect 553084 552 553090 604
rect 553121 595 553179 601
rect 553121 561 553133 595
rect 553167 592 553179 595
rect 568022 592 568028 604
rect 553167 564 568028 592
rect 553167 561 553179 564
rect 553121 555 553179 561
rect 568022 552 568028 564
rect 568080 552 568086 604
rect 543366 524 543372 536
rect 531332 496 543372 524
rect 543366 484 543372 496
rect 543424 484 543430 536
rect 546218 524 546224 536
rect 546179 496 546224 524
rect 546218 484 546224 496
rect 546276 484 546282 536
rect 548886 524 548892 536
rect 548847 496 548892 524
rect 548886 484 548892 496
rect 548944 484 548950 536
rect 550082 484 550088 536
rect 550140 524 550146 536
rect 552937 527 552995 533
rect 552937 524 552949 527
rect 550140 496 552949 524
rect 550140 484 550146 496
rect 552937 493 552949 496
rect 552983 493 552995 527
rect 565446 524 565452 536
rect 552937 487 552995 493
rect 553136 496 565452 524
rect 524386 428 529152 456
rect 529477 459 529535 465
rect 529477 425 529489 459
rect 529523 456 529535 459
rect 533430 456 533436 468
rect 529523 428 533436 456
rect 529523 425 529535 428
rect 529477 419 529535 425
rect 533430 416 533436 428
rect 533488 416 533494 468
rect 534166 416 534172 468
rect 534224 456 534230 468
rect 545666 456 545672 468
rect 534224 428 545672 456
rect 534224 416 534230 428
rect 545666 416 545672 428
rect 545724 416 545730 468
rect 547690 416 547696 468
rect 547748 456 547754 468
rect 553136 456 553164 496
rect 565446 484 565452 496
rect 565504 484 565510 536
rect 563054 456 563060 468
rect 547748 428 553164 456
rect 553228 428 563060 456
rect 547748 416 547754 428
rect 490926 388 490932 400
rect 488506 360 490932 388
rect 490926 348 490932 360
rect 490984 348 490990 400
rect 495342 348 495348 400
rect 495400 388 495406 400
rect 511534 388 511540 400
rect 495400 360 511540 388
rect 495400 348 495406 360
rect 511534 348 511540 360
rect 511592 348 511598 400
rect 513282 348 513288 400
rect 513340 388 513346 400
rect 514757 391 514815 397
rect 514757 388 514769 391
rect 513340 360 514769 388
rect 513340 348 513346 360
rect 514757 357 514769 360
rect 514803 357 514815 391
rect 514938 388 514944 400
rect 514899 360 514944 388
rect 514757 351 514815 357
rect 514938 348 514944 360
rect 514996 348 515002 400
rect 515398 388 515404 400
rect 515359 360 515404 388
rect 515398 348 515404 360
rect 515456 348 515462 400
rect 522850 348 522856 400
rect 522908 388 522914 400
rect 539778 388 539784 400
rect 522908 360 539784 388
rect 522908 348 522914 360
rect 539778 348 539784 360
rect 539836 348 539842 400
rect 540701 391 540759 397
rect 540701 357 540713 391
rect 540747 388 540759 391
rect 542170 388 542176 400
rect 540747 360 542176 388
rect 540747 357 540759 360
rect 540701 351 540759 357
rect 542170 348 542176 360
rect 542228 348 542234 400
rect 542630 348 542636 400
rect 542688 388 542694 400
rect 544194 388 544200 400
rect 542688 360 544200 388
rect 542688 348 542694 360
rect 544194 348 544200 360
rect 544252 348 544258 400
rect 545114 348 545120 400
rect 545172 388 545178 400
rect 553228 388 553256 428
rect 563054 416 563060 428
rect 563112 416 563118 468
rect 545172 360 553256 388
rect 553305 391 553363 397
rect 545172 348 545178 360
rect 553305 357 553317 391
rect 553351 388 553363 391
rect 561766 388 561772 400
rect 553351 360 561772 388
rect 553351 357 553363 360
rect 553305 351 553363 357
rect 561766 348 561772 360
rect 561824 348 561830 400
rect 313700 292 320956 320
rect 321480 292 321554 320
rect 313700 280 313706 292
rect 264882 212 264888 264
rect 264940 252 264946 264
rect 271046 252 271052 264
rect 264940 224 271052 252
rect 264940 212 264946 224
rect 271046 212 271052 224
rect 271104 212 271110 264
rect 282914 212 282920 264
rect 282972 252 282978 264
rect 289998 252 290004 264
rect 282972 224 290004 252
rect 282972 212 282978 224
rect 289998 212 290004 224
rect 290056 212 290062 264
rect 302418 212 302424 264
rect 302476 252 302482 264
rect 310241 255 310299 261
rect 310241 252 310253 255
rect 302476 224 310253 252
rect 302476 212 302482 224
rect 310241 221 310253 224
rect 310287 221 310299 255
rect 310241 215 310299 221
rect 319438 212 319444 264
rect 319496 252 319502 264
rect 321480 252 321508 292
rect 334250 280 334256 332
rect 334308 320 334314 332
rect 343634 320 343640 332
rect 334308 292 343640 320
rect 334308 280 334314 292
rect 343634 280 343640 292
rect 343692 280 343698 332
rect 351270 280 351276 332
rect 351328 320 351334 332
rect 360838 320 360844 332
rect 351328 292 360844 320
rect 351328 280 351334 292
rect 360838 280 360844 292
rect 360896 280 360902 332
rect 362678 280 362684 332
rect 362736 320 362742 332
rect 364978 320 364984 332
rect 362736 292 364984 320
rect 362736 280 362742 292
rect 364978 280 364984 292
rect 365036 280 365042 332
rect 376294 280 376300 332
rect 376352 320 376358 332
rect 386966 320 386972 332
rect 376352 292 386972 320
rect 376352 280 376358 292
rect 386966 280 386972 292
rect 387024 280 387030 332
rect 387610 280 387616 332
rect 387668 320 387674 332
rect 399202 320 399208 332
rect 387668 292 399208 320
rect 387668 280 387674 292
rect 399202 280 399208 292
rect 399260 280 399266 332
rect 399297 323 399355 329
rect 399297 289 399309 323
rect 399343 320 399355 323
rect 401502 320 401508 332
rect 399343 292 401508 320
rect 399343 289 399355 292
rect 399297 283 399355 289
rect 401502 280 401508 292
rect 401560 280 401566 332
rect 402330 280 402336 332
rect 402388 320 402394 332
rect 414014 320 414020 332
rect 402388 292 414020 320
rect 402388 280 402394 292
rect 414014 280 414020 292
rect 414072 280 414078 332
rect 416685 323 416743 329
rect 416685 320 416697 323
rect 414860 292 416697 320
rect 319496 224 321508 252
rect 319496 212 319502 224
rect 321554 212 321560 264
rect 321612 252 321618 264
rect 330110 252 330116 264
rect 321612 224 330116 252
rect 321612 212 321618 224
rect 330110 212 330116 224
rect 330168 212 330174 264
rect 346762 212 346768 264
rect 346820 252 346826 264
rect 356054 252 356060 264
rect 346820 224 356060 252
rect 346820 212 346826 224
rect 356054 212 356060 224
rect 356112 212 356118 264
rect 358078 212 358084 264
rect 358136 252 358142 264
rect 360749 255 360807 261
rect 360749 252 360761 255
rect 358136 224 360761 252
rect 358136 212 358142 224
rect 360749 221 360761 224
rect 360795 221 360807 255
rect 360749 215 360807 221
rect 364886 212 364892 264
rect 364944 252 364950 264
rect 374270 252 374276 264
rect 364944 224 374276 252
rect 364944 212 364950 224
rect 374270 212 374276 224
rect 374328 212 374334 264
rect 375098 212 375104 264
rect 375156 252 375162 264
rect 385957 255 386015 261
rect 385957 252 385969 255
rect 375156 224 385969 252
rect 375156 212 375162 224
rect 385957 221 385969 224
rect 386003 221 386015 255
rect 385957 215 386015 221
rect 386506 212 386512 264
rect 386564 252 386570 264
rect 398006 252 398012 264
rect 386564 224 398012 252
rect 386564 212 386570 224
rect 398006 212 398012 224
rect 398064 212 398070 264
rect 398558 212 398564 264
rect 398616 252 398622 264
rect 410518 252 410524 264
rect 398616 224 410524 252
rect 398616 212 398622 224
rect 410518 212 410524 224
rect 410576 212 410582 264
rect 411530 212 411536 264
rect 411588 252 411594 264
rect 414860 252 414888 292
rect 416685 289 416697 292
rect 416731 289 416743 323
rect 416685 283 416743 289
rect 419442 280 419448 332
rect 419500 320 419506 332
rect 431034 320 431040 332
rect 419500 292 431040 320
rect 419500 280 419506 292
rect 431034 280 431040 292
rect 431092 280 431098 332
rect 434254 280 434260 332
rect 434312 320 434318 332
rect 447134 320 447140 332
rect 434312 292 447140 320
rect 434312 280 434318 292
rect 447134 280 447140 292
rect 447192 280 447198 332
rect 448974 280 448980 332
rect 449032 320 449038 332
rect 449032 292 456104 320
rect 449032 280 449038 292
rect 411588 224 414888 252
rect 411588 212 411594 224
rect 414934 212 414940 264
rect 414992 252 414998 264
rect 427265 255 427323 261
rect 427265 252 427277 255
rect 414992 224 427277 252
rect 414992 212 414998 224
rect 427265 221 427277 224
rect 427311 221 427323 255
rect 427265 215 427323 221
rect 439866 212 439872 264
rect 439924 252 439930 264
rect 453482 252 453488 264
rect 439924 224 453488 252
rect 439924 212 439930 224
rect 453482 212 453488 224
rect 453540 212 453546 264
rect 186958 184 186964 196
rect 184906 156 186964 184
rect 17402 76 17408 128
rect 17460 116 17466 128
rect 20070 116 20076 128
rect 17460 88 20076 116
rect 17460 76 17466 88
rect 20070 76 20076 88
rect 20128 76 20134 128
rect 45738 76 45744 128
rect 45796 116 45802 128
rect 47394 116 47400 128
rect 45796 88 47400 116
rect 45796 76 45802 88
rect 47394 76 47400 88
rect 47452 76 47458 128
rect 129826 76 129832 128
rect 129884 116 129890 128
rect 130286 116 130292 128
rect 129884 88 130292 116
rect 129884 76 129890 88
rect 130286 76 130292 88
rect 130344 76 130350 128
rect 155954 76 155960 128
rect 156012 116 156018 128
rect 157518 116 157524 128
rect 156012 88 157524 116
rect 156012 76 156018 88
rect 157518 76 157524 88
rect 157576 76 157582 128
rect 159358 76 159364 128
rect 159416 116 159422 128
rect 161474 116 161480 128
rect 159416 88 161480 116
rect 159416 76 159422 88
rect 161474 76 161480 88
rect 161532 76 161538 128
rect 184290 76 184296 128
rect 184348 116 184354 128
rect 184906 116 184934 156
rect 186958 144 186964 156
rect 187016 144 187022 196
rect 227346 144 227352 196
rect 227404 184 227410 196
rect 232038 184 232044 196
rect 227404 156 232044 184
rect 227404 144 227410 156
rect 232038 144 232044 156
rect 232096 144 232102 196
rect 257982 144 257988 196
rect 258040 184 258046 196
rect 263870 184 263876 196
rect 258040 156 263876 184
rect 258040 144 258046 156
rect 263870 144 263876 156
rect 263928 144 263934 196
rect 274082 144 274088 196
rect 274140 184 274146 196
rect 280709 187 280767 193
rect 280709 184 280721 187
rect 274140 156 280721 184
rect 274140 144 274146 156
rect 280709 153 280721 156
rect 280755 153 280767 187
rect 280709 147 280767 153
rect 284110 144 284116 196
rect 284168 184 284174 196
rect 291194 184 291200 196
rect 284168 156 291200 184
rect 284168 144 284174 156
rect 291194 144 291200 156
rect 291252 144 291258 196
rect 296806 144 296812 196
rect 296864 184 296870 196
rect 303982 184 303988 196
rect 296864 156 303988 184
rect 296864 144 296870 156
rect 303982 144 303988 156
rect 304040 144 304046 196
rect 320634 144 320640 196
rect 320692 184 320698 196
rect 329006 184 329012 196
rect 320692 156 329012 184
rect 320692 144 320698 156
rect 329006 144 329012 156
rect 329064 144 329070 196
rect 329742 144 329748 196
rect 329800 184 329806 196
rect 338669 187 338727 193
rect 338669 184 338681 187
rect 329800 156 338681 184
rect 329800 144 329806 156
rect 338669 153 338681 156
rect 338715 153 338727 187
rect 338669 147 338727 153
rect 344370 144 344376 196
rect 344428 184 344434 196
rect 352558 184 352564 196
rect 344428 156 352564 184
rect 344428 144 344434 156
rect 352558 144 352564 156
rect 352616 144 352622 196
rect 355870 144 355876 196
rect 355928 184 355934 196
rect 365990 184 365996 196
rect 355928 156 365996 184
rect 355928 144 355934 156
rect 365990 144 365996 156
rect 366048 144 366054 196
rect 367830 144 367836 196
rect 367888 184 367894 196
rect 375466 184 375472 196
rect 367888 156 375472 184
rect 367888 144 367894 156
rect 375466 144 375472 156
rect 375524 144 375530 196
rect 380802 144 380808 196
rect 380860 184 380866 196
rect 391566 184 391572 196
rect 380860 156 391572 184
rect 380860 144 380866 156
rect 391566 144 391572 156
rect 391624 144 391630 196
rect 396258 144 396264 196
rect 396316 184 396322 196
rect 405642 184 405648 196
rect 396316 156 405648 184
rect 396316 144 396322 156
rect 405642 144 405648 156
rect 405700 144 405706 196
rect 406930 144 406936 196
rect 406988 184 406994 196
rect 418798 184 418804 196
rect 406988 156 418804 184
rect 406988 144 406994 156
rect 418798 144 418804 156
rect 418856 144 418862 196
rect 423490 144 423496 196
rect 423548 184 423554 196
rect 436462 184 436468 196
rect 423548 156 436468 184
rect 423548 144 423554 156
rect 436462 144 436468 156
rect 436520 144 436526 196
rect 437474 144 437480 196
rect 437532 184 437538 196
rect 450630 184 450636 196
rect 437532 156 450636 184
rect 437532 144 437538 156
rect 450630 144 450636 156
rect 450688 144 450694 196
rect 456076 184 456104 292
rect 456518 280 456524 332
rect 456576 320 456582 332
rect 470870 320 470876 332
rect 456576 292 470876 320
rect 456576 280 456582 292
rect 470870 280 470876 292
rect 470928 280 470934 332
rect 471698 280 471704 332
rect 471756 320 471762 332
rect 486421 323 486479 329
rect 486421 320 486433 323
rect 471756 292 486433 320
rect 471756 280 471762 292
rect 486421 289 486433 292
rect 486467 289 486479 323
rect 501598 320 501604 332
rect 486421 283 486479 289
rect 490852 292 501604 320
rect 457533 255 457591 261
rect 457533 221 457545 255
rect 457579 252 457591 255
rect 457579 224 461624 252
rect 457579 221 457591 224
rect 457533 215 457591 221
rect 460934 184 460940 196
rect 456076 156 460940 184
rect 460934 144 460940 156
rect 460992 144 460998 196
rect 184348 88 184934 116
rect 184348 76 184354 88
rect 185486 76 185492 128
rect 185544 116 185550 128
rect 188246 116 188252 128
rect 185544 88 188252 116
rect 185544 76 185550 88
rect 188246 76 188252 88
rect 188304 76 188310 128
rect 215018 76 215024 128
rect 215076 116 215082 128
rect 219434 116 219440 128
rect 215076 88 219440 116
rect 215076 76 215082 88
rect 219434 76 219440 88
rect 219492 76 219498 128
rect 228542 76 228548 128
rect 228600 116 228606 128
rect 233234 116 233240 128
rect 228600 88 233240 116
rect 228600 76 228606 88
rect 233234 76 233240 88
rect 233292 76 233298 128
rect 236546 76 236552 128
rect 236604 116 236610 128
rect 241422 116 241428 128
rect 236604 88 241428 116
rect 236604 76 236610 88
rect 241422 76 241428 88
rect 241480 76 241486 128
rect 266078 76 266084 128
rect 266136 116 266142 128
rect 272150 116 272156 128
rect 266136 88 272156 116
rect 266136 76 266142 88
rect 272150 76 272156 88
rect 272208 76 272214 128
rect 299014 76 299020 128
rect 299072 116 299078 128
rect 303798 116 303804 128
rect 299072 88 303804 116
rect 299072 76 299078 88
rect 303798 76 303804 88
rect 303856 76 303862 128
rect 322842 76 322848 128
rect 322900 116 322906 128
rect 331214 116 331220 128
rect 322900 88 331220 116
rect 322900 76 322906 88
rect 331214 76 331220 88
rect 331272 76 331278 128
rect 331950 76 331956 128
rect 332008 116 332014 128
rect 340969 119 341027 125
rect 340969 116 340981 119
rect 332008 88 340981 116
rect 332008 76 332014 88
rect 340969 85 340981 88
rect 341015 85 341027 119
rect 340969 79 341027 85
rect 341794 76 341800 128
rect 341852 116 341858 128
rect 349430 116 349436 128
rect 341852 88 349436 116
rect 341852 76 341858 88
rect 349430 76 349436 88
rect 349488 76 349494 128
rect 357805 119 357863 125
rect 357805 85 357817 119
rect 357851 116 357863 119
rect 363690 116 363696 128
rect 357851 88 363696 116
rect 357851 85 357863 88
rect 357805 79 357863 85
rect 363690 76 363696 88
rect 363748 76 363754 128
rect 366726 76 366732 128
rect 366784 116 366790 128
rect 371881 119 371939 125
rect 371881 116 371893 119
rect 366784 88 371893 116
rect 366784 76 366790 88
rect 371881 85 371893 88
rect 371927 85 371939 119
rect 371881 79 371939 85
rect 385402 76 385408 128
rect 385460 116 385466 128
rect 396810 116 396816 128
rect 385460 88 396816 116
rect 385460 76 385466 88
rect 396810 76 396816 88
rect 396868 76 396874 128
rect 404630 76 404636 128
rect 404688 116 404694 128
rect 416406 116 416412 128
rect 404688 88 416412 116
rect 404688 76 404694 88
rect 416406 76 416412 88
rect 416464 76 416470 128
rect 424686 76 424692 128
rect 424744 116 424750 128
rect 437750 116 437756 128
rect 424744 88 437756 116
rect 424744 76 424750 88
rect 437750 76 437756 88
rect 437808 76 437814 128
rect 451274 76 451280 128
rect 451332 116 451338 128
rect 461489 119 461547 125
rect 461489 116 461501 119
rect 451332 88 461501 116
rect 451332 76 451338 88
rect 461489 85 461501 88
rect 461535 85 461547 119
rect 461596 116 461624 224
rect 462406 212 462412 264
rect 462464 252 462470 264
rect 476758 252 476764 264
rect 462464 224 476764 252
rect 462464 212 462470 224
rect 476758 212 476764 224
rect 476816 212 476822 264
rect 479518 252 479524 264
rect 479479 224 479524 252
rect 479518 212 479524 224
rect 479576 212 479582 264
rect 482646 212 482652 264
rect 482704 252 482710 264
rect 484949 255 485007 261
rect 484949 252 484961 255
rect 482704 224 484961 252
rect 482704 212 482710 224
rect 484949 221 484961 224
rect 484995 221 485007 255
rect 484949 215 485007 221
rect 486050 212 486056 264
rect 486108 252 486114 264
rect 490852 252 490880 292
rect 501598 280 501604 292
rect 501656 280 501662 332
rect 506934 280 506940 332
rect 506992 320 506998 332
rect 508961 323 509019 329
rect 508961 320 508973 323
rect 506992 292 508973 320
rect 506992 280 506998 292
rect 508961 289 508973 292
rect 509007 289 509019 323
rect 508961 283 509019 289
rect 516962 280 516968 332
rect 517020 320 517026 332
rect 529477 323 529535 329
rect 529477 320 529489 323
rect 517020 292 529489 320
rect 517020 280 517026 292
rect 529477 289 529489 292
rect 529523 289 529535 323
rect 529477 283 529535 289
rect 529569 323 529627 329
rect 529569 289 529581 323
rect 529615 320 529627 323
rect 534534 320 534540 332
rect 529615 292 534540 320
rect 529615 289 529627 292
rect 529569 283 529627 289
rect 534534 280 534540 292
rect 534592 280 534598 332
rect 539410 280 539416 332
rect 539468 320 539474 332
rect 557166 320 557172 332
rect 539468 292 557172 320
rect 539468 280 539474 292
rect 557166 280 557172 292
rect 557224 280 557230 332
rect 560202 280 560208 332
rect 560260 320 560266 332
rect 578326 320 578332 332
rect 560260 292 578332 320
rect 560260 280 560266 292
rect 578326 280 578332 292
rect 578384 280 578390 332
rect 486108 224 490880 252
rect 486108 212 486114 224
rect 490926 212 490932 264
rect 490984 252 490990 264
rect 506198 252 506204 264
rect 490984 224 506204 252
rect 490984 212 490990 224
rect 506198 212 506204 224
rect 506256 212 506262 264
rect 508590 252 508596 264
rect 508551 224 508596 252
rect 508590 212 508596 224
rect 508648 212 508654 264
rect 508869 255 508927 261
rect 508869 221 508881 255
rect 508915 252 508927 255
rect 510246 252 510252 264
rect 508915 224 510252 252
rect 508915 221 508927 224
rect 508869 215 508927 221
rect 510246 212 510252 224
rect 510304 212 510310 264
rect 521562 212 521568 264
rect 521620 252 521626 264
rect 538030 252 538036 264
rect 521620 224 538036 252
rect 521620 212 521626 224
rect 538030 212 538036 224
rect 538088 212 538094 264
rect 538766 212 538772 264
rect 538824 252 538830 264
rect 555878 252 555884 264
rect 538824 224 555884 252
rect 538824 212 538830 224
rect 555878 212 555884 224
rect 555936 212 555942 264
rect 557994 212 558000 264
rect 558052 252 558058 264
rect 563790 252 563796 264
rect 558052 224 563796 252
rect 558052 212 558058 224
rect 563790 212 563796 224
rect 563848 212 563854 264
rect 463602 144 463608 196
rect 463660 184 463666 196
rect 477862 184 477868 196
rect 463660 156 477868 184
rect 463660 144 463666 156
rect 477862 144 477868 156
rect 477920 144 477926 196
rect 478506 144 478512 196
rect 478564 184 478570 196
rect 493505 187 493563 193
rect 493505 184 493517 187
rect 478564 156 493517 184
rect 478564 144 478570 156
rect 493505 153 493517 156
rect 493551 153 493563 187
rect 493505 147 493563 153
rect 496722 144 496728 196
rect 496780 184 496786 196
rect 509878 184 509884 196
rect 496780 156 509884 184
rect 496780 144 496786 156
rect 509878 144 509884 156
rect 509936 144 509942 196
rect 518066 184 518072 196
rect 517486 156 518072 184
rect 469582 116 469588 128
rect 461596 88 469588 116
rect 461489 79 461547 85
rect 469582 76 469588 88
rect 469640 76 469646 128
rect 470594 76 470600 128
rect 470652 116 470658 128
rect 482968 125 482974 128
rect 480901 119 480959 125
rect 480901 116 480913 119
rect 470652 88 480913 116
rect 470652 76 470658 88
rect 480901 85 480913 88
rect 480947 85 480959 119
rect 480901 79 480959 85
rect 482925 119 482974 125
rect 482925 85 482937 119
rect 482971 85 482974 119
rect 482925 79 482974 85
rect 482968 76 482974 79
rect 483026 76 483032 128
rect 484949 119 485007 125
rect 484949 85 484961 119
rect 484995 116 485007 119
rect 498197 119 498255 125
rect 498197 116 498209 119
rect 484995 88 498209 116
rect 484995 85 485007 88
rect 484949 79 485007 85
rect 498197 85 498209 88
rect 498243 85 498255 119
rect 498197 79 498255 85
rect 502334 76 502340 128
rect 502392 116 502398 128
rect 517486 116 517514 156
rect 518066 144 518072 156
rect 518124 144 518130 196
rect 520366 144 520372 196
rect 520424 184 520430 196
rect 536926 184 536932 196
rect 520424 156 536932 184
rect 520424 144 520430 156
rect 536926 144 536932 156
rect 536984 144 536990 196
rect 537570 144 537576 196
rect 537628 184 537634 196
rect 543458 184 543464 196
rect 537628 156 543464 184
rect 537628 144 537634 156
rect 543458 144 543464 156
rect 543516 144 543522 196
rect 544194 144 544200 196
rect 544252 184 544258 196
rect 553305 187 553363 193
rect 553305 184 553317 187
rect 544252 156 553317 184
rect 544252 144 544258 156
rect 553305 153 553317 156
rect 553351 153 553363 187
rect 553305 147 553363 153
rect 554590 144 554596 196
rect 554648 184 554654 196
rect 572898 184 572904 196
rect 554648 156 572904 184
rect 554648 144 554654 156
rect 572898 144 572904 156
rect 572956 144 572962 196
rect 502392 88 517514 116
rect 502392 76 502398 88
rect 518158 76 518164 128
rect 518216 116 518222 128
rect 529569 119 529627 125
rect 529569 116 529581 119
rect 518216 88 529581 116
rect 518216 76 518222 88
rect 529569 85 529581 88
rect 529615 85 529627 119
rect 529569 79 529627 85
rect 529658 76 529664 128
rect 529716 116 529722 128
rect 529716 88 533108 116
rect 529716 76 529722 88
rect 16298 8 16304 60
rect 16356 48 16362 60
rect 18966 48 18972 60
rect 16356 20 18972 48
rect 16356 8 16362 20
rect 18966 8 18972 20
rect 19024 8 19030 60
rect 44082 8 44088 60
rect 44140 48 44146 60
rect 46198 48 46204 60
rect 44140 20 46204 48
rect 44140 8 44146 20
rect 46198 8 46204 20
rect 46256 8 46262 60
rect 213822 8 213828 60
rect 213880 48 213886 60
rect 217778 48 217784 60
rect 213880 20 217784 48
rect 213880 8 213886 20
rect 217778 8 217784 20
rect 217836 8 217842 60
rect 241146 8 241152 60
rect 241204 48 241210 60
rect 246022 48 246028 60
rect 241204 20 246028 48
rect 241204 8 241210 20
rect 246022 8 246028 20
rect 246080 8 246086 60
rect 314746 8 314752 60
rect 314804 48 314810 60
rect 322934 48 322940 60
rect 314804 20 322940 48
rect 314804 8 314810 20
rect 322934 8 322940 20
rect 322992 8 322998 60
rect 324038 8 324044 60
rect 324096 48 324102 60
rect 332502 48 332508 60
rect 324096 20 332508 48
rect 324096 8 324102 20
rect 332502 8 332508 20
rect 332560 8 332566 60
rect 333146 8 333152 60
rect 333204 48 333210 60
rect 342346 48 342352 60
rect 333204 20 342352 48
rect 333204 8 333210 20
rect 342346 8 342352 20
rect 342404 8 342410 60
rect 349062 8 349068 60
rect 349120 48 349126 60
rect 358446 48 358452 60
rect 349120 20 358452 48
rect 349120 8 349126 20
rect 358446 8 358452 20
rect 358504 8 358510 60
rect 360749 51 360807 57
rect 360749 17 360761 51
rect 360795 48 360807 51
rect 368201 51 368259 57
rect 368201 48 368213 51
rect 360795 20 368213 48
rect 360795 17 360807 20
rect 360749 11 360807 17
rect 368201 17 368213 20
rect 368247 17 368259 51
rect 368201 11 368259 17
rect 369026 8 369032 60
rect 369084 48 369090 60
rect 376754 48 376760 60
rect 369084 20 376760 48
rect 369084 8 369090 20
rect 376754 8 376760 20
rect 376812 8 376818 60
rect 378594 8 378600 60
rect 378652 48 378658 60
rect 389174 48 389180 60
rect 378652 20 389180 48
rect 378652 8 378658 20
rect 389174 8 389180 20
rect 389232 8 389238 60
rect 389910 8 389916 60
rect 389968 48 389974 60
rect 399297 51 399355 57
rect 399297 48 399309 51
rect 389968 20 399309 48
rect 389968 8 389974 20
rect 399297 17 399309 20
rect 399343 17 399355 51
rect 399297 11 399355 17
rect 399938 8 399944 60
rect 399996 48 400002 60
rect 411622 48 411628 60
rect 399996 20 411628 48
rect 399996 8 400002 20
rect 411622 8 411628 20
rect 411680 8 411686 60
rect 422386 8 422392 60
rect 422444 48 422450 60
rect 435545 51 435603 57
rect 435545 48 435557 51
rect 422444 20 435557 48
rect 422444 8 422450 20
rect 435545 17 435557 20
rect 435591 17 435603 51
rect 435545 11 435603 17
rect 436462 8 436468 60
rect 436520 48 436526 60
rect 449986 48 449992 60
rect 436520 20 449992 48
rect 436520 8 436526 20
rect 449986 8 449992 20
rect 450044 8 450050 60
rect 454218 8 454224 60
rect 454276 48 454282 60
rect 456981 51 457039 57
rect 456981 48 456993 51
rect 454276 20 456993 48
rect 454276 8 454282 20
rect 456981 17 456993 20
rect 457027 17 457039 51
rect 456981 11 457039 17
rect 459002 8 459008 60
rect 459060 48 459066 60
rect 473262 48 473268 60
rect 459060 20 473268 48
rect 459060 8 459066 20
rect 473262 8 473268 20
rect 473320 8 473326 60
rect 473998 8 474004 60
rect 474056 48 474062 60
rect 483566 48 483572 60
rect 474056 20 483572 48
rect 474056 8 474062 20
rect 483566 8 483572 20
rect 483624 8 483630 60
rect 488534 8 488540 60
rect 488592 48 488598 60
rect 503990 48 503996 60
rect 488592 20 503996 48
rect 488592 8 488598 20
rect 503990 8 503996 20
rect 504048 8 504054 60
rect 515582 8 515588 60
rect 515640 48 515646 60
rect 532326 48 532332 60
rect 515640 20 532332 48
rect 515640 8 515646 20
rect 532326 8 532332 20
rect 532384 8 532390 60
rect 533080 48 533108 88
rect 535270 76 535276 128
rect 535328 116 535334 128
rect 552661 119 552719 125
rect 552661 116 552673 119
rect 535328 88 552673 116
rect 535328 76 535334 88
rect 552661 85 552673 88
rect 552707 85 552719 119
rect 552661 79 552719 85
rect 561398 76 561404 128
rect 561456 116 561462 128
rect 580718 116 580724 128
rect 561456 88 580724 116
rect 561456 76 561462 88
rect 580718 76 580724 88
rect 580776 76 580782 128
rect 546494 48 546500 60
rect 533080 20 546500 48
rect 546494 8 546500 20
rect 546552 8 546558 60
rect 552382 8 552388 60
rect 552440 48 552446 60
rect 566921 51 566979 57
rect 566921 48 566933 51
rect 552440 20 566933 48
rect 552440 8 552446 20
rect 566921 17 566933 20
rect 566967 17 566979 51
rect 566921 11 566979 17
<< via1 >>
rect 235448 703808 235500 703860
rect 300860 703808 300912 703860
rect 271788 703740 271840 703792
rect 364708 703740 364760 703792
rect 257252 703672 257304 703724
rect 429476 703672 429528 703724
rect 242440 703604 242492 703656
rect 430028 703604 430080 703656
rect 170496 703536 170548 703588
rect 315488 703536 315540 703588
rect 227628 703468 227680 703520
rect 464436 703468 464488 703520
rect 105452 703400 105504 703452
rect 330300 703400 330352 703452
rect 40500 703332 40552 703384
rect 345020 703332 345072 703384
rect 1492 703264 1544 703316
rect 359740 703264 359792 703316
rect 213000 703196 213052 703248
rect 576400 703196 576452 703248
rect 1584 703128 1636 703180
rect 374460 703128 374512 703180
rect 198280 703060 198332 703112
rect 575020 703060 575072 703112
rect 1676 702992 1728 703044
rect 389180 702992 389232 703044
rect 183376 702924 183428 702976
rect 573640 702924 573692 702976
rect 1768 702856 1820 702908
rect 403900 702856 403952 702908
rect 139308 702788 139360 702840
rect 578976 702788 579028 702840
rect 2596 702720 2648 702772
rect 448152 702720 448204 702772
rect 2228 702652 2280 702704
rect 477592 702652 477644 702704
rect 204 702584 256 702636
rect 507124 702584 507176 702636
rect 20 702516 72 702568
rect 536840 702516 536892 702568
rect 21456 702448 21508 702500
rect 576124 702448 576176 702500
rect 85304 702380 85356 702432
rect 569408 702380 569460 702432
rect 247408 702312 247460 702364
rect 299388 702312 299440 702364
rect 217876 702244 217928 702296
rect 313372 702244 313424 702296
rect 154028 702176 154080 702228
rect 292580 702176 292632 702228
rect 299112 702176 299164 702228
rect 320456 702176 320508 702228
rect 178592 702108 178644 702160
rect 329196 702108 329248 702160
rect 329748 702108 329800 702160
rect 349896 702108 349948 702160
rect 75460 702040 75512 702092
rect 266452 702040 266504 702092
rect 305000 702040 305052 702092
rect 438308 702040 438360 702092
rect 90180 701972 90232 702024
rect 343640 701972 343692 702024
rect 349068 701972 349120 702024
rect 467840 701972 467892 702024
rect 192944 701904 192996 701956
rect 577596 701904 577648 701956
rect 4436 701836 4488 701888
rect 414204 701836 414256 701888
rect 1952 701768 2004 701820
rect 423680 701768 423732 701820
rect 144276 701700 144328 701752
rect 572168 701700 572220 701752
rect 134432 701632 134484 701684
rect 578884 701632 578936 701684
rect 129464 701564 129516 701616
rect 573456 701564 573508 701616
rect 572 701496 624 701548
rect 453028 701496 453080 701548
rect 119712 701428 119764 701480
rect 574836 701428 574888 701480
rect 664 701360 716 701412
rect 458180 701360 458232 701412
rect 2412 701292 2464 701344
rect 472716 701292 472768 701344
rect 104808 701224 104860 701276
rect 577504 701224 577556 701276
rect 480 701156 532 701208
rect 482560 701156 482612 701208
rect 4344 701088 4396 701140
rect 487436 701088 487488 701140
rect 556896 701088 556948 701140
rect 564440 701088 564492 701140
rect 281264 701020 281316 701072
rect 305736 701020 305788 701072
rect 313280 701020 313332 701072
rect 335360 701020 335412 701072
rect 424968 701020 425020 701072
rect 443276 701020 443328 701072
rect 8116 700952 8168 701004
rect 329748 700952 329800 701004
rect 464436 700952 464488 701004
rect 559656 700952 559708 701004
rect 72976 700884 73028 700936
rect 313280 700884 313332 700936
rect 252284 700816 252336 700868
rect 478512 700816 478564 700868
rect 89168 700748 89220 700800
rect 340052 700748 340104 700800
rect 343640 700748 343692 700800
rect 580540 700748 580592 700800
rect 137836 700680 137888 700732
rect 299112 700680 299164 700732
rect 299388 700680 299440 700732
rect 329196 700680 329248 700732
rect 580724 700680 580776 700732
rect 154120 700612 154172 700664
rect 325332 700612 325384 700664
rect 326068 700612 326120 700664
rect 580448 700612 580500 700664
rect 3608 700544 3660 700596
rect 260840 700544 260892 700596
rect 267648 700544 267700 700596
rect 291384 700544 291436 700596
rect 292580 700544 292632 700596
rect 295340 700544 295392 700596
rect 300124 700544 300176 700596
rect 310612 700544 310664 700596
rect 313372 700544 313424 700596
rect 580080 700544 580132 700596
rect 3700 700476 3752 700528
rect 266360 700476 266412 700528
rect 283840 700476 283892 700528
rect 295892 700476 295944 700528
rect 580632 700476 580684 700528
rect 232688 700408 232740 700460
rect 527180 700408 527232 700460
rect 237104 700340 237156 700392
rect 543464 700340 543516 700392
rect 24308 700272 24360 700324
rect 354956 700272 355008 700324
rect 430028 700272 430080 700324
rect 494796 700272 494848 700324
rect 267004 700204 267056 700256
rect 413652 700204 413704 700256
rect 261806 700136 261858 700188
rect 397460 700136 397512 700188
rect 202788 700068 202840 700120
rect 218980 700068 219032 700120
rect 462320 700068 462372 700120
rect 281264 700000 281316 700052
rect 281356 700000 281408 700052
rect 348792 700000 348844 700052
rect 276848 699932 276900 699984
rect 332508 699932 332560 699984
rect 222844 699864 222896 699916
rect 577688 699864 577740 699916
rect 4252 699796 4304 699848
rect 364616 699796 364668 699848
rect 208124 699728 208176 699780
rect 570880 699728 570932 699780
rect 2964 699660 3016 699712
rect 369768 699660 369820 699712
rect 3332 699592 3384 699644
rect 305000 699592 305052 699644
rect 266452 699524 266504 699576
rect 580356 699524 580408 699576
rect 3976 699456 4028 699508
rect 349068 699456 349120 699508
rect 379520 699499 379572 699508
rect 379520 699465 379529 699499
rect 379529 699465 379563 699499
rect 379563 699465 379572 699499
rect 379520 699456 379572 699465
rect 394148 699499 394200 699508
rect 394148 699465 394157 699499
rect 394157 699465 394191 699499
rect 394191 699465 394200 699499
rect 394148 699456 394200 699465
rect 408868 699499 408920 699508
rect 408868 699465 408877 699499
rect 408877 699465 408911 699499
rect 408911 699465 408920 699499
rect 408868 699456 408920 699465
rect 453948 699499 454000 699508
rect 453948 699465 453957 699499
rect 453957 699465 453991 699499
rect 453991 699465 454000 699499
rect 453948 699456 454000 699465
rect 3240 699388 3292 699440
rect 424968 699388 425020 699440
rect 521844 699431 521896 699440
rect 521844 699397 521853 699431
rect 521853 699397 521887 699431
rect 521887 699397 521896 699431
rect 521844 699388 521896 699397
rect 551284 699431 551336 699440
rect 551284 699397 551293 699431
rect 551293 699397 551327 699431
rect 551327 699397 551336 699431
rect 551284 699388 551336 699397
rect 35992 699363 36044 699372
rect 35992 699329 36001 699363
rect 36001 699329 36035 699363
rect 36035 699329 36044 699363
rect 35992 699320 36044 699329
rect 65616 699363 65668 699372
rect 65616 699329 65625 699363
rect 65625 699329 65659 699363
rect 65659 699329 65668 699363
rect 65616 699320 65668 699329
rect 80152 699363 80204 699372
rect 80152 699329 80161 699363
rect 80161 699329 80195 699363
rect 80195 699329 80204 699363
rect 80152 699320 80204 699329
rect 95148 699363 95200 699372
rect 95148 699329 95157 699363
rect 95157 699329 95191 699363
rect 95191 699329 95200 699363
rect 95148 699320 95200 699329
rect 100024 699363 100076 699372
rect 100024 699329 100033 699363
rect 100033 699329 100067 699363
rect 100067 699329 100076 699363
rect 100024 699320 100076 699329
rect 109868 699363 109920 699372
rect 109868 699329 109877 699363
rect 109877 699329 109911 699363
rect 109911 699329 109920 699363
rect 109868 699320 109920 699329
rect 114560 699363 114612 699372
rect 114560 699329 114569 699363
rect 114569 699329 114603 699363
rect 114603 699329 114612 699363
rect 114560 699320 114612 699329
rect 148968 699363 149020 699372
rect 148968 699329 148977 699363
rect 148977 699329 149011 699363
rect 149011 699329 149020 699363
rect 148968 699320 149020 699329
rect 158812 699363 158864 699372
rect 158812 699329 158821 699363
rect 158821 699329 158855 699363
rect 158855 699329 158864 699363
rect 158812 699320 158864 699329
rect 163872 699363 163924 699372
rect 163872 699329 163881 699363
rect 163881 699329 163915 699363
rect 163915 699329 163924 699363
rect 163872 699320 163924 699329
rect 168840 699363 168892 699372
rect 168840 699329 168849 699363
rect 168849 699329 168883 699363
rect 168883 699329 168892 699363
rect 168840 699320 168892 699329
rect 173716 699363 173768 699372
rect 173716 699329 173725 699363
rect 173725 699329 173759 699363
rect 173759 699329 173768 699363
rect 173716 699320 173768 699329
rect 188436 699363 188488 699372
rect 188436 699329 188445 699363
rect 188445 699329 188479 699363
rect 188479 699329 188488 699363
rect 188436 699320 188488 699329
rect 202972 699320 203024 699372
rect 572260 699320 572312 699372
rect 940 699252 992 699304
rect 569592 699184 569644 699236
rect 848 699116 900 699168
rect 565360 699048 565412 699100
rect 573548 698980 573600 699032
rect 756 698912 808 698964
rect 576308 698844 576360 698896
rect 570788 698776 570840 698828
rect 576216 698708 576268 698760
rect 569500 698640 569552 698692
rect 574928 698572 574980 698624
rect 570696 698504 570748 698556
rect 565268 698436 565320 698488
rect 566740 698368 566792 698420
rect 566556 698300 566608 698352
rect 112 697688 164 697740
rect 574744 697620 574796 697672
rect 2044 697552 2096 697604
rect 3424 697484 3476 697536
rect 577688 684428 577740 684480
rect 580816 684428 580868 684480
rect 576400 671984 576452 672036
rect 579620 671984 579672 672036
rect 572260 644376 572312 644428
rect 580172 644376 580224 644428
rect 570880 632000 570932 632052
rect 580172 632000 580224 632052
rect 575020 618196 575072 618248
rect 580172 618196 580224 618248
rect 569592 591948 569644 592000
rect 580172 591948 580224 592000
rect 577596 578144 577648 578196
rect 580816 578144 580868 578196
rect 573640 564340 573692 564392
rect 580172 564340 580224 564392
rect 573548 538160 573600 538212
rect 580172 538160 580224 538212
rect 2780 514836 2832 514888
rect 4436 514836 4488 514888
rect 565360 511912 565412 511964
rect 580172 511912 580224 511964
rect 570788 485732 570840 485784
rect 579620 485732 579672 485784
rect 576308 471928 576360 471980
rect 579804 471928 579856 471980
rect 572168 431876 572220 431928
rect 579712 431876 579764 431928
rect 576216 419432 576268 419484
rect 580172 419432 580224 419484
rect 573456 379448 573508 379500
rect 579620 379448 579672 379500
rect 572076 353200 572128 353252
rect 580172 353200 580224 353252
rect 574928 325592 574980 325644
rect 580172 325592 580224 325644
rect 574836 313216 574888 313268
rect 580172 313216 580224 313268
rect 569500 299412 569552 299464
rect 580172 299412 580224 299464
rect 570696 273164 570748 273216
rect 579620 273164 579672 273216
rect 577504 259360 577556 259412
rect 580632 259360 580684 259412
rect 565268 245556 565320 245608
rect 580172 245556 580224 245608
rect 569408 233180 569460 233232
rect 579988 233180 580040 233232
rect 566740 206932 566792 206984
rect 580172 206932 580224 206984
rect 566556 166948 566608 167000
rect 580172 166948 580224 167000
rect 569316 153144 569368 153196
rect 579804 153144 579856 153196
rect 573364 139340 573416 139392
rect 580172 139340 580224 139392
rect 565176 126896 565228 126948
rect 580172 126896 580224 126948
rect 566648 113092 566700 113144
rect 580172 113092 580224 113144
rect 571984 100648 572036 100700
rect 580172 100648 580224 100700
rect 574744 86912 574796 86964
rect 580172 86912 580224 86964
rect 565084 73108 565136 73160
rect 579988 73108 580040 73160
rect 570604 60664 570656 60716
rect 580172 60664 580224 60716
rect 576124 46860 576176 46912
rect 580172 46860 580224 46912
rect 566464 33056 566516 33108
rect 580172 33056 580224 33108
rect 569224 20612 569276 20664
rect 580172 20612 580224 20664
rect 569132 3068 569184 3120
rect 577412 3068 577464 3120
rect 563704 3000 563756 3052
rect 583392 3000 583444 3052
rect 563520 2932 563572 2984
rect 573916 2932 573968 2984
rect 563796 2864 563848 2916
rect 575480 2864 575532 2916
rect 582196 2864 582248 2916
rect 576308 2796 576360 2848
rect 2964 2048 3016 2100
rect 564440 2048 564492 2100
rect 565820 1368 565872 1420
rect 569040 1368 569092 1420
rect 564440 1232 564492 1284
rect 571524 1164 571576 1216
rect 1676 620 1728 672
rect 5356 620 5408 672
rect 6460 620 6512 672
rect 10048 620 10100 672
rect 572 552 624 604
rect 4344 552 4396 604
rect 5264 552 5316 604
rect 8852 552 8904 604
rect 7472 527 7524 536
rect 7472 493 7481 527
rect 7481 493 7515 527
rect 7515 493 7524 527
rect 7472 484 7524 493
rect 8576 484 8628 536
rect 11152 552 11204 604
rect 11520 620 11572 672
rect 12624 620 12676 672
rect 13360 620 13412 672
rect 16672 620 16724 672
rect 20628 620 20680 672
rect 23480 620 23532 672
rect 12348 552 12400 604
rect 15568 552 15620 604
rect 19432 552 19484 604
rect 22376 552 22428 604
rect 23020 552 23072 604
rect 25780 620 25832 672
rect 28816 620 28868 672
rect 31668 620 31720 672
rect 34796 620 34848 672
rect 37280 620 37332 672
rect 38384 620 38436 672
rect 24860 552 24912 604
rect 25320 552 25372 604
rect 28080 552 28132 604
rect 28724 552 28776 604
rect 29184 552 29236 604
rect 30104 552 30156 604
rect 32588 552 32640 604
rect 37188 552 37240 604
rect 39580 552 39632 604
rect 40684 620 40736 672
rect 42800 620 42852 672
rect 46664 620 46716 672
rect 48504 620 48556 672
rect 48964 620 49016 672
rect 50804 620 50856 672
rect 63224 620 63276 672
rect 40776 552 40828 604
rect 41880 552 41932 604
rect 43996 552 44048 604
rect 47860 552 47912 604
rect 49608 552 49660 604
rect 50160 552 50212 604
rect 51356 552 51408 604
rect 53012 552 53064 604
rect 54944 552 54996 604
rect 56416 552 56468 604
rect 62028 552 62080 604
rect 63316 552 63368 604
rect 64328 620 64380 672
rect 65616 620 65668 672
rect 66720 620 66772 672
rect 68008 620 68060 672
rect 69112 620 69164 672
rect 70584 620 70636 672
rect 133236 620 133288 672
rect 134156 620 134208 672
rect 136180 620 136232 672
rect 137652 620 137704 672
rect 138756 620 138808 672
rect 140044 620 140096 672
rect 151360 620 151412 672
rect 153016 620 153068 672
rect 153660 620 153712 672
rect 155408 620 155460 672
rect 162768 620 162820 672
rect 164884 620 164936 672
rect 64420 552 64472 604
rect 65524 552 65576 604
rect 66812 552 66864 604
rect 70308 552 70360 604
rect 71228 552 71280 604
rect 76196 552 76248 604
rect 76932 552 76984 604
rect 77392 552 77444 604
rect 78036 552 78088 604
rect 78588 552 78640 604
rect 79140 552 79192 604
rect 79692 552 79744 604
rect 80336 552 80388 604
rect 80888 552 80940 604
rect 81440 552 81492 604
rect 82084 552 82136 604
rect 82728 552 82780 604
rect 121828 552 121880 604
rect 122288 552 122340 604
rect 124128 552 124180 604
rect 124680 552 124732 604
rect 125232 552 125284 604
rect 125876 552 125928 604
rect 126428 552 126480 604
rect 126980 552 127032 604
rect 127532 552 127584 604
rect 128176 552 128228 604
rect 128636 552 128688 604
rect 129372 552 129424 604
rect 133880 552 133932 604
rect 135260 552 135312 604
rect 136456 552 136508 604
rect 137560 552 137612 604
rect 138848 552 138900 604
rect 139952 552 140004 604
rect 141240 552 141292 604
rect 144552 552 144604 604
rect 145932 552 145984 604
rect 146852 552 146904 604
rect 148324 552 148376 604
rect 152556 552 152608 604
rect 154212 552 154264 604
rect 154764 552 154816 604
rect 156604 552 156656 604
rect 157064 552 157116 604
rect 158904 552 158956 604
rect 161572 552 161624 604
rect 163688 552 163740 604
rect 14464 484 14516 536
rect 18512 484 18564 536
rect 21272 484 21324 536
rect 22008 484 22060 536
rect 3240 416 3292 468
rect 6644 416 6696 468
rect 24860 416 24912 468
rect 26884 416 26936 468
rect 51908 484 51960 536
rect 67732 484 67784 536
rect 69388 484 69440 536
rect 134984 484 135036 536
rect 141056 484 141108 536
rect 142068 484 142120 536
rect 158168 484 158220 536
rect 159732 484 159784 536
rect 14556 348 14608 400
rect 17868 348 17920 400
rect 42156 416 42208 468
rect 163412 416 163464 468
rect 166080 620 166132 672
rect 167092 620 167144 672
rect 169576 620 169628 672
rect 180892 620 180944 672
rect 183744 620 183796 672
rect 165988 552 166040 604
rect 168380 552 168432 604
rect 170680 552 170732 604
rect 173164 552 173216 604
rect 179788 552 179840 604
rect 182548 552 182600 604
rect 183192 552 183244 604
rect 186136 620 186188 672
rect 191104 620 191156 672
rect 194416 620 194468 672
rect 211620 620 211672 672
rect 215668 620 215720 672
rect 219532 620 219584 672
rect 226156 620 226208 672
rect 231032 620 231084 672
rect 190000 552 190052 604
rect 193220 552 193272 604
rect 196808 552 196860 604
rect 187700 484 187752 536
rect 191012 484 191064 536
rect 192944 484 192996 536
rect 39856 348 39908 400
rect 42892 348 42944 400
rect 45100 348 45152 400
rect 71320 348 71372 400
rect 72332 348 72384 400
rect 72424 348 72476 400
rect 73528 348 73580 400
rect 73620 348 73672 400
rect 74632 348 74684 400
rect 130936 348 130988 400
rect 131948 348 132000 400
rect 132040 348 132092 400
rect 133144 348 133196 400
rect 160468 348 160520 400
rect 162676 348 162728 400
rect 195244 348 195296 400
rect 199108 552 199160 604
rect 203616 552 203668 604
rect 204168 552 204220 604
rect 205732 552 205784 604
rect 209780 552 209832 604
rect 210424 552 210476 604
rect 212172 552 212224 604
rect 214472 552 214524 604
rect 218428 552 218480 604
rect 222752 552 222804 604
rect 223948 552 224000 604
rect 225052 552 225104 604
rect 208400 484 208452 536
rect 225328 484 225380 536
rect 226524 484 226576 536
rect 229836 552 229888 604
rect 229652 484 229704 536
rect 234620 620 234672 672
rect 235448 620 235500 672
rect 237748 620 237800 672
rect 242900 620 242952 672
rect 247960 620 248012 672
rect 253480 620 253532 672
rect 255780 620 255832 672
rect 261760 620 261812 672
rect 262680 620 262732 672
rect 268844 620 268896 672
rect 275836 620 275888 672
rect 277492 620 277544 672
rect 284300 620 284352 672
rect 286600 620 286652 672
rect 288992 620 289044 672
rect 291108 620 291160 672
rect 293408 620 293460 672
rect 231860 552 231912 604
rect 237012 552 237064 604
rect 238116 552 238168 604
rect 233148 484 233200 536
rect 212540 416 212592 468
rect 216588 416 216640 468
rect 221832 416 221884 468
rect 234344 416 234396 468
rect 239312 552 239364 604
rect 240508 595 240560 604
rect 240508 561 240517 595
rect 240517 561 240551 595
rect 240551 561 240560 595
rect 240508 552 240560 561
rect 249984 552 250036 604
rect 251180 595 251232 604
rect 251180 561 251189 595
rect 251189 561 251223 595
rect 251223 561 251232 595
rect 251180 552 251232 561
rect 252284 552 252336 604
rect 244556 484 244608 536
rect 254584 552 254636 604
rect 260656 552 260708 604
rect 258080 484 258132 536
rect 260472 484 260524 536
rect 266544 552 266596 604
rect 267740 552 267792 604
rect 261576 484 261628 536
rect 239956 416 240008 468
rect 244924 416 244976 468
rect 246764 416 246816 468
rect 252560 416 252612 468
rect 259092 416 259144 468
rect 263692 416 263744 468
rect 270040 552 270092 604
rect 271788 552 271840 604
rect 279516 552 279568 604
rect 280712 595 280764 604
rect 280712 561 280721 595
rect 280721 561 280755 595
rect 280755 561 280764 595
rect 280712 552 280764 561
rect 281816 595 281868 604
rect 281816 561 281825 595
rect 281825 561 281859 595
rect 281859 561 281868 595
rect 281816 552 281868 561
rect 283104 595 283156 604
rect 283104 561 283113 595
rect 283113 561 283147 595
rect 283147 561 283156 595
rect 283104 552 283156 561
rect 288808 552 288860 604
rect 296076 552 296128 604
rect 297272 595 297324 604
rect 297272 561 297281 595
rect 297281 561 297315 595
rect 297315 561 297324 595
rect 297272 552 297324 561
rect 298468 620 298520 672
rect 300768 620 300820 672
rect 301320 620 301372 672
rect 307668 663 307720 672
rect 307668 629 307677 663
rect 307677 629 307711 663
rect 307711 629 307720 663
rect 307668 620 307720 629
rect 309048 620 309100 672
rect 311348 620 311400 672
rect 315948 620 316000 672
rect 299664 552 299716 604
rect 268384 484 268436 536
rect 274548 484 274600 536
rect 278504 484 278556 536
rect 270684 416 270736 468
rect 276756 416 276808 468
rect 217232 348 217284 400
rect 221740 348 221792 400
rect 222476 348 222528 400
rect 227260 348 227312 400
rect 245660 348 245712 400
rect 253112 348 253164 400
rect 259276 348 259328 400
rect 264980 348 265032 400
rect 272892 348 272944 400
rect 292212 484 292264 536
rect 280436 416 280488 468
rect 285680 416 285732 468
rect 287612 416 287664 468
rect 293868 416 293920 468
rect 294512 348 294564 400
rect 301964 552 302016 604
rect 308036 552 308088 604
rect 310244 595 310296 604
rect 310244 561 310253 595
rect 310253 561 310287 595
rect 310287 561 310296 595
rect 310244 552 310296 561
rect 311440 595 311492 604
rect 311440 561 311449 595
rect 311449 561 311483 595
rect 311483 561 311492 595
rect 311440 552 311492 561
rect 312636 595 312688 604
rect 312636 561 312645 595
rect 312645 561 312679 595
rect 312679 561 312688 595
rect 312636 552 312688 561
rect 300216 484 300268 536
rect 308772 484 308824 536
rect 317328 552 317380 604
rect 318340 620 318392 672
rect 326804 620 326856 672
rect 327448 620 327500 672
rect 324412 552 324464 604
rect 325608 552 325660 604
rect 326344 552 326396 604
rect 335268 552 335320 604
rect 316040 527 316092 536
rect 316040 493 316049 527
rect 316049 493 316083 527
rect 316083 493 316092 527
rect 316040 484 316092 493
rect 317144 484 317196 536
rect 339776 620 339828 672
rect 336648 552 336700 604
rect 337476 552 337528 604
rect 338672 595 338724 604
rect 338672 561 338681 595
rect 338681 561 338715 595
rect 338715 561 338724 595
rect 338672 552 338724 561
rect 339868 595 339920 604
rect 339868 561 339877 595
rect 339877 561 339911 595
rect 339911 561 339920 595
rect 339868 552 339920 561
rect 340972 595 341024 604
rect 340972 561 340981 595
rect 340981 561 341015 595
rect 341015 561 341024 595
rect 340972 552 341024 561
rect 343180 620 343232 672
rect 352840 620 352892 672
rect 349252 552 349304 604
rect 336464 484 336516 536
rect 337200 484 337252 536
rect 346768 484 346820 536
rect 347688 484 347740 536
rect 357532 552 357584 604
rect 359280 620 359332 672
rect 360384 620 360436 672
rect 363788 620 363840 672
rect 366088 620 366140 672
rect 371608 620 371660 672
rect 373908 620 373960 672
rect 361948 552 362000 604
rect 367008 595 367060 604
rect 367008 561 367017 595
rect 367017 561 367051 595
rect 367051 561 367060 595
rect 367008 552 367060 561
rect 368204 595 368256 604
rect 368204 561 368213 595
rect 368213 561 368247 595
rect 368247 561 368256 595
rect 368204 552 368256 561
rect 369400 595 369452 604
rect 369400 561 369409 595
rect 369409 561 369443 595
rect 369443 561 369452 595
rect 369400 552 369452 561
rect 371700 552 371752 604
rect 376484 552 376536 604
rect 379520 552 379572 604
rect 352472 484 352524 536
rect 354680 484 354732 536
rect 303620 416 303672 468
rect 312452 416 312504 468
rect 320732 416 320784 468
rect 304724 348 304776 400
rect 220176 280 220228 332
rect 243360 280 243412 332
rect 248972 280 249024 332
rect 249708 280 249760 332
rect 255228 280 255280 332
rect 256884 280 256936 332
rect 262772 280 262824 332
rect 279240 280 279292 332
rect 289820 280 289872 332
rect 297916 280 297968 332
rect 305736 280 305788 332
rect 307024 280 307076 332
rect 314844 348 314896 400
rect 318892 348 318944 400
rect 313648 280 313700 332
rect 321836 416 321888 468
rect 325148 416 325200 468
rect 327816 348 327868 400
rect 330852 416 330904 468
rect 340604 416 340656 468
rect 348424 416 348476 468
rect 353576 416 353628 468
rect 361488 484 361540 536
rect 364800 416 364852 468
rect 374368 484 374420 536
rect 377404 484 377456 536
rect 382372 620 382424 672
rect 383108 620 383160 672
rect 390284 620 390336 672
rect 392216 663 392268 672
rect 392216 629 392225 663
rect 392225 629 392259 663
rect 392259 629 392268 663
rect 392216 620 392268 629
rect 394240 620 394292 672
rect 395620 620 395672 672
rect 385960 595 386012 604
rect 385960 561 385969 595
rect 385969 561 386003 595
rect 386003 561 386012 595
rect 385960 552 386012 561
rect 372712 416 372764 468
rect 379612 416 379664 468
rect 382004 484 382056 536
rect 388260 552 388312 604
rect 393320 552 393372 604
rect 388812 484 388864 536
rect 400128 552 400180 604
rect 403072 620 403124 672
rect 403440 620 403492 672
rect 563520 1028 563572 1080
rect 569132 960 569184 1012
rect 404820 552 404872 604
rect 405372 595 405424 604
rect 405372 561 405381 595
rect 405381 561 405415 595
rect 405415 561 405424 595
rect 405372 552 405424 561
rect 407212 620 407264 672
rect 408132 620 408184 672
rect 415492 620 415544 672
rect 409236 595 409288 604
rect 409236 561 409245 595
rect 409245 561 409279 595
rect 409279 561 409288 595
rect 409236 552 409288 561
rect 412640 552 412692 604
rect 421012 620 421064 672
rect 421104 620 421156 672
rect 421748 620 421800 672
rect 426072 620 426124 672
rect 426348 663 426400 672
rect 426348 629 426357 663
rect 426357 629 426391 663
rect 426391 629 426400 663
rect 426992 663 427044 672
rect 426348 620 426400 629
rect 426992 629 427001 663
rect 427001 629 427035 663
rect 427035 629 427044 663
rect 426992 620 427044 629
rect 427268 663 427320 672
rect 427268 629 427277 663
rect 427277 629 427311 663
rect 427311 629 427320 663
rect 427268 620 427320 629
rect 427912 663 427964 672
rect 427912 629 427921 663
rect 427921 629 427955 663
rect 427955 629 427964 663
rect 427912 620 427964 629
rect 417148 595 417200 604
rect 417148 561 417157 595
rect 417157 561 417191 595
rect 417191 561 417200 595
rect 417148 552 417200 561
rect 417884 595 417936 604
rect 417884 561 417893 595
rect 417893 561 417927 595
rect 417927 561 417936 595
rect 417884 552 417936 561
rect 418620 595 418672 604
rect 418620 561 418629 595
rect 418629 561 418663 595
rect 418663 561 418672 595
rect 418620 552 418672 561
rect 419908 595 419960 604
rect 419908 561 419917 595
rect 419917 561 419951 595
rect 419951 561 419960 595
rect 419908 552 419960 561
rect 420552 552 420604 604
rect 428372 620 428424 672
rect 431868 663 431920 672
rect 431868 629 431877 663
rect 431877 629 431911 663
rect 431911 629 431920 663
rect 431868 620 431920 629
rect 434444 663 434496 672
rect 434444 629 434453 663
rect 434453 629 434487 663
rect 434487 629 434496 663
rect 434444 620 434496 629
rect 428464 552 428516 604
rect 433248 552 433300 604
rect 407488 484 407540 536
rect 413744 527 413796 536
rect 413744 493 413753 527
rect 413753 493 413787 527
rect 413787 493 413796 527
rect 413744 484 413796 493
rect 393964 416 394016 468
rect 333612 348 333664 400
rect 336556 348 336608 400
rect 344744 348 344796 400
rect 345572 348 345624 400
rect 355048 348 355100 400
rect 356980 348 357032 400
rect 370412 348 370464 400
rect 379060 348 379112 400
rect 381912 348 381964 400
rect 393228 348 393280 400
rect 397460 348 397512 400
rect 401140 416 401192 468
rect 412916 416 412968 468
rect 405832 348 405884 400
rect 410340 348 410392 400
rect 422760 484 422812 536
rect 416136 416 416188 468
rect 429476 484 429528 536
rect 435548 595 435600 604
rect 435548 561 435557 595
rect 435557 561 435591 595
rect 435591 561 435600 595
rect 435548 552 435600 561
rect 438768 595 438820 604
rect 438768 561 438777 595
rect 438777 561 438811 595
rect 438811 561 438820 595
rect 438768 552 438820 561
rect 439136 595 439188 604
rect 439136 561 439145 595
rect 439145 561 439179 595
rect 439179 561 439188 595
rect 439136 552 439188 561
rect 440332 552 440384 604
rect 441068 595 441120 604
rect 441068 561 441077 595
rect 441077 561 441111 595
rect 441111 561 441120 595
rect 441068 552 441120 561
rect 441528 620 441580 672
rect 442172 620 442224 672
rect 443276 620 443328 672
rect 445024 663 445076 672
rect 445024 629 445033 663
rect 445033 629 445067 663
rect 445067 629 445076 663
rect 445024 620 445076 629
rect 445576 620 445628 672
rect 452384 663 452436 672
rect 452384 629 452393 663
rect 452393 629 452427 663
rect 452427 629 452436 663
rect 452384 620 452436 629
rect 454500 620 454552 672
rect 442632 552 442684 604
rect 444472 552 444524 604
rect 457076 663 457128 672
rect 457076 629 457085 663
rect 457085 629 457119 663
rect 457119 629 457128 663
rect 457996 663 458048 672
rect 457076 620 457128 629
rect 457996 629 458005 663
rect 458005 629 458039 663
rect 458039 629 458048 663
rect 457996 620 458048 629
rect 458180 620 458232 672
rect 459192 663 459244 672
rect 459192 629 459201 663
rect 459201 629 459235 663
rect 459235 629 459244 663
rect 459192 620 459244 629
rect 460296 663 460348 672
rect 460296 629 460305 663
rect 460305 629 460339 663
rect 460339 629 460348 663
rect 460296 620 460348 629
rect 461952 663 462004 672
rect 461952 629 461961 663
rect 461961 629 461995 663
rect 461995 629 462004 663
rect 461952 620 462004 629
rect 464712 620 464764 672
rect 466276 663 466328 672
rect 466276 629 466285 663
rect 466285 629 466319 663
rect 466319 629 466328 663
rect 466276 620 466328 629
rect 472256 620 472308 672
rect 472808 663 472860 672
rect 472808 629 472817 663
rect 472817 629 472851 663
rect 472851 629 472860 663
rect 472808 620 472860 629
rect 474556 663 474608 672
rect 474556 629 474565 663
rect 474565 629 474599 663
rect 474599 629 474608 663
rect 474556 620 474608 629
rect 455604 552 455656 604
rect 435364 484 435416 536
rect 448244 484 448296 536
rect 449624 527 449676 536
rect 449624 493 449633 527
rect 449633 493 449667 527
rect 449667 493 449676 527
rect 449624 484 449676 493
rect 452292 527 452344 536
rect 452292 493 452301 527
rect 452301 493 452335 527
rect 452335 493 452344 527
rect 452292 484 452344 493
rect 455880 527 455932 536
rect 455880 493 455889 527
rect 455889 493 455923 527
rect 455923 493 455932 527
rect 455880 484 455932 493
rect 461492 552 461544 604
rect 461768 552 461820 604
rect 467472 552 467524 604
rect 468300 595 468352 604
rect 468300 561 468309 595
rect 468309 561 468343 595
rect 468343 561 468352 595
rect 468300 552 468352 561
rect 430396 416 430448 468
rect 443644 416 443696 468
rect 446680 416 446732 468
rect 456064 416 456116 468
rect 418344 348 418396 400
rect 430672 348 430724 400
rect 433064 348 433116 400
rect 446036 348 446088 400
rect 447876 348 447928 400
rect 468484 484 468536 536
rect 469220 484 469272 536
rect 484032 620 484084 672
rect 485136 620 485188 672
rect 487436 663 487488 672
rect 487436 629 487445 663
rect 487445 629 487479 663
rect 487479 629 487488 663
rect 487436 620 487488 629
rect 487712 663 487764 672
rect 487712 629 487721 663
rect 487721 629 487755 663
rect 487755 629 487764 663
rect 492680 663 492732 672
rect 487712 620 487764 629
rect 492680 629 492689 663
rect 492689 629 492723 663
rect 492723 629 492732 663
rect 492680 620 492732 629
rect 475752 595 475804 604
rect 475752 561 475761 595
rect 475761 561 475795 595
rect 475795 561 475804 595
rect 475752 552 475804 561
rect 479156 595 479208 604
rect 479156 561 479165 595
rect 479165 561 479199 595
rect 479199 561 479208 595
rect 479156 552 479208 561
rect 480628 595 480680 604
rect 480628 561 480637 595
rect 480637 561 480671 595
rect 480671 561 480680 595
rect 480628 552 480680 561
rect 480812 595 480864 604
rect 480812 561 480821 595
rect 480821 561 480855 595
rect 480855 561 480864 595
rect 480812 552 480864 561
rect 485228 552 485280 604
rect 486424 595 486476 604
rect 486424 561 486433 595
rect 486433 561 486467 595
rect 486467 561 486476 595
rect 486424 552 486476 561
rect 489920 595 489972 604
rect 489920 561 489929 595
rect 489929 561 489963 595
rect 489963 561 489972 595
rect 489920 552 489972 561
rect 492588 552 492640 604
rect 475108 484 475160 536
rect 476212 484 476264 536
rect 481456 527 481508 536
rect 461400 416 461452 468
rect 466000 416 466052 468
rect 481456 493 481465 527
rect 481465 493 481499 527
rect 481499 493 481508 527
rect 481456 484 481508 493
rect 483756 527 483808 536
rect 483756 493 483765 527
rect 483765 493 483799 527
rect 483799 493 483808 527
rect 483756 484 483808 493
rect 489736 484 489788 536
rect 493324 663 493376 672
rect 493324 629 493333 663
rect 493333 629 493367 663
rect 493367 629 493376 663
rect 493324 620 493376 629
rect 494428 620 494480 672
rect 493508 595 493560 604
rect 493508 561 493517 595
rect 493517 561 493551 595
rect 493551 561 493560 595
rect 493508 552 493560 561
rect 494704 595 494756 604
rect 494704 561 494713 595
rect 494713 561 494747 595
rect 494747 561 494756 595
rect 494704 552 494756 561
rect 464988 348 465040 400
rect 467196 348 467248 400
rect 480720 391 480772 400
rect 480720 357 480729 391
rect 480729 357 480763 391
rect 480763 357 480772 391
rect 480720 348 480772 357
rect 492128 416 492180 468
rect 505192 663 505244 672
rect 505192 629 505201 663
rect 505201 629 505235 663
rect 505235 629 505244 663
rect 505744 663 505796 672
rect 505192 620 505244 629
rect 505744 629 505753 663
rect 505753 629 505787 663
rect 505787 629 505796 663
rect 505744 620 505796 629
rect 507860 663 507912 672
rect 507860 629 507869 663
rect 507869 629 507903 663
rect 507903 629 507912 663
rect 507860 620 507912 629
rect 517152 620 517204 672
rect 518992 620 519044 672
rect 520740 663 520792 672
rect 498108 595 498160 604
rect 498108 561 498117 595
rect 498117 561 498151 595
rect 498151 561 498160 595
rect 498108 552 498160 561
rect 498200 595 498252 604
rect 498200 561 498209 595
rect 498209 561 498243 595
rect 498243 561 498252 595
rect 498936 595 498988 604
rect 498200 552 498252 561
rect 498936 561 498945 595
rect 498945 561 498979 595
rect 498979 561 498988 595
rect 498936 552 498988 561
rect 499396 595 499448 604
rect 499396 561 499405 595
rect 499405 561 499439 595
rect 499439 561 499448 595
rect 499396 552 499448 561
rect 500132 595 500184 604
rect 500132 561 500141 595
rect 500141 561 500175 595
rect 500175 561 500184 595
rect 500132 552 500184 561
rect 502984 595 503036 604
rect 502984 561 502993 595
rect 502993 561 503027 595
rect 503027 561 503036 595
rect 502984 552 503036 561
rect 503536 552 503588 604
rect 519268 552 519320 604
rect 520740 629 520749 663
rect 520749 629 520783 663
rect 520783 629 520792 663
rect 520740 620 520792 629
rect 521844 663 521896 672
rect 521844 629 521853 663
rect 521853 629 521887 663
rect 521887 629 521896 663
rect 521844 620 521896 629
rect 523040 620 523092 672
rect 523316 620 523368 672
rect 523960 620 524012 672
rect 526260 663 526312 672
rect 526260 629 526269 663
rect 526269 629 526303 663
rect 526303 629 526312 663
rect 526260 620 526312 629
rect 524236 595 524288 604
rect 524236 561 524245 595
rect 524245 561 524279 595
rect 524279 561 524288 595
rect 524236 552 524288 561
rect 526628 595 526680 604
rect 526628 561 526637 595
rect 526637 561 526671 595
rect 526671 561 526680 595
rect 526628 552 526680 561
rect 533068 663 533120 672
rect 529020 595 529072 604
rect 529020 561 529029 595
rect 529029 561 529063 595
rect 529063 561 529072 595
rect 529020 552 529072 561
rect 497832 484 497884 536
rect 504640 527 504692 536
rect 504640 493 504649 527
rect 504649 493 504683 527
rect 504683 493 504692 527
rect 504640 484 504692 493
rect 507308 484 507360 536
rect 509240 484 509292 536
rect 512184 527 512236 536
rect 501236 416 501288 468
rect 510344 459 510396 468
rect 510344 425 510353 459
rect 510353 425 510387 459
rect 510387 425 510396 459
rect 510344 416 510396 425
rect 510988 459 511040 468
rect 510988 425 510997 459
rect 510997 425 511031 459
rect 511031 425 511040 459
rect 510988 416 511040 425
rect 512184 493 512193 527
rect 512193 493 512227 527
rect 512227 493 512236 527
rect 512184 484 512236 493
rect 513748 527 513800 536
rect 513748 493 513757 527
rect 513757 493 513791 527
rect 513791 493 513800 527
rect 513748 484 513800 493
rect 525064 527 525116 536
rect 523224 416 523276 468
rect 525064 493 525073 527
rect 525073 493 525107 527
rect 525107 493 525116 527
rect 525064 484 525116 493
rect 530124 552 530176 604
rect 533068 629 533077 663
rect 533077 629 533111 663
rect 533111 629 533120 663
rect 533068 620 533120 629
rect 535828 620 535880 672
rect 565820 824 565872 876
rect 540980 620 541032 672
rect 566832 756 566884 808
rect 570328 756 570380 808
rect 575112 688 575164 740
rect 553768 620 553820 672
rect 555792 663 555844 672
rect 555792 629 555801 663
rect 555801 629 555835 663
rect 555835 629 555844 663
rect 555792 620 555844 629
rect 556896 620 556948 672
rect 558736 663 558788 672
rect 558736 629 558745 663
rect 558745 629 558779 663
rect 558779 629 558788 663
rect 558736 620 558788 629
rect 562600 620 562652 672
rect 575480 620 575532 672
rect 531872 552 531924 604
rect 540796 552 540848 604
rect 549076 552 549128 604
rect 550272 595 550324 604
rect 550272 561 550281 595
rect 550281 561 550315 595
rect 550315 561 550324 595
rect 550272 552 550324 561
rect 551192 595 551244 604
rect 551192 561 551201 595
rect 551201 561 551235 595
rect 551235 561 551244 595
rect 551192 552 551244 561
rect 552664 595 552716 604
rect 552664 561 552673 595
rect 552673 561 552707 595
rect 552707 561 552716 595
rect 552664 552 552716 561
rect 553032 595 553084 604
rect 553032 561 553041 595
rect 553041 561 553075 595
rect 553075 561 553084 595
rect 553032 552 553084 561
rect 568028 552 568080 604
rect 543372 484 543424 536
rect 546224 527 546276 536
rect 546224 493 546233 527
rect 546233 493 546267 527
rect 546267 493 546276 527
rect 546224 484 546276 493
rect 548892 527 548944 536
rect 548892 493 548901 527
rect 548901 493 548935 527
rect 548935 493 548944 527
rect 548892 484 548944 493
rect 550088 484 550140 536
rect 533436 416 533488 468
rect 534172 416 534224 468
rect 545672 416 545724 468
rect 547696 416 547748 468
rect 565452 484 565504 536
rect 490932 348 490984 400
rect 495348 348 495400 400
rect 511540 348 511592 400
rect 513288 348 513340 400
rect 514944 391 514996 400
rect 514944 357 514953 391
rect 514953 357 514987 391
rect 514987 357 514996 391
rect 514944 348 514996 357
rect 515404 391 515456 400
rect 515404 357 515413 391
rect 515413 357 515447 391
rect 515447 357 515456 391
rect 515404 348 515456 357
rect 522856 348 522908 400
rect 539784 348 539836 400
rect 542176 348 542228 400
rect 542636 348 542688 400
rect 544200 348 544252 400
rect 545120 348 545172 400
rect 563060 416 563112 468
rect 561772 348 561824 400
rect 264888 212 264940 264
rect 271052 212 271104 264
rect 282920 212 282972 264
rect 290004 212 290056 264
rect 302424 212 302476 264
rect 319444 212 319496 264
rect 334256 280 334308 332
rect 343640 280 343692 332
rect 351276 280 351328 332
rect 360844 280 360896 332
rect 362684 280 362736 332
rect 364984 280 365036 332
rect 376300 280 376352 332
rect 386972 280 387024 332
rect 387616 280 387668 332
rect 399208 280 399260 332
rect 401508 280 401560 332
rect 402336 280 402388 332
rect 414020 280 414072 332
rect 321560 212 321612 264
rect 330116 212 330168 264
rect 346768 212 346820 264
rect 356060 212 356112 264
rect 358084 212 358136 264
rect 364892 212 364944 264
rect 374276 212 374328 264
rect 375104 212 375156 264
rect 386512 212 386564 264
rect 398012 212 398064 264
rect 398564 212 398616 264
rect 410524 212 410576 264
rect 411536 212 411588 264
rect 419448 280 419500 332
rect 431040 280 431092 332
rect 434260 280 434312 332
rect 447140 280 447192 332
rect 448980 280 449032 332
rect 414940 212 414992 264
rect 439872 212 439924 264
rect 453488 212 453540 264
rect 17408 76 17460 128
rect 20076 76 20128 128
rect 45744 76 45796 128
rect 47400 76 47452 128
rect 129832 76 129884 128
rect 130292 76 130344 128
rect 155960 76 156012 128
rect 157524 76 157576 128
rect 159364 76 159416 128
rect 161480 76 161532 128
rect 184296 76 184348 128
rect 186964 144 187016 196
rect 227352 144 227404 196
rect 232044 144 232096 196
rect 257988 144 258040 196
rect 263876 144 263928 196
rect 274088 144 274140 196
rect 284116 144 284168 196
rect 291200 144 291252 196
rect 296812 144 296864 196
rect 303988 144 304040 196
rect 320640 144 320692 196
rect 329012 144 329064 196
rect 329748 144 329800 196
rect 344376 144 344428 196
rect 352564 144 352616 196
rect 355876 144 355928 196
rect 365996 144 366048 196
rect 367836 144 367888 196
rect 375472 144 375524 196
rect 380808 144 380860 196
rect 391572 144 391624 196
rect 396264 144 396316 196
rect 405648 144 405700 196
rect 406936 144 406988 196
rect 418804 144 418856 196
rect 423496 144 423548 196
rect 436468 144 436520 196
rect 437480 144 437532 196
rect 450636 144 450688 196
rect 456524 280 456576 332
rect 470876 280 470928 332
rect 471704 280 471756 332
rect 460940 144 460992 196
rect 185492 76 185544 128
rect 188252 76 188304 128
rect 215024 76 215076 128
rect 219440 76 219492 128
rect 228548 76 228600 128
rect 233240 76 233292 128
rect 236552 76 236604 128
rect 241428 76 241480 128
rect 266084 76 266136 128
rect 272156 76 272208 128
rect 299020 76 299072 128
rect 303804 76 303856 128
rect 322848 76 322900 128
rect 331220 76 331272 128
rect 331956 76 332008 128
rect 341800 76 341852 128
rect 349436 76 349488 128
rect 363696 76 363748 128
rect 366732 76 366784 128
rect 385408 76 385460 128
rect 396816 76 396868 128
rect 404636 76 404688 128
rect 416412 76 416464 128
rect 424692 76 424744 128
rect 437756 76 437808 128
rect 451280 76 451332 128
rect 462412 212 462464 264
rect 476764 212 476816 264
rect 479524 255 479576 264
rect 479524 221 479533 255
rect 479533 221 479567 255
rect 479567 221 479576 255
rect 479524 212 479576 221
rect 482652 212 482704 264
rect 486056 212 486108 264
rect 501604 280 501656 332
rect 506940 280 506992 332
rect 516968 280 517020 332
rect 534540 280 534592 332
rect 539416 280 539468 332
rect 557172 280 557224 332
rect 560208 280 560260 332
rect 578332 280 578384 332
rect 490932 212 490984 264
rect 506204 212 506256 264
rect 508596 255 508648 264
rect 508596 221 508605 255
rect 508605 221 508639 255
rect 508639 221 508648 255
rect 508596 212 508648 221
rect 510252 212 510304 264
rect 521568 212 521620 264
rect 538036 212 538088 264
rect 538772 212 538824 264
rect 555884 212 555936 264
rect 558000 212 558052 264
rect 563796 212 563848 264
rect 463608 144 463660 196
rect 477868 144 477920 196
rect 478512 144 478564 196
rect 496728 144 496780 196
rect 509884 144 509936 196
rect 469588 76 469640 128
rect 470600 76 470652 128
rect 482974 76 483026 128
rect 502340 76 502392 128
rect 518072 144 518124 196
rect 520372 144 520424 196
rect 536932 144 536984 196
rect 537576 144 537628 196
rect 543464 144 543516 196
rect 544200 144 544252 196
rect 554596 144 554648 196
rect 572904 144 572956 196
rect 518164 76 518216 128
rect 529664 76 529716 128
rect 16304 8 16356 60
rect 18972 8 19024 60
rect 44088 8 44140 60
rect 46204 8 46256 60
rect 213828 8 213880 60
rect 217784 8 217836 60
rect 241152 8 241204 60
rect 246028 8 246080 60
rect 314752 8 314804 60
rect 322940 8 322992 60
rect 324044 8 324096 60
rect 332508 8 332560 60
rect 333152 8 333204 60
rect 342352 8 342404 60
rect 349068 8 349120 60
rect 358452 8 358504 60
rect 369032 8 369084 60
rect 376760 8 376812 60
rect 378600 8 378652 60
rect 389180 8 389232 60
rect 389916 8 389968 60
rect 399944 8 399996 60
rect 411628 8 411680 60
rect 422392 8 422444 60
rect 436468 8 436520 60
rect 449992 8 450044 60
rect 454224 8 454276 60
rect 459008 8 459060 60
rect 473268 8 473320 60
rect 474004 8 474056 60
rect 483572 8 483624 60
rect 488540 8 488592 60
rect 503996 8 504048 60
rect 515588 8 515640 60
rect 532332 8 532384 60
rect 535276 76 535328 128
rect 561404 76 561456 128
rect 580724 76 580776 128
rect 546500 8 546552 60
rect 552388 8 552440 60
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 170496 703588 170548 703594
rect 170496 703530 170548 703536
rect 1492 703316 1544 703322
rect 1492 703258 1544 703264
rect 204 702636 256 702642
rect 204 702578 256 702584
rect 20 702568 72 702574
rect 20 702510 72 702516
rect 32 71913 60 702510
rect 112 697740 164 697746
rect 112 697682 164 697688
rect 124 111217 152 697682
rect 216 163441 244 702578
rect 572 701548 624 701554
rect 572 701490 624 701496
rect 294 701448 350 701457
rect 294 701383 350 701392
rect 308 209774 336 701383
rect 480 701208 532 701214
rect 480 701150 532 701156
rect 386 697640 442 697649
rect 386 697575 442 697584
rect 400 229094 428 697575
rect 492 241074 520 701150
rect 584 345409 612 701490
rect 664 701412 716 701418
rect 664 701354 716 701360
rect 676 358465 704 701354
rect 940 699304 992 699310
rect 940 699246 992 699252
rect 848 699168 900 699174
rect 848 699110 900 699116
rect 756 698964 808 698970
rect 756 698906 808 698912
rect 768 501809 796 698906
rect 860 553897 888 699110
rect 952 606121 980 699246
rect 1504 684321 1532 703258
rect 1584 703180 1636 703186
rect 1584 703122 1636 703128
rect 1490 684312 1546 684321
rect 1490 684247 1546 684256
rect 1596 632097 1624 703122
rect 1676 703044 1728 703050
rect 1676 702986 1728 702992
rect 1582 632088 1638 632097
rect 1582 632023 1638 632032
rect 938 606112 994 606121
rect 938 606047 994 606056
rect 1688 580009 1716 702986
rect 1768 702908 1820 702914
rect 1768 702850 1820 702856
rect 1674 580000 1730 580009
rect 1674 579935 1730 579944
rect 846 553888 902 553897
rect 846 553823 902 553832
rect 1780 527921 1808 702850
rect 2596 702772 2648 702778
rect 2596 702714 2648 702720
rect 2228 702704 2280 702710
rect 2228 702646 2280 702652
rect 1952 701820 2004 701826
rect 1952 701762 2004 701768
rect 1858 698184 1914 698193
rect 1858 698119 1914 698128
rect 1766 527912 1822 527921
rect 1766 527847 1822 527856
rect 754 501800 810 501809
rect 754 501735 810 501744
rect 1872 475697 1900 698119
rect 1858 475688 1914 475697
rect 1858 475623 1914 475632
rect 1964 449585 1992 701762
rect 2134 701312 2190 701321
rect 2134 701247 2190 701256
rect 2044 697604 2096 697610
rect 2044 697546 2096 697552
rect 1950 449576 2006 449585
rect 1950 449511 2006 449520
rect 662 358456 718 358465
rect 662 358391 718 358400
rect 570 345400 626 345409
rect 570 345335 626 345344
rect 570 241088 626 241097
rect 492 241046 570 241074
rect 570 241023 626 241032
rect 400 229066 612 229094
rect 584 214985 612 229066
rect 570 214976 626 214985
rect 570 214911 626 214920
rect 308 209746 612 209774
rect 584 201929 612 209746
rect 570 201920 626 201929
rect 570 201855 626 201864
rect 202 163432 258 163441
rect 202 163367 258 163376
rect 110 111208 166 111217
rect 110 111143 166 111152
rect 18 71904 74 71913
rect 18 71839 74 71848
rect 2056 32473 2084 697546
rect 2148 97617 2176 701247
rect 2240 267209 2268 702646
rect 2318 701584 2374 701593
rect 2318 701519 2374 701528
rect 2226 267200 2282 267209
rect 2226 267135 2282 267144
rect 2332 188873 2360 701519
rect 2412 701344 2464 701350
rect 2412 701286 2464 701292
rect 2424 306241 2452 701286
rect 2502 697776 2558 697785
rect 2502 697711 2558 697720
rect 2516 319297 2544 697711
rect 2608 371385 2636 702714
rect 4436 701888 4488 701894
rect 4436 701830 4488 701836
rect 4344 701140 4396 701146
rect 4344 701082 4396 701088
rect 4066 700632 4122 700641
rect 3608 700596 3660 700602
rect 4066 700567 4122 700576
rect 3608 700538 3660 700544
rect 3146 700496 3202 700505
rect 3146 700431 3202 700440
rect 2964 699712 3016 699718
rect 2964 699654 3016 699660
rect 2686 698048 2742 698057
rect 2686 697983 2742 697992
rect 2700 423609 2728 697983
rect 2976 671265 3004 699654
rect 3054 697912 3110 697921
rect 3054 697847 3110 697856
rect 2962 671256 3018 671265
rect 2962 671191 3018 671200
rect 3068 566953 3096 697847
rect 3054 566944 3110 566953
rect 3054 566879 3110 566888
rect 2780 514888 2832 514894
rect 2778 514856 2780 514865
rect 2832 514856 2834 514865
rect 2778 514791 2834 514800
rect 3160 462641 3188 700431
rect 3332 699644 3384 699650
rect 3332 699586 3384 699592
rect 3240 699440 3292 699446
rect 3240 699382 3292 699388
rect 3146 462632 3202 462641
rect 3146 462567 3202 462576
rect 2686 423600 2742 423609
rect 2686 423535 2742 423544
rect 3252 410553 3280 699382
rect 3238 410544 3294 410553
rect 3238 410479 3294 410488
rect 3344 397497 3372 699586
rect 3514 698456 3570 698465
rect 3514 698391 3570 698400
rect 3424 697536 3476 697542
rect 3424 697478 3476 697484
rect 3330 397488 3386 397497
rect 3330 397423 3386 397432
rect 2594 371376 2650 371385
rect 2594 371311 2650 371320
rect 2502 319288 2558 319297
rect 2502 319223 2558 319232
rect 2410 306232 2466 306241
rect 2410 306167 2466 306176
rect 2318 188864 2374 188873
rect 2318 188799 2374 188808
rect 2134 97608 2190 97617
rect 2134 97543 2190 97552
rect 2042 32464 2098 32473
rect 2042 32399 2098 32408
rect 3436 19417 3464 697478
rect 3528 45529 3556 698391
rect 3620 58585 3648 700538
rect 3700 700528 3752 700534
rect 3700 700470 3752 700476
rect 3712 84697 3740 700470
rect 3882 700360 3938 700369
rect 3882 700295 3938 700304
rect 3790 699000 3846 699009
rect 3790 698935 3846 698944
rect 3804 136785 3832 698935
rect 3896 149841 3924 700295
rect 3976 699508 4028 699514
rect 3976 699450 4028 699456
rect 3988 293185 4016 699450
rect 4080 619177 4108 700567
rect 4252 699848 4304 699854
rect 4252 699790 4304 699796
rect 4264 658209 4292 699790
rect 4250 658200 4306 658209
rect 4250 658135 4306 658144
rect 4066 619168 4122 619177
rect 4066 619103 4122 619112
rect 4356 586514 4384 701082
rect 4172 586486 4384 586514
rect 4172 583794 4200 586486
rect 4080 583766 4200 583794
rect 3974 293176 4030 293185
rect 3974 293111 4030 293120
rect 4080 254153 4108 583766
rect 4448 514894 4476 701830
rect 6642 701720 6698 701729
rect 6642 701655 6698 701664
rect 6656 699938 6684 701655
rect 8128 701010 8156 703520
rect 21456 702500 21508 702506
rect 21456 702442 21508 702448
rect 16302 702128 16358 702137
rect 16302 702063 16358 702072
rect 8116 701004 8168 701010
rect 8116 700946 8168 700952
rect 16316 699938 16344 702063
rect 21468 699938 21496 702442
rect 24320 700330 24348 703520
rect 40512 703390 40540 703520
rect 40500 703384 40552 703390
rect 40500 703326 40552 703332
rect 70122 701992 70178 702001
rect 70122 701927 70178 701936
rect 24308 700324 24360 700330
rect 24308 700266 24360 700272
rect 60416 700224 60472 700233
rect 60416 700159 60472 700168
rect 46018 700088 46074 700097
rect 46018 700023 46074 700032
rect 31206 699952 31262 699961
rect 6440 699910 6684 699938
rect 16192 699910 16344 699938
rect 21160 699910 21496 699938
rect 30912 699910 31206 699938
rect 46032 699938 46060 700023
rect 45724 699910 46060 699938
rect 60430 699924 60458 700159
rect 31206 699887 31262 699896
rect 26146 699816 26202 699825
rect 26036 699774 26146 699802
rect 26146 699751 26202 699760
rect 70136 699666 70164 701927
rect 72988 700942 73016 703520
rect 85304 702432 85356 702438
rect 85304 702374 85356 702380
rect 75460 702092 75512 702098
rect 75460 702034 75512 702040
rect 72976 700936 73028 700942
rect 72976 700878 73028 700884
rect 75472 699938 75500 702034
rect 85316 699938 85344 702374
rect 89180 700806 89208 703520
rect 105464 703458 105492 703520
rect 105452 703452 105504 703458
rect 105452 703394 105504 703400
rect 90180 702024 90232 702030
rect 90180 701966 90232 701972
rect 89168 700800 89220 700806
rect 89168 700742 89220 700748
rect 90192 699938 90220 701966
rect 134432 701684 134484 701690
rect 134432 701626 134484 701632
rect 129464 701616 129516 701622
rect 129464 701558 129516 701564
rect 119712 701480 119764 701486
rect 119712 701422 119764 701428
rect 104808 701276 104860 701282
rect 104808 701218 104860 701224
rect 104820 699938 104848 701218
rect 119724 699938 119752 701422
rect 129476 699938 129504 701558
rect 134444 699938 134472 701626
rect 137848 700738 137876 703520
rect 139308 702840 139360 702846
rect 139308 702782 139360 702788
rect 137836 700732 137888 700738
rect 137836 700674 137888 700680
rect 139320 699938 139348 702782
rect 154028 702228 154080 702234
rect 154028 702170 154080 702176
rect 144276 701752 144328 701758
rect 144276 701694 144328 701700
rect 144288 699938 144316 701694
rect 154040 699938 154068 702170
rect 154132 700670 154160 703520
rect 170324 703474 170352 703520
rect 170508 703474 170536 703530
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 227628 703520 227680 703526
rect 235142 703520 235254 704960
rect 235448 703860 235500 703866
rect 235448 703802 235500 703808
rect 235460 703610 235488 703802
rect 235368 703582 235488 703610
rect 242440 703656 242492 703662
rect 242440 703598 242492 703604
rect 170324 703446 170536 703474
rect 198280 703112 198332 703118
rect 198280 703054 198332 703060
rect 183376 702976 183428 702982
rect 183376 702918 183428 702924
rect 178592 702160 178644 702166
rect 178592 702102 178644 702108
rect 154120 700664 154172 700670
rect 154120 700606 154172 700612
rect 178604 699938 178632 702102
rect 183388 699938 183416 702918
rect 192944 701956 192996 701962
rect 192944 701898 192996 701904
rect 75164 699910 75500 699938
rect 85008 699910 85344 699938
rect 89884 699910 90220 699938
rect 104604 699910 104848 699938
rect 119416 699910 119752 699938
rect 129168 699910 129504 699938
rect 134136 699910 134472 699938
rect 139012 699910 139348 699938
rect 143980 699910 144316 699938
rect 153732 699910 154068 699938
rect 178296 699910 178632 699938
rect 183264 699910 183416 699938
rect 192956 699666 192984 701898
rect 198292 699938 198320 703054
rect 202800 700126 202828 703520
rect 213000 703248 213052 703254
rect 213000 703190 213052 703196
rect 202788 700120 202840 700126
rect 202788 700062 202840 700068
rect 213012 699938 213040 703190
rect 217876 702296 217928 702302
rect 217876 702238 217928 702244
rect 217888 699938 217916 702238
rect 218992 700126 219020 703520
rect 227628 703462 227680 703468
rect 235184 703474 235212 703520
rect 235368 703474 235396 703582
rect 218980 700120 219032 700126
rect 218980 700062 219032 700068
rect 227640 699938 227668 703462
rect 235184 703446 235396 703474
rect 232688 700460 232740 700466
rect 232688 700402 232740 700408
rect 232700 699938 232728 700402
rect 237104 700392 237156 700398
rect 237104 700334 237156 700340
rect 197984 699910 198320 699938
rect 212704 699910 213040 699938
rect 217580 699910 217916 699938
rect 222548 699922 222884 699938
rect 222548 699916 222896 699922
rect 222548 699910 222844 699916
rect 227424 699910 227668 699938
rect 232392 699910 232728 699938
rect 222844 699858 222896 699864
rect 207828 699786 208164 699802
rect 207828 699780 208176 699786
rect 207828 699774 208124 699780
rect 208124 699722 208176 699728
rect 237116 699666 237144 700334
rect 242452 699938 242480 703598
rect 251426 703520 251538 704960
rect 257252 703724 257304 703730
rect 257252 703666 257304 703672
rect 247408 702364 247460 702370
rect 247408 702306 247460 702312
rect 247420 699938 247448 702306
rect 252284 700868 252336 700874
rect 252284 700810 252336 700816
rect 252296 699938 252324 700810
rect 257264 699938 257292 703666
rect 267618 703520 267730 704960
rect 271788 703792 271840 703798
rect 271788 703734 271840 703740
rect 266452 702092 266504 702098
rect 266452 702034 266504 702040
rect 266358 701856 266414 701865
rect 266358 701791 266414 701800
rect 260838 701720 260894 701729
rect 260838 701655 260894 701664
rect 260852 700602 260880 701655
rect 260840 700596 260892 700602
rect 260840 700538 260892 700544
rect 266372 700534 266400 701791
rect 266360 700528 266412 700534
rect 266360 700470 266412 700476
rect 261806 700188 261858 700194
rect 261806 700130 261858 700136
rect 242144 699910 242480 699938
rect 247112 699910 247448 699938
rect 251988 699910 252324 699938
rect 256956 699910 257292 699938
rect 261818 699924 261846 700130
rect 70136 699638 70288 699666
rect 192956 699638 193108 699666
rect 237116 699638 237268 699666
rect 266464 699582 266492 702034
rect 267660 700602 267688 703520
rect 267648 700596 267700 700602
rect 267648 700538 267700 700544
rect 267004 700256 267056 700262
rect 267004 700198 267056 700204
rect 267016 699938 267044 700198
rect 271800 699938 271828 703734
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 300860 703860 300912 703866
rect 300860 703802 300912 703808
rect 281264 701072 281316 701078
rect 281264 701014 281316 701020
rect 281276 700058 281304 701014
rect 283852 700534 283880 703520
rect 299388 702364 299440 702370
rect 299388 702306 299440 702312
rect 292580 702228 292632 702234
rect 292580 702170 292632 702176
rect 299112 702228 299164 702234
rect 299112 702170 299164 702176
rect 286690 701176 286746 701185
rect 286690 701111 286746 701120
rect 283840 700528 283892 700534
rect 283840 700470 283892 700476
rect 281264 700052 281316 700058
rect 281264 699994 281316 700000
rect 281356 700052 281408 700058
rect 281356 699994 281408 700000
rect 276848 699984 276900 699990
rect 266708 699910 267044 699938
rect 271676 699910 271828 699938
rect 276552 699932 276848 699938
rect 276552 699926 276900 699932
rect 281368 699938 281396 699994
rect 286704 699938 286732 701111
rect 292592 700602 292620 702170
rect 295338 701176 295394 701185
rect 295338 701111 295394 701120
rect 295352 700602 295380 701111
rect 299124 700738 299152 702170
rect 299400 700738 299428 702306
rect 299112 700732 299164 700738
rect 299112 700674 299164 700680
rect 299388 700732 299440 700738
rect 299388 700674 299440 700680
rect 300136 700602 300164 703520
rect 291384 700596 291436 700602
rect 291384 700538 291436 700544
rect 292580 700596 292632 700602
rect 292580 700538 292632 700544
rect 295340 700596 295392 700602
rect 295340 700538 295392 700544
rect 300124 700596 300176 700602
rect 300124 700538 300176 700544
rect 276552 699910 276888 699926
rect 281368 699910 281520 699938
rect 286396 699910 286732 699938
rect 291396 699666 291424 700538
rect 295892 700528 295944 700534
rect 295892 700470 295944 700476
rect 295904 699938 295932 700470
rect 300872 699938 300900 703802
rect 315488 703588 315540 703594
rect 315488 703530 315540 703536
rect 313372 702296 313424 702302
rect 313372 702238 313424 702244
rect 305000 702092 305052 702098
rect 305000 702034 305052 702040
rect 295904 699910 296240 699938
rect 300872 699910 301116 699938
rect 291272 699638 291424 699666
rect 305012 699650 305040 702034
rect 305736 701072 305788 701078
rect 305736 701014 305788 701020
rect 313280 701072 313332 701078
rect 313280 701014 313332 701020
rect 305748 699938 305776 701014
rect 313292 700942 313320 701014
rect 313280 700936 313332 700942
rect 313280 700878 313332 700884
rect 313384 700602 313412 702238
rect 310612 700596 310664 700602
rect 310612 700538 310664 700544
rect 313372 700596 313424 700602
rect 313372 700538 313424 700544
rect 310624 699938 310652 700538
rect 315500 699938 315528 703530
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364708 703792 364760 703798
rect 364708 703734 364760 703740
rect 364720 703610 364748 703734
rect 364720 703582 364840 703610
rect 330300 703452 330352 703458
rect 330300 703394 330352 703400
rect 320456 702228 320508 702234
rect 320456 702170 320508 702176
rect 320468 699938 320496 702170
rect 329196 702160 329248 702166
rect 329196 702102 329248 702108
rect 329748 702160 329800 702166
rect 329748 702102 329800 702108
rect 326066 701992 326122 702001
rect 326066 701927 326122 701936
rect 326250 701992 326306 702001
rect 326250 701927 326306 701936
rect 326080 700670 326108 701927
rect 325332 700664 325384 700670
rect 325332 700606 325384 700612
rect 326068 700664 326120 700670
rect 326068 700606 326120 700612
rect 325344 699938 325372 700606
rect 305748 699910 306084 699938
rect 310624 699910 310960 699938
rect 315500 699910 315836 699938
rect 320468 699910 320804 699938
rect 325344 699910 325680 699938
rect 305000 699644 305052 699650
rect 305000 699586 305052 699592
rect 266452 699576 266504 699582
rect 266452 699518 266504 699524
rect 326264 699417 326292 701927
rect 329208 700738 329236 702102
rect 329760 701010 329788 702102
rect 329748 701004 329800 701010
rect 329748 700946 329800 700952
rect 329196 700732 329248 700738
rect 329196 700674 329248 700680
rect 330312 699938 330340 703394
rect 332520 699990 332548 703520
rect 345020 703384 345072 703390
rect 345020 703326 345072 703332
rect 343640 702024 343692 702030
rect 343640 701966 343692 701972
rect 335360 701072 335412 701078
rect 335360 701014 335412 701020
rect 332508 699984 332560 699990
rect 330312 699910 330648 699938
rect 332508 699926 332560 699932
rect 335372 699802 335400 701014
rect 343652 700806 343680 701966
rect 340052 700800 340104 700806
rect 340052 700742 340104 700748
rect 343640 700800 343692 700806
rect 343640 700742 343692 700748
rect 340064 699938 340092 700742
rect 345032 699938 345060 703326
rect 348804 700058 348832 703520
rect 364812 703474 364840 703582
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429476 703724 429528 703730
rect 429476 703666 429528 703672
rect 429488 703610 429516 703666
rect 429488 703582 429700 703610
rect 364996 703474 365024 703520
rect 364812 703446 365024 703474
rect 359740 703316 359792 703322
rect 359740 703258 359792 703264
rect 349896 702160 349948 702166
rect 349896 702102 349948 702108
rect 349068 702024 349120 702030
rect 349068 701966 349120 701972
rect 348792 700052 348844 700058
rect 348792 699994 348844 700000
rect 340064 699910 340400 699938
rect 345032 699910 345368 699938
rect 335372 699774 335524 699802
rect 349080 699514 349108 701966
rect 349908 699938 349936 702102
rect 354956 700324 355008 700330
rect 354956 700266 355008 700272
rect 354968 699938 354996 700266
rect 359752 699938 359780 703258
rect 374460 703180 374512 703186
rect 374460 703122 374512 703128
rect 374472 699938 374500 703122
rect 389180 703044 389232 703050
rect 389180 702986 389232 702992
rect 384302 700632 384358 700641
rect 384302 700567 384358 700576
rect 384316 699938 384344 700567
rect 389192 699938 389220 702986
rect 397472 700194 397500 703520
rect 403900 702908 403952 702914
rect 403900 702850 403952 702856
rect 399022 701992 399078 702001
rect 399022 701927 399078 701936
rect 397460 700188 397512 700194
rect 397460 700130 397512 700136
rect 399036 699938 399064 701927
rect 403912 699938 403940 702850
rect 413664 700262 413692 703520
rect 429672 703474 429700 703582
rect 429814 703520 429926 704960
rect 430028 703656 430080 703662
rect 430028 703598 430080 703604
rect 429856 703474 429884 703520
rect 429672 703446 429884 703474
rect 414204 701888 414256 701894
rect 414204 701830 414256 701836
rect 413652 700256 413704 700262
rect 413652 700198 413704 700204
rect 349908 699910 350244 699938
rect 354968 699910 355212 699938
rect 359752 699910 360088 699938
rect 374472 699910 374808 699938
rect 384316 699910 384652 699938
rect 389192 699910 389528 699938
rect 399036 699910 399372 699938
rect 403912 699910 404248 699938
rect 364616 699848 364668 699854
rect 364668 699796 364964 699802
rect 364616 699790 364964 699796
rect 364628 699774 364964 699790
rect 369768 699712 369820 699718
rect 414216 699666 414244 701830
rect 423680 701820 423732 701826
rect 423680 701762 423732 701768
rect 423692 699938 423720 701762
rect 424968 701072 425020 701078
rect 424968 701014 425020 701020
rect 423692 699910 423936 699938
rect 369820 699660 369932 699666
rect 369768 699654 369932 699660
rect 369780 699638 369932 699654
rect 414092 699638 414244 699666
rect 379532 699514 379776 699530
rect 394160 699514 394496 699530
rect 408880 699514 409216 699530
rect 349068 699508 349120 699514
rect 349068 699450 349120 699456
rect 379520 699508 379776 699514
rect 379572 699502 379776 699508
rect 394148 699508 394496 699514
rect 379520 699450 379572 699456
rect 394200 699502 394496 699508
rect 408868 699508 409216 699514
rect 394148 699450 394200 699456
rect 408920 699502 409216 699508
rect 408868 699450 408920 699456
rect 424980 699446 425008 701014
rect 428462 700496 428518 700505
rect 428462 700431 428518 700440
rect 428476 699938 428504 700431
rect 430040 700330 430068 703598
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 464436 703520 464488 703526
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 448152 702772 448204 702778
rect 448152 702714 448204 702720
rect 438308 702092 438360 702098
rect 438308 702034 438360 702040
rect 430028 700324 430080 700330
rect 430028 700266 430080 700272
rect 438320 699938 438348 702034
rect 443276 701072 443328 701078
rect 443276 701014 443328 701020
rect 443288 699938 443316 701014
rect 448164 699938 448192 702714
rect 453028 701548 453080 701554
rect 453028 701490 453080 701496
rect 453040 699938 453068 701490
rect 458180 701412 458232 701418
rect 458180 701354 458232 701360
rect 458192 699938 458220 701354
rect 462332 700126 462360 703520
rect 464436 703462 464488 703468
rect 464448 701010 464476 703462
rect 477592 702704 477644 702710
rect 477592 702646 477644 702652
rect 467840 702024 467892 702030
rect 467840 701966 467892 701972
rect 464436 701004 464488 701010
rect 464436 700946 464488 700952
rect 462320 700120 462372 700126
rect 462320 700062 462372 700068
rect 467852 699938 467880 701966
rect 472716 701344 472768 701350
rect 472716 701286 472768 701292
rect 472728 699938 472756 701286
rect 477604 699938 477632 702646
rect 478524 700874 478552 703520
rect 482560 701208 482612 701214
rect 482560 701150 482612 701156
rect 478512 700868 478564 700874
rect 478512 700810 478564 700816
rect 482572 699938 482600 701150
rect 487436 701140 487488 701146
rect 487436 701082 487488 701088
rect 487448 699938 487476 701082
rect 494808 700330 494836 703520
rect 507124 702636 507176 702642
rect 507124 702578 507176 702584
rect 497278 701584 497334 701593
rect 497278 701519 497334 701528
rect 494796 700324 494848 700330
rect 494796 700266 494848 700272
rect 497292 699938 497320 701519
rect 502338 701448 502394 701457
rect 502338 701383 502394 701392
rect 502352 699938 502380 701383
rect 507136 699938 507164 702578
rect 526718 701856 526774 701865
rect 526718 701791 526774 701800
rect 516966 700360 517022 700369
rect 516966 700295 517022 700304
rect 516980 699938 517008 700295
rect 526732 699938 526760 701791
rect 527192 700466 527220 703520
rect 536840 702568 536892 702574
rect 536840 702510 536892 702516
rect 531686 701312 531742 701321
rect 531686 701247 531742 701256
rect 527180 700460 527232 700466
rect 527180 700402 527232 700408
rect 531700 699938 531728 701247
rect 536852 700210 536880 702510
rect 543476 700398 543504 703520
rect 546498 701720 546554 701729
rect 546498 701655 546554 701664
rect 543464 700392 543516 700398
rect 543464 700334 543516 700340
rect 536852 700182 536926 700210
rect 428476 699910 428812 699938
rect 438320 699910 438656 699938
rect 443288 699910 443624 699938
rect 448164 699910 448500 699938
rect 453040 699910 453376 699938
rect 458192 699910 458344 699938
rect 467852 699910 468188 699938
rect 472728 699910 473064 699938
rect 477604 699910 477940 699938
rect 482572 699910 482908 699938
rect 487448 699910 487784 699938
rect 497292 699910 497628 699938
rect 502352 699910 502504 699938
rect 507136 699910 507472 699938
rect 516980 699910 517316 699938
rect 526732 699910 527068 699938
rect 531700 699910 532036 699938
rect 536898 699924 536926 700182
rect 546512 699938 546540 701655
rect 556896 701140 556948 701146
rect 556896 701082 556948 701088
rect 556908 699938 556936 701082
rect 559668 701010 559696 703520
rect 576400 703248 576452 703254
rect 576400 703190 576452 703196
rect 575020 703112 575072 703118
rect 575020 703054 575072 703060
rect 573640 702976 573692 702982
rect 573640 702918 573692 702924
rect 569408 702432 569460 702438
rect 569408 702374 569460 702380
rect 569222 702128 569278 702137
rect 569222 702063 569278 702072
rect 561126 701992 561182 702001
rect 561126 701927 561182 701936
rect 559656 701004 559708 701010
rect 559656 700946 559708 700952
rect 546512 699910 546756 699938
rect 556600 699910 556936 699938
rect 561140 699938 561168 701927
rect 564440 701140 564492 701146
rect 564440 701082 564492 701088
rect 561140 699910 561476 699938
rect 453946 699544 454002 699553
rect 453946 699479 453948 699488
rect 454000 699479 454002 699488
rect 453948 699450 454000 699456
rect 424968 699440 425020 699446
rect 11610 699408 11666 699417
rect 11316 699366 11610 699394
rect 41050 699408 41106 699417
rect 35880 699378 36032 699394
rect 35880 699372 36044 699378
rect 35880 699366 35992 699372
rect 11610 699343 11666 699352
rect 40756 699366 41050 699394
rect 50894 699408 50950 699417
rect 50600 699366 50894 699394
rect 41050 699343 41106 699352
rect 55770 699408 55826 699417
rect 55476 699366 55770 699394
rect 50894 699343 50950 699352
rect 124586 699408 124642 699417
rect 65320 699378 65656 699394
rect 80040 699378 80192 699394
rect 94852 699378 95188 699394
rect 99728 699378 100064 699394
rect 109572 699378 109908 699394
rect 114448 699378 114600 699394
rect 65320 699372 65668 699378
rect 65320 699366 65616 699372
rect 55770 699343 55826 699352
rect 35992 699314 36044 699320
rect 80040 699372 80204 699378
rect 80040 699366 80152 699372
rect 65616 699314 65668 699320
rect 94852 699372 95200 699378
rect 94852 699366 95148 699372
rect 80152 699314 80204 699320
rect 99728 699372 100076 699378
rect 99728 699366 100024 699372
rect 95148 699314 95200 699320
rect 109572 699372 109920 699378
rect 109572 699366 109868 699372
rect 100024 699314 100076 699320
rect 114448 699372 114612 699378
rect 114448 699366 114560 699372
rect 109868 699314 109920 699320
rect 124292 699366 124586 699394
rect 326250 699408 326306 699417
rect 148856 699378 149008 699394
rect 158700 699378 158852 699394
rect 163576 699378 163912 699394
rect 168544 699378 168880 699394
rect 173420 699378 173756 699394
rect 188140 699378 188476 699394
rect 202860 699378 203012 699394
rect 148856 699372 149020 699378
rect 148856 699366 148968 699372
rect 124586 699343 124642 699352
rect 114560 699314 114612 699320
rect 158700 699372 158864 699378
rect 158700 699366 158812 699372
rect 148968 699314 149020 699320
rect 163576 699372 163924 699378
rect 163576 699366 163872 699372
rect 158812 699314 158864 699320
rect 168544 699372 168892 699378
rect 168544 699366 168840 699372
rect 163872 699314 163924 699320
rect 173420 699372 173768 699378
rect 173420 699366 173716 699372
rect 168840 699314 168892 699320
rect 188140 699372 188488 699378
rect 188140 699366 188436 699372
rect 173716 699314 173768 699320
rect 202860 699372 203024 699378
rect 202860 699366 202972 699372
rect 188436 699314 188488 699320
rect 326250 699343 326306 699352
rect 418710 699408 418766 699417
rect 418766 699366 419060 699394
rect 521844 699440 521896 699446
rect 424968 699382 425020 699388
rect 433430 699408 433486 699417
rect 418710 699343 418766 699352
rect 462870 699408 462926 699417
rect 433486 699366 433780 699394
rect 433430 699343 433486 699352
rect 492586 699408 492642 699417
rect 462926 699366 463220 699394
rect 462870 699343 462926 699352
rect 511998 699408 512054 699417
rect 492642 699366 492752 699394
rect 492586 699343 492642 699352
rect 512054 699366 512348 699394
rect 551284 699440 551336 699446
rect 541530 699408 541586 699417
rect 521896 699388 522192 699394
rect 521844 699382 522192 699388
rect 521856 699366 522192 699382
rect 511998 699343 512054 699352
rect 541586 699366 541880 699394
rect 551336 699388 551632 699394
rect 551284 699382 551632 699388
rect 551296 699366 551632 699382
rect 541530 699343 541586 699352
rect 202972 699314 203024 699320
rect 4436 514888 4488 514894
rect 4436 514830 4488 514836
rect 4066 254144 4122 254153
rect 4066 254079 4122 254088
rect 3882 149832 3938 149841
rect 3882 149767 3938 149776
rect 3790 136776 3846 136785
rect 3790 136711 3846 136720
rect 3698 84688 3754 84697
rect 3698 84623 3754 84632
rect 3606 58576 3662 58585
rect 3606 58511 3662 58520
rect 3514 45520 3570 45529
rect 3514 45455 3570 45464
rect 3422 19408 3478 19417
rect 3422 19343 3478 19352
rect 2962 6488 3018 6497
rect 2962 6423 3018 6432
rect 2976 2106 3004 6423
rect 563704 3052 563756 3058
rect 563704 2994 563756 3000
rect 563520 2984 563572 2990
rect 563520 2926 563572 2932
rect 2964 2100 3016 2106
rect 2964 2042 3016 2048
rect 563532 1086 563560 2926
rect 563520 1080 563572 1086
rect 563520 1022 563572 1028
rect 563716 762 563744 2994
rect 563796 2916 563848 2922
rect 563796 2858 563848 2864
rect 563408 734 563744 762
rect 1676 672 1728 678
rect 5356 672 5408 678
rect 1676 614 1728 620
rect 4066 640 4122 649
rect 572 604 624 610
rect 572 546 624 552
rect 584 480 612 546
rect 1688 480 1716 614
rect 2884 564 3096 592
rect 4356 610 4600 626
rect 6460 672 6512 678
rect 5408 620 5704 626
rect 5356 614 5704 620
rect 10048 672 10100 678
rect 7838 640 7894 649
rect 6460 614 6512 620
rect 4066 575 4122 584
rect 4344 604 4600 610
rect 2884 480 2912 564
rect 3068 490 3096 564
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 3068 474 3280 490
rect 4080 480 4108 575
rect 4396 598 4600 604
rect 5264 604 5316 610
rect 4344 546 4396 552
rect 5368 598 5704 614
rect 5264 546 5316 552
rect 5276 480 5304 546
rect 6472 480 6500 614
rect 7484 598 7696 626
rect 7484 542 7512 598
rect 7472 536 7524 542
rect 3068 468 3292 474
rect 3068 462 3240 468
rect 3240 410 3292 416
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 6656 474 6808 490
rect 7472 478 7524 484
rect 7668 480 7696 598
rect 9954 640 10010 649
rect 7894 598 8004 626
rect 8588 598 8800 626
rect 8864 610 9108 626
rect 7838 575 7894 584
rect 8588 542 8616 598
rect 8576 536 8628 542
rect 6644 468 6808 474
rect 6696 462 6808 468
rect 6644 410 6696 416
rect 7626 -960 7738 480
rect 8576 478 8628 484
rect 8772 480 8800 598
rect 8852 604 9108 610
rect 8904 598 9108 604
rect 11520 672 11572 678
rect 10100 620 10212 626
rect 10048 614 10212 620
rect 10060 598 10212 614
rect 11408 620 11520 626
rect 12624 672 12676 678
rect 11408 614 11572 620
rect 12512 620 12624 626
rect 12512 614 12676 620
rect 13360 672 13412 678
rect 16672 672 16724 678
rect 13726 640 13782 649
rect 13360 614 13412 620
rect 11152 604 11204 610
rect 9954 575 10010 584
rect 8852 546 8904 552
rect 9968 480 9996 575
rect 11408 598 11560 614
rect 12348 604 12400 610
rect 11152 546 11204 552
rect 12512 598 12664 614
rect 12348 546 12400 552
rect 11164 480 11192 546
rect 12360 480 12388 546
rect 8730 -960 8842 480
rect 9926 -960 10038 480
rect 11122 -960 11234 480
rect 12318 -960 12430 480
rect 13372 218 13400 614
rect 13616 598 13726 626
rect 13726 575 13782 584
rect 14476 598 14812 626
rect 15580 610 15916 626
rect 20628 672 20680 678
rect 16724 620 17020 626
rect 16672 614 17020 620
rect 15568 604 15916 610
rect 14476 542 14504 598
rect 15620 598 15916 604
rect 16684 598 17020 614
rect 17880 598 18216 626
rect 23480 672 23532 678
rect 20628 614 20680 620
rect 19432 604 19484 610
rect 15568 546 15620 552
rect 14464 536 14516 542
rect 13514 218 13626 480
rect 14464 478 14516 484
rect 14556 400 14608 406
rect 14710 354 14822 480
rect 14608 348 14822 354
rect 14556 342 14822 348
rect 14568 326 14822 342
rect 13372 190 13626 218
rect 13514 -960 13626 190
rect 14710 -960 14822 326
rect 15906 82 16018 480
rect 17010 82 17122 480
rect 17880 406 17908 598
rect 19432 546 19484 552
rect 18512 536 18564 542
rect 17868 400 17920 406
rect 17868 342 17920 348
rect 18206 218 18318 480
rect 18512 478 18564 484
rect 19444 480 19472 546
rect 20640 480 20668 614
rect 21836 598 22048 626
rect 22388 610 22724 626
rect 25780 672 25832 678
rect 23532 620 23828 626
rect 23480 614 23828 620
rect 21272 536 21324 542
rect 21324 484 21620 490
rect 18524 218 18552 478
rect 18206 190 18552 218
rect 17408 128 17460 134
rect 15906 66 16344 82
rect 17010 76 17408 82
rect 17010 70 17460 76
rect 15906 60 16356 66
rect 15906 54 16304 60
rect 15906 -960 16018 54
rect 16304 2 16356 8
rect 17010 54 17448 70
rect 17010 -960 17122 54
rect 18206 -960 18318 190
rect 18984 66 19320 82
rect 18972 60 19320 66
rect 19024 54 19320 60
rect 18972 2 19024 8
rect 19402 -960 19514 480
rect 20076 128 20128 134
rect 20128 76 20424 82
rect 20076 70 20424 76
rect 20088 54 20424 70
rect 20598 -960 20710 480
rect 21272 478 21620 484
rect 21836 480 21864 598
rect 22020 542 22048 598
rect 22376 604 22724 610
rect 22428 598 22724 604
rect 23020 604 23072 610
rect 22376 546 22428 552
rect 23492 598 23828 614
rect 24872 610 25024 626
rect 28816 672 28868 678
rect 26514 640 26570 649
rect 25832 620 26128 626
rect 25780 614 26128 620
rect 24860 604 25024 610
rect 23020 546 23072 552
rect 24228 564 24440 592
rect 22008 536 22060 542
rect 21284 462 21620 478
rect 21794 -960 21906 480
rect 22008 478 22060 484
rect 23032 480 23060 546
rect 24228 480 24256 564
rect 24412 490 24440 564
rect 24912 598 25024 604
rect 25320 604 25372 610
rect 24860 546 24912 552
rect 25792 598 26128 614
rect 28722 640 28778 649
rect 28092 610 28428 626
rect 28080 604 28428 610
rect 26514 575 26570 584
rect 25320 546 25372 552
rect 22990 -960 23102 480
rect 24186 -960 24298 480
rect 24412 474 24900 490
rect 25332 480 25360 546
rect 26528 480 26556 575
rect 27724 564 27936 592
rect 24412 468 24912 474
rect 24412 462 24860 468
rect 24860 410 24912 416
rect 25290 -960 25402 480
rect 26486 -960 26598 480
rect 26896 474 27232 490
rect 27724 480 27752 564
rect 27908 513 27936 564
rect 28132 598 28428 604
rect 31668 672 31720 678
rect 30286 640 30342 649
rect 28868 620 28948 626
rect 28816 614 28948 620
rect 28828 598 28948 614
rect 29196 610 29532 626
rect 28722 575 28724 584
rect 28080 546 28132 552
rect 28776 575 28778 584
rect 28724 546 28776 552
rect 27894 504 27950 513
rect 26884 468 27232 474
rect 26936 462 27232 468
rect 26884 410 26936 416
rect 27682 -960 27794 480
rect 28920 480 28948 598
rect 29184 604 29532 610
rect 29236 598 29532 604
rect 30104 604 30156 610
rect 29184 546 29236 552
rect 31298 640 31354 649
rect 30342 598 30636 626
rect 30286 575 30342 584
rect 34796 672 34848 678
rect 33598 640 33654 649
rect 31720 620 31832 626
rect 31668 614 31832 620
rect 31680 598 31832 614
rect 32232 598 32444 626
rect 32600 610 32936 626
rect 31298 575 31354 584
rect 30104 546 30156 552
rect 30116 480 30144 546
rect 31312 480 31340 575
rect 27894 439 27950 448
rect 28878 -960 28990 480
rect 30074 -960 30186 480
rect 31270 -960 31382 480
rect 32232 377 32260 598
rect 32416 480 32444 598
rect 32588 604 32936 610
rect 32640 598 32936 604
rect 37280 672 37332 678
rect 34796 614 34848 620
rect 35990 640 36046 649
rect 33598 575 33654 584
rect 32588 546 32640 552
rect 33612 480 33640 575
rect 33874 504 33930 513
rect 32218 368 32274 377
rect 32218 303 32274 312
rect 32374 -960 32486 480
rect 33570 -960 33682 480
rect 33930 462 34132 490
rect 34808 480 34836 614
rect 38384 672 38436 678
rect 37332 620 37536 626
rect 37280 614 37536 620
rect 40684 672 40736 678
rect 38384 614 38436 620
rect 38474 640 38530 649
rect 35990 575 36046 584
rect 37188 604 37240 610
rect 36004 480 36032 575
rect 37292 598 37536 614
rect 37188 546 37240 552
rect 36174 504 36230 513
rect 33874 439 33930 448
rect 34766 -960 34878 480
rect 34978 368 35034 377
rect 35034 326 35236 354
rect 34978 303 35034 312
rect 35962 -960 36074 480
rect 36230 462 36340 490
rect 37200 480 37228 546
rect 38396 480 38424 614
rect 38530 598 38640 626
rect 42800 672 42852 678
rect 40684 614 40736 620
rect 39580 604 39632 610
rect 38474 575 38530 584
rect 39580 546 39632 552
rect 39592 480 39620 546
rect 40696 480 40724 614
rect 40788 610 40940 626
rect 46664 672 46716 678
rect 42852 620 43148 626
rect 42800 614 43148 620
rect 40776 604 40940 610
rect 40828 598 40940 604
rect 41880 604 41932 610
rect 40776 546 40828 552
rect 42812 598 43148 614
rect 44008 610 44344 626
rect 43996 604 44344 610
rect 41880 546 41932 552
rect 44048 598 44344 604
rect 45112 598 45448 626
rect 46664 614 46716 620
rect 48504 672 48556 678
rect 48964 672 49016 678
rect 48556 620 48852 626
rect 48504 614 48852 620
rect 50804 672 50856 678
rect 48964 614 49016 620
rect 43996 546 44048 552
rect 41892 480 41920 546
rect 36174 439 36230 448
rect 37158 -960 37270 480
rect 38354 -960 38466 480
rect 39550 -960 39662 480
rect 39856 400 39908 406
rect 39744 348 39856 354
rect 39744 342 39908 348
rect 39744 326 39896 342
rect 40654 -960 40766 480
rect 41850 -960 41962 480
rect 42044 474 42196 490
rect 42044 468 42208 474
rect 42044 462 42156 468
rect 42156 410 42208 416
rect 42892 400 42944 406
rect 43046 354 43158 480
rect 42944 348 43158 354
rect 42892 342 43158 348
rect 42904 326 43158 342
rect 43046 -960 43158 326
rect 44242 82 44354 480
rect 45112 406 45140 598
rect 46676 480 46704 614
rect 47860 604 47912 610
rect 48516 598 48852 614
rect 47860 546 47912 552
rect 47872 480 47900 546
rect 48976 480 49004 614
rect 49620 610 49956 626
rect 63224 672 63276 678
rect 52550 640 52606 649
rect 50856 620 51152 626
rect 50804 614 51152 620
rect 49608 604 49956 610
rect 49660 598 49956 604
rect 50160 604 50212 610
rect 49608 546 49660 552
rect 50816 598 51152 614
rect 51356 604 51408 610
rect 50160 546 50212 552
rect 54206 640 54262 649
rect 53024 610 53360 626
rect 52550 575 52606 584
rect 53012 604 53360 610
rect 51356 546 51408 552
rect 50172 480 50200 546
rect 51368 480 51396 546
rect 51908 536 51960 542
rect 51960 484 52256 490
rect 45100 400 45152 406
rect 45100 342 45152 348
rect 44100 66 44354 82
rect 44088 60 44354 66
rect 44140 54 44354 60
rect 44088 2 44140 8
rect 44242 -960 44354 54
rect 45438 82 45550 480
rect 45744 128 45796 134
rect 45438 76 45744 82
rect 45438 70 45796 76
rect 45438 54 45784 70
rect 46216 66 46552 82
rect 46204 60 46552 66
rect 45438 -960 45550 54
rect 46256 54 46552 60
rect 46204 2 46256 8
rect 46634 -960 46746 480
rect 47400 128 47452 134
rect 47452 76 47748 82
rect 47400 70 47748 76
rect 47412 54 47748 70
rect 47830 -960 47942 480
rect 48934 -960 49046 480
rect 50130 -960 50242 480
rect 51326 -960 51438 480
rect 51908 478 52256 484
rect 52564 480 52592 575
rect 53064 598 53360 604
rect 53576 598 53788 626
rect 53012 546 53064 552
rect 53576 513 53604 598
rect 53562 504 53618 513
rect 51920 462 52256 478
rect 52522 -960 52634 480
rect 53760 480 53788 598
rect 56046 640 56102 649
rect 54262 598 54556 626
rect 54944 604 54996 610
rect 54206 575 54262 584
rect 57610 640 57666 649
rect 56428 610 56764 626
rect 56046 575 56102 584
rect 56416 604 56764 610
rect 54944 546 54996 552
rect 54956 480 54984 546
rect 55310 504 55366 513
rect 53562 439 53618 448
rect 53718 -960 53830 480
rect 54914 -960 55026 480
rect 55366 462 55660 490
rect 56060 480 56088 575
rect 56468 598 56764 604
rect 56416 546 56468 552
rect 57256 564 57468 592
rect 58438 640 58494 649
rect 57666 598 57960 626
rect 57610 575 57666 584
rect 59818 640 59874 649
rect 58438 575 58494 584
rect 57256 480 57284 564
rect 57440 513 57468 564
rect 57426 504 57482 513
rect 55310 439 55366 448
rect 56018 -960 56130 480
rect 57214 -960 57326 480
rect 58452 480 58480 575
rect 59464 564 59676 592
rect 60830 640 60886 649
rect 59874 598 60168 626
rect 59818 575 59874 584
rect 62118 640 62174 649
rect 60830 575 60886 584
rect 62028 604 62080 610
rect 59464 513 59492 564
rect 58806 504 58862 513
rect 57426 439 57482 448
rect 58410 -960 58522 480
rect 59450 504 59506 513
rect 58862 462 59064 490
rect 58806 439 58862 448
rect 59648 480 59676 564
rect 60844 480 60872 575
rect 62174 598 62468 626
rect 64328 672 64380 678
rect 63224 614 63276 620
rect 62118 575 62174 584
rect 62028 546 62080 552
rect 61106 504 61162 513
rect 59450 439 59506 448
rect 59606 -960 59718 480
rect 60802 -960 60914 480
rect 61162 462 61364 490
rect 62040 480 62068 546
rect 63236 480 63264 614
rect 63328 610 63664 626
rect 65616 672 65668 678
rect 64328 614 64380 620
rect 63316 604 63664 610
rect 63368 598 63664 604
rect 63316 546 63368 552
rect 64340 480 64368 614
rect 64432 610 64768 626
rect 66720 672 66772 678
rect 65668 620 65872 626
rect 65616 614 65872 620
rect 68008 672 68060 678
rect 66720 614 66772 620
rect 64420 604 64768 610
rect 64472 598 64768 604
rect 65524 604 65576 610
rect 64420 546 64472 552
rect 65628 598 65872 614
rect 65524 546 65576 552
rect 65536 480 65564 546
rect 66732 480 66760 614
rect 66824 610 67068 626
rect 66812 604 67068 610
rect 66864 598 67068 604
rect 67744 598 67956 626
rect 69112 672 69164 678
rect 68060 620 68172 626
rect 68008 614 68172 620
rect 70584 672 70636 678
rect 69112 614 69164 620
rect 70472 620 70584 626
rect 133236 672 133288 678
rect 70472 614 70636 620
rect 68020 598 68172 614
rect 66812 546 66864 552
rect 67744 542 67772 598
rect 67732 536 67784 542
rect 61106 439 61162 448
rect 61998 -960 62110 480
rect 63194 -960 63306 480
rect 64298 -960 64410 480
rect 65494 -960 65606 480
rect 66690 -960 66802 480
rect 67732 478 67784 484
rect 67928 480 67956 598
rect 69124 480 69152 614
rect 70308 604 70360 610
rect 70472 598 70624 614
rect 71240 610 71576 626
rect 71228 604 71576 610
rect 70308 546 70360 552
rect 71280 598 71576 604
rect 72344 598 72680 626
rect 73540 598 73876 626
rect 74644 598 74980 626
rect 76944 610 77280 626
rect 78048 610 78384 626
rect 79152 610 79488 626
rect 80348 610 80684 626
rect 81452 610 81788 626
rect 82740 610 82892 626
rect 76196 604 76248 610
rect 71228 546 71280 552
rect 69388 536 69440 542
rect 69276 484 69388 490
rect 67886 -960 67998 480
rect 69082 -960 69194 480
rect 69276 478 69440 484
rect 70320 480 70348 546
rect 69276 462 69428 478
rect 70278 -960 70390 480
rect 71320 400 71372 406
rect 71474 354 71586 480
rect 72344 406 72372 598
rect 71372 348 71586 354
rect 71320 342 71586 348
rect 72332 400 72384 406
rect 72332 342 72384 348
rect 72424 400 72476 406
rect 72578 354 72690 480
rect 73540 406 73568 598
rect 72476 348 72690 354
rect 72424 342 72690 348
rect 73528 400 73580 406
rect 73528 342 73580 348
rect 73620 400 73672 406
rect 73774 354 73886 480
rect 74644 406 74672 598
rect 76196 546 76248 552
rect 76932 604 77280 610
rect 76984 598 77280 604
rect 77392 604 77444 610
rect 76932 546 76984 552
rect 77392 546 77444 552
rect 78036 604 78384 610
rect 78088 598 78384 604
rect 78588 604 78640 610
rect 78036 546 78088 552
rect 78588 546 78640 552
rect 79140 604 79488 610
rect 79192 598 79488 604
rect 79692 604 79744 610
rect 79140 546 79192 552
rect 79692 546 79744 552
rect 80336 604 80684 610
rect 80388 598 80684 604
rect 80888 604 80940 610
rect 80336 546 80388 552
rect 80888 546 80940 552
rect 81440 604 81788 610
rect 81492 598 81788 604
rect 82084 604 82136 610
rect 81440 546 81492 552
rect 82084 546 82136 552
rect 82728 604 82892 610
rect 82780 598 82892 604
rect 83292 598 83504 626
rect 82728 546 82780 552
rect 76208 480 76236 546
rect 77404 480 77432 546
rect 78600 480 78628 546
rect 79704 480 79732 546
rect 80900 480 80928 546
rect 82096 480 82124 546
rect 83292 480 83320 598
rect 83476 490 83504 598
rect 84488 598 85192 626
rect 85684 598 85896 626
rect 73672 348 73886 354
rect 73620 342 73886 348
rect 74632 400 74684 406
rect 74632 342 74684 348
rect 71332 326 71586 342
rect 72436 326 72690 342
rect 73632 326 73886 342
rect 71474 -960 71586 326
rect 72578 -960 72690 326
rect 73774 -960 73886 326
rect 74970 82 75082 480
rect 74970 54 76084 82
rect 74970 -960 75082 54
rect 76166 -960 76278 480
rect 77362 -960 77474 480
rect 78558 -960 78670 480
rect 79662 -960 79774 480
rect 80858 -960 80970 480
rect 82054 -960 82166 480
rect 83250 -960 83362 480
rect 83476 462 84088 490
rect 84488 480 84516 598
rect 85684 480 85712 598
rect 85868 490 85896 598
rect 86880 598 87492 626
rect 87984 598 88596 626
rect 89180 598 89392 626
rect 84446 -960 84558 480
rect 85642 -960 85754 480
rect 85868 462 86296 490
rect 86880 480 86908 598
rect 87984 480 88012 598
rect 89180 480 89208 598
rect 89364 490 89392 598
rect 90376 598 90896 626
rect 91572 598 92000 626
rect 92768 598 93196 626
rect 93964 598 94300 626
rect 95160 598 95404 626
rect 96264 598 96600 626
rect 97460 598 97704 626
rect 98656 598 98808 626
rect 99852 598 100004 626
rect 105616 598 105768 626
rect 106812 598 106964 626
rect 107916 598 108160 626
rect 109020 598 109356 626
rect 110216 598 110552 626
rect 111320 598 111656 626
rect 112424 598 112852 626
rect 113620 598 114048 626
rect 114724 598 115244 626
rect 115828 598 116440 626
rect 86838 -960 86950 480
rect 87942 -960 88054 480
rect 89138 -960 89250 480
rect 89364 462 89792 490
rect 90376 480 90404 598
rect 91572 480 91600 598
rect 92768 480 92796 598
rect 93964 480 93992 598
rect 95160 480 95188 598
rect 96264 480 96292 598
rect 97460 480 97488 598
rect 98656 480 98684 598
rect 99852 480 99880 598
rect 105740 480 105768 598
rect 106936 480 106964 598
rect 108132 480 108160 598
rect 109328 480 109356 598
rect 110524 480 110552 598
rect 111628 480 111656 598
rect 112824 480 112852 598
rect 114020 480 114048 598
rect 115216 480 115244 598
rect 116412 480 116440 598
rect 117424 598 117636 626
rect 118128 598 118832 626
rect 119324 598 119936 626
rect 117424 490 117452 598
rect 90334 -960 90446 480
rect 91530 -960 91642 480
rect 92726 -960 92838 480
rect 93922 -960 94034 480
rect 95118 -960 95230 480
rect 96222 -960 96334 480
rect 97418 -960 97530 480
rect 98614 -960 98726 480
rect 99810 -960 99922 480
rect 101006 -960 101118 480
rect 102202 -960 102314 480
rect 103306 -960 103418 480
rect 104502 -960 104614 480
rect 105698 -960 105810 480
rect 106894 -960 107006 480
rect 108090 -960 108202 480
rect 109286 -960 109398 480
rect 110482 -960 110594 480
rect 111586 -960 111698 480
rect 112782 -960 112894 480
rect 113978 -960 114090 480
rect 115174 -960 115286 480
rect 116370 -960 116482 480
rect 117024 462 117452 490
rect 117608 480 117636 598
rect 118804 480 118832 598
rect 119908 480 119936 598
rect 120920 598 121132 626
rect 121532 610 121868 626
rect 121532 604 121880 610
rect 121532 598 121828 604
rect 120920 490 120948 598
rect 117566 -960 117678 480
rect 118762 -960 118874 480
rect 119866 -960 119978 480
rect 120428 462 120948 490
rect 121104 480 121132 598
rect 121828 546 121880 552
rect 122288 604 122340 610
rect 122288 546 122340 552
rect 123312 598 123524 626
rect 123832 610 124168 626
rect 124936 610 125272 626
rect 126132 610 126468 626
rect 127236 610 127572 626
rect 128340 610 128676 626
rect 123832 604 124180 610
rect 123832 598 124128 604
rect 122300 480 122328 546
rect 123312 490 123340 598
rect 121062 -960 121174 480
rect 122258 -960 122370 480
rect 122728 462 123340 490
rect 123496 480 123524 598
rect 124128 546 124180 552
rect 124680 604 124732 610
rect 124936 604 125284 610
rect 124936 598 125232 604
rect 124680 546 124732 552
rect 125232 546 125284 552
rect 125876 604 125928 610
rect 126132 604 126480 610
rect 126132 598 126428 604
rect 125876 546 125928 552
rect 126428 546 126480 552
rect 126980 604 127032 610
rect 127236 604 127584 610
rect 127236 598 127532 604
rect 126980 546 127032 552
rect 127532 546 127584 552
rect 128176 604 128228 610
rect 128340 604 128688 610
rect 128340 598 128636 604
rect 128176 546 128228 552
rect 128636 546 128688 552
rect 129372 604 129424 610
rect 130640 598 130976 626
rect 131744 598 132080 626
rect 132940 620 133236 626
rect 134156 672 134208 678
rect 132940 614 133288 620
rect 132940 598 133276 614
rect 133892 610 134044 626
rect 134156 614 134208 620
rect 136180 672 136232 678
rect 137652 672 137704 678
rect 136232 620 136344 626
rect 136180 614 136344 620
rect 133880 604 134044 610
rect 129372 546 129424 552
rect 124692 480 124720 546
rect 125888 480 125916 546
rect 126992 480 127020 546
rect 128188 480 128216 546
rect 129384 480 129412 546
rect 123454 -960 123566 480
rect 124650 -960 124762 480
rect 125846 -960 125958 480
rect 126950 -960 127062 480
rect 128146 -960 128258 480
rect 129342 -960 129454 480
rect 129832 128 129884 134
rect 129536 76 129832 82
rect 129536 70 129884 76
rect 130292 128 130344 134
rect 130538 82 130650 480
rect 130948 406 130976 598
rect 130936 400 130988 406
rect 130936 342 130988 348
rect 131734 354 131846 480
rect 132052 406 132080 598
rect 133932 598 134044 604
rect 133880 546 133932 552
rect 134168 480 134196 614
rect 135260 604 135312 610
rect 136192 598 136344 614
rect 137448 610 137600 626
rect 138756 672 138808 678
rect 137652 614 137704 620
rect 138552 620 138756 626
rect 140044 672 140096 678
rect 138552 614 138808 620
rect 136456 604 136508 610
rect 135260 546 135312 552
rect 137448 604 137612 610
rect 137448 598 137560 604
rect 136456 546 136508 552
rect 137560 546 137612 552
rect 134984 536 135036 542
rect 135036 484 135148 490
rect 131948 400 132000 406
rect 131734 348 131948 354
rect 131734 342 132000 348
rect 132040 400 132092 406
rect 132040 342 132092 348
rect 132930 354 133042 480
rect 133144 400 133196 406
rect 132930 348 133144 354
rect 132930 342 133196 348
rect 130344 76 130650 82
rect 130292 70 130650 76
rect 129536 54 129872 70
rect 130304 54 130650 70
rect 130538 -960 130650 54
rect 131734 326 131988 342
rect 132930 326 133184 342
rect 131734 -960 131846 326
rect 132930 -960 133042 326
rect 134126 -960 134238 480
rect 134984 478 135148 484
rect 135272 480 135300 546
rect 136468 480 136496 546
rect 137664 480 137692 614
rect 138552 598 138796 614
rect 139748 610 139992 626
rect 151360 672 151412 678
rect 142066 640 142122 649
rect 140044 614 140096 620
rect 138848 604 138900 610
rect 139748 604 140004 610
rect 139748 598 139952 604
rect 138848 546 138900 552
rect 139952 546 140004 552
rect 138860 480 138888 546
rect 140056 480 140084 614
rect 141240 604 141292 610
rect 141956 598 142066 626
rect 143446 640 143502 649
rect 142066 575 142122 584
rect 142264 598 142476 626
rect 143152 598 143446 626
rect 141240 546 141292 552
rect 141056 536 141108 542
rect 140852 484 141056 490
rect 134996 462 135148 478
rect 135230 -960 135342 480
rect 136426 -960 136538 480
rect 137622 -960 137734 480
rect 138818 -960 138930 480
rect 140014 -960 140126 480
rect 140852 478 141108 484
rect 141252 480 141280 546
rect 142068 536 142120 542
rect 142264 490 142292 598
rect 142120 484 142292 490
rect 140852 462 141096 478
rect 141210 -960 141322 480
rect 142068 478 142292 484
rect 142448 480 142476 598
rect 144734 640 144790 649
rect 143446 575 143502 584
rect 143552 598 143764 626
rect 144256 610 144592 626
rect 144256 604 144604 610
rect 144256 598 144552 604
rect 143552 480 143580 598
rect 143736 513 143764 598
rect 145746 640 145802 649
rect 145452 598 145746 626
rect 144734 575 144790 584
rect 147126 640 147182 649
rect 146556 610 146892 626
rect 145746 575 145802 584
rect 145932 604 145984 610
rect 144552 546 144604 552
rect 143722 504 143778 513
rect 142080 462 142292 478
rect 142406 -960 142518 480
rect 143510 -960 143622 480
rect 144748 480 144776 575
rect 146556 604 146904 610
rect 146556 598 146852 604
rect 145932 546 145984 552
rect 148966 640 149022 649
rect 147126 575 147182 584
rect 148324 604 148376 610
rect 146852 546 146904 552
rect 145944 480 145972 546
rect 147140 480 147168 575
rect 148856 598 148966 626
rect 150622 640 150678 649
rect 148966 575 149022 584
rect 149348 598 149560 626
rect 148324 546 148376 552
rect 147770 504 147826 513
rect 143722 439 143778 448
rect 144706 -960 144818 480
rect 145902 -960 146014 480
rect 147098 -960 147210 480
rect 147660 462 147770 490
rect 148336 480 148364 546
rect 149348 513 149376 598
rect 149334 504 149390 513
rect 147770 439 147826 448
rect 148294 -960 148406 480
rect 149532 480 149560 598
rect 151064 620 151360 626
rect 153016 672 153068 678
rect 151064 614 151412 620
rect 151818 640 151874 649
rect 151064 598 151400 614
rect 150622 575 150678 584
rect 152260 610 152596 626
rect 153660 672 153712 678
rect 153016 614 153068 620
rect 153364 620 153660 626
rect 155408 672 155460 678
rect 153364 614 153712 620
rect 152260 604 152608 610
rect 152260 598 152556 604
rect 151818 575 151874 584
rect 150254 504 150310 513
rect 149334 439 149390 448
rect 149490 -960 149602 480
rect 149960 462 150254 490
rect 150636 480 150664 575
rect 151832 480 151860 575
rect 152556 546 152608 552
rect 153028 480 153056 614
rect 153364 598 153700 614
rect 154468 610 154804 626
rect 162768 672 162820 678
rect 155408 614 155460 620
rect 154212 604 154264 610
rect 154468 604 154816 610
rect 154468 598 154764 604
rect 154212 546 154264 552
rect 154764 546 154816 552
rect 154224 480 154252 546
rect 155420 480 155448 614
rect 156768 610 157104 626
rect 156604 604 156656 610
rect 156768 604 157116 610
rect 156768 598 157064 604
rect 156604 546 156656 552
rect 157872 598 158208 626
rect 157064 546 157116 552
rect 156616 480 156644 546
rect 158180 542 158208 598
rect 158904 604 158956 610
rect 160172 598 160508 626
rect 161276 610 161612 626
rect 162472 620 162768 626
rect 164884 672 164936 678
rect 164790 640 164846 649
rect 162472 614 162820 620
rect 161276 604 161624 610
rect 161276 598 161572 604
rect 158904 546 158956 552
rect 158168 536 158220 542
rect 150254 439 150310 448
rect 150594 -960 150706 480
rect 151790 -960 151902 480
rect 152986 -960 153098 480
rect 154182 -960 154294 480
rect 155378 -960 155490 480
rect 155960 128 156012 134
rect 155664 76 155960 82
rect 155664 70 156012 76
rect 155664 54 156000 70
rect 156574 -960 156686 480
rect 157524 128 157576 134
rect 157770 82 157882 480
rect 158168 478 158220 484
rect 158916 480 158944 546
rect 159732 536 159784 542
rect 157576 76 157882 82
rect 157524 70 157882 76
rect 157536 54 157882 70
rect 157770 -960 157882 54
rect 158874 -960 158986 480
rect 159732 478 159784 484
rect 159744 354 159772 478
rect 160070 354 160182 480
rect 160480 406 160508 598
rect 162472 598 162808 614
rect 163688 604 163740 610
rect 161572 546 161624 552
rect 164680 598 164790 626
rect 166080 672 166132 678
rect 164884 614 164936 620
rect 164790 575 164846 584
rect 163688 546 163740 552
rect 159744 326 160182 354
rect 160468 400 160520 406
rect 160468 342 160520 348
rect 159364 128 159416 134
rect 159068 76 159364 82
rect 159068 70 159416 76
rect 159068 54 159404 70
rect 160070 -960 160182 326
rect 161266 82 161378 480
rect 162462 354 162574 480
rect 163424 474 163576 490
rect 163700 480 163728 546
rect 164896 480 164924 614
rect 165876 610 166028 626
rect 167092 672 167144 678
rect 166080 614 166132 620
rect 166980 620 167092 626
rect 169576 672 169628 678
rect 167366 640 167422 649
rect 166980 614 167144 620
rect 165876 604 166040 610
rect 165876 598 165988 604
rect 165988 546 166040 552
rect 166092 480 166120 614
rect 166980 598 167132 614
rect 167196 598 167366 626
rect 167196 480 167224 598
rect 169482 640 169538 649
rect 167366 575 167422 584
rect 168380 604 168432 610
rect 169280 598 169482 626
rect 180892 672 180944 678
rect 171966 640 172022 649
rect 169576 614 169628 620
rect 169482 575 169538 584
rect 168380 546 168432 552
rect 168392 480 168420 546
rect 169588 480 169616 614
rect 170384 610 170720 626
rect 170384 604 170732 610
rect 170384 598 170680 604
rect 170680 546 170732 552
rect 170784 598 170996 626
rect 170784 480 170812 598
rect 163412 468 163576 474
rect 163464 462 163576 468
rect 163412 410 163464 416
rect 162676 400 162728 406
rect 162462 348 162676 354
rect 162462 342 162728 348
rect 162462 326 162716 342
rect 161480 128 161532 134
rect 161266 76 161480 82
rect 161266 70 161532 76
rect 161266 54 161520 70
rect 161266 -960 161378 54
rect 162462 -960 162574 326
rect 163658 -960 163770 480
rect 164854 -960 164966 480
rect 166050 -960 166162 480
rect 167154 -960 167266 480
rect 168194 368 168250 377
rect 168084 326 168194 354
rect 168194 303 168250 312
rect 168350 -960 168462 480
rect 169546 -960 169658 480
rect 170742 -960 170854 480
rect 170968 377 170996 598
rect 172978 640 173034 649
rect 172684 598 172978 626
rect 171966 575 172022 584
rect 175462 640 175518 649
rect 172978 575 173034 584
rect 173164 604 173216 610
rect 171980 480 172008 575
rect 173164 546 173216 552
rect 174096 598 174308 626
rect 173176 480 173204 546
rect 173898 504 173954 513
rect 170954 368 171010 377
rect 171690 368 171746 377
rect 171488 326 171690 354
rect 170954 303 171010 312
rect 171690 303 171746 312
rect 171938 -960 172050 480
rect 173134 -960 173246 480
rect 173788 462 173898 490
rect 174096 490 174124 598
rect 173898 439 173954 448
rect 174004 462 174124 490
rect 174280 480 174308 598
rect 176382 640 176438 649
rect 176088 598 176382 626
rect 175462 575 175518 584
rect 179050 640 179106 649
rect 176382 575 176438 584
rect 176672 598 176884 626
rect 175476 480 175504 575
rect 176672 480 176700 598
rect 176856 513 176884 598
rect 177684 598 177896 626
rect 176842 504 176898 513
rect 174004 377 174032 462
rect 173990 368 174046 377
rect 173990 303 174046 312
rect 174238 -960 174350 480
rect 175186 368 175242 377
rect 174984 326 175186 354
rect 175186 303 175242 312
rect 175434 -960 175546 480
rect 176630 -960 176742 480
rect 177486 504 177542 513
rect 177192 462 177486 490
rect 176842 439 176898 448
rect 177486 439 177542 448
rect 177684 377 177712 598
rect 177868 480 177896 598
rect 180246 640 180302 649
rect 179492 610 179828 626
rect 179492 604 179840 610
rect 179492 598 179788 604
rect 179050 575 179106 584
rect 179064 480 179092 575
rect 180596 620 180892 626
rect 183744 672 183796 678
rect 182086 640 182142 649
rect 180596 614 180944 620
rect 180596 598 180932 614
rect 181272 598 181484 626
rect 181792 598 182086 626
rect 180246 575 180302 584
rect 179788 546 179840 552
rect 180260 480 180288 575
rect 177670 368 177726 377
rect 177670 303 177726 312
rect 177826 -960 177938 480
rect 178682 368 178738 377
rect 178388 326 178682 354
rect 178682 303 178738 312
rect 179022 -960 179134 480
rect 180218 -960 180330 480
rect 181272 377 181300 598
rect 181456 480 181484 598
rect 182896 610 183232 626
rect 186136 672 186188 678
rect 183744 614 183796 620
rect 184938 640 184994 649
rect 182086 575 182142 584
rect 182548 604 182600 610
rect 182896 604 183244 610
rect 182896 598 183192 604
rect 182548 546 182600 552
rect 183192 546 183244 552
rect 182560 480 182588 546
rect 183756 480 183784 614
rect 191104 672 191156 678
rect 186136 614 186188 620
rect 184938 575 184994 584
rect 184952 480 184980 575
rect 186148 480 186176 614
rect 187404 598 187740 626
rect 188600 598 188844 626
rect 189704 610 190040 626
rect 190808 620 191104 626
rect 194416 672 194468 678
rect 192298 640 192354 649
rect 190808 614 191156 620
rect 189704 604 190052 610
rect 189704 598 190000 604
rect 187712 542 187740 598
rect 187700 536 187752 542
rect 186594 504 186650 513
rect 181258 368 181314 377
rect 181258 303 181314 312
rect 181414 -960 181526 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184296 128 184348 134
rect 184000 76 184296 82
rect 184000 70 184348 76
rect 184000 54 184336 70
rect 184910 -960 185022 480
rect 185492 128 185544 134
rect 185196 76 185492 82
rect 185196 70 185544 76
rect 185196 54 185532 70
rect 186106 -960 186218 480
rect 186300 462 186594 490
rect 186594 439 186650 448
rect 187302 218 187414 480
rect 187700 478 187752 484
rect 186976 202 187414 218
rect 186964 196 187414 202
rect 187016 190 187414 196
rect 186964 138 187016 144
rect 187302 -960 187414 190
rect 188252 128 188304 134
rect 188498 82 188610 480
rect 188816 377 188844 598
rect 190808 598 191144 614
rect 192004 598 192298 626
rect 211620 672 211672 678
rect 194416 614 194468 620
rect 195610 640 195666 649
rect 192298 575 192354 584
rect 193220 604 193272 610
rect 190000 546 190052 552
rect 193220 546 193272 552
rect 191012 536 191064 542
rect 189906 504 189962 513
rect 188802 368 188858 377
rect 188802 303 188858 312
rect 188304 76 188610 82
rect 188252 70 188610 76
rect 188264 54 188610 70
rect 188498 -960 188610 54
rect 189694 218 189806 480
rect 189906 439 189962 448
rect 189920 218 189948 439
rect 189694 190 189948 218
rect 190798 354 190910 480
rect 191012 478 191064 484
rect 192944 536 192996 542
rect 192996 484 193108 490
rect 191024 354 191052 478
rect 190798 326 191052 354
rect 191994 354 192106 480
rect 192944 478 193108 484
rect 193232 480 193260 546
rect 194046 504 194102 513
rect 192956 462 193108 478
rect 192206 368 192262 377
rect 191994 326 192206 354
rect 189694 -960 189806 190
rect 190798 -960 190910 326
rect 191994 -960 192106 326
rect 192206 303 192262 312
rect 193190 -960 193302 480
rect 194102 462 194212 490
rect 194428 480 194456 614
rect 197910 640 197966 649
rect 195610 575 195666 584
rect 196808 604 196860 610
rect 195624 480 195652 575
rect 200026 640 200082 649
rect 197910 575 197966 584
rect 199108 604 199160 610
rect 196808 546 196860 552
rect 196820 480 196848 546
rect 197924 480 197952 575
rect 199916 598 200026 626
rect 203890 640 203946 649
rect 203320 610 203656 626
rect 203320 604 203668 610
rect 203320 598 203616 604
rect 200026 575 200082 584
rect 199108 546 199160 552
rect 200132 564 200344 592
rect 198922 504 198978 513
rect 194046 439 194102 448
rect 194386 -960 194498 480
rect 195244 400 195296 406
rect 195296 348 195408 354
rect 195244 342 195408 348
rect 195256 326 195408 342
rect 195582 -960 195694 480
rect 196622 368 196678 377
rect 196512 326 196622 354
rect 196622 303 196678 312
rect 196778 -960 196890 480
rect 197726 96 197782 105
rect 197616 54 197726 82
rect 197726 31 197782 40
rect 197882 -960 197994 480
rect 198812 462 198922 490
rect 199120 480 199148 546
rect 198922 439 198978 448
rect 199078 -960 199190 480
rect 200132 377 200160 564
rect 200316 480 200344 564
rect 201512 564 201724 592
rect 201314 504 201370 513
rect 200118 368 200174 377
rect 200118 303 200174 312
rect 200274 -960 200386 480
rect 201112 462 201314 490
rect 201512 480 201540 564
rect 201314 439 201370 448
rect 201470 -960 201582 480
rect 201696 105 201724 564
rect 202524 564 202736 592
rect 202524 377 202552 564
rect 202708 480 202736 564
rect 203890 575 203946 584
rect 204166 640 204222 649
rect 207386 640 207442 649
rect 205620 610 205772 626
rect 205620 604 205784 610
rect 205620 598 205732 604
rect 204166 575 204168 584
rect 203616 546 203668 552
rect 203904 480 203932 575
rect 204220 575 204222 584
rect 204168 546 204220 552
rect 204916 564 205128 592
rect 204916 513 204944 564
rect 204902 504 204958 513
rect 202510 368 202566 377
rect 202510 303 202566 312
rect 202418 232 202474 241
rect 202216 190 202418 218
rect 202418 167 202474 176
rect 201682 96 201738 105
rect 201682 31 201738 40
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205100 480 205128 564
rect 205732 546 205784 552
rect 206020 564 206232 592
rect 208214 640 208270 649
rect 207920 598 208214 626
rect 207386 575 207442 584
rect 208214 575 208270 584
rect 208398 640 208454 649
rect 209318 640 209374 649
rect 208398 575 208454 584
rect 208596 598 208808 626
rect 209024 598 209318 626
rect 206020 513 206048 564
rect 206006 504 206062 513
rect 204902 439 204958 448
rect 204810 368 204866 377
rect 204516 326 204810 354
rect 204810 303 204866 312
rect 205058 -960 205170 480
rect 206204 480 206232 564
rect 206926 504 206982 513
rect 206006 439 206062 448
rect 206162 -960 206274 480
rect 206724 462 206926 490
rect 207400 480 207428 575
rect 208412 542 208440 575
rect 208400 536 208452 542
rect 206926 439 206982 448
rect 207358 -960 207470 480
rect 208400 478 208452 484
rect 208596 480 208624 598
rect 208554 -960 208666 480
rect 208780 377 208808 598
rect 210128 610 210464 626
rect 209318 575 209374 584
rect 209780 604 209832 610
rect 210128 604 210476 610
rect 210128 598 210424 604
rect 209780 546 209832 552
rect 210424 546 210476 552
rect 210804 598 211016 626
rect 211324 620 211620 626
rect 215668 672 215720 678
rect 211324 614 211672 620
rect 213366 640 213422 649
rect 211324 598 211660 614
rect 212172 604 212224 610
rect 209792 480 209820 546
rect 210804 513 210832 598
rect 210790 504 210846 513
rect 208766 368 208822 377
rect 208766 303 208822 312
rect 209750 -960 209862 480
rect 210988 480 211016 598
rect 219532 672 219584 678
rect 216126 640 216182 649
rect 215668 614 215720 620
rect 213366 575 213422 584
rect 214472 604 214524 610
rect 212172 546 212224 552
rect 212184 480 212212 546
rect 210790 439 210846 448
rect 210946 -960 211058 480
rect 212142 -960 212254 480
rect 212428 474 212580 490
rect 213380 480 213408 575
rect 214472 546 214524 552
rect 214484 480 214512 546
rect 215680 480 215708 614
rect 215832 598 216126 626
rect 216936 598 217272 626
rect 218132 610 218468 626
rect 219236 620 219532 626
rect 226156 672 226208 678
rect 219236 614 219584 620
rect 220450 640 220506 649
rect 218132 604 218480 610
rect 218132 598 218428 604
rect 216126 575 216182 584
rect 212428 468 212592 474
rect 212428 462 212540 468
rect 212540 410 212592 416
rect 213338 -960 213450 480
rect 213532 66 213868 82
rect 213532 60 213880 66
rect 213532 54 213828 60
rect 213828 2 213880 8
rect 214442 -960 214554 480
rect 215024 128 215076 134
rect 214728 76 215024 82
rect 214728 70 215076 76
rect 214728 54 215064 70
rect 215638 -960 215750 480
rect 216588 468 216640 474
rect 216588 410 216640 416
rect 216600 354 216628 410
rect 216834 354 216946 480
rect 217244 406 217272 598
rect 219236 598 219572 614
rect 223854 640 223910 649
rect 221536 598 221872 626
rect 220450 575 220506 584
rect 218428 546 218480 552
rect 220464 480 220492 575
rect 216600 326 216946 354
rect 217232 400 217284 406
rect 217232 342 217284 348
rect 216834 -960 216946 326
rect 218030 82 218142 480
rect 217796 66 218142 82
rect 217784 60 218142 66
rect 217836 54 218142 60
rect 217784 2 217836 8
rect 218030 -960 218142 54
rect 219226 82 219338 480
rect 220188 338 220340 354
rect 220176 332 220340 338
rect 220228 326 220340 332
rect 220176 274 220228 280
rect 219440 128 219492 134
rect 219226 76 219440 82
rect 219226 70 219492 76
rect 219226 54 219480 70
rect 219226 -960 219338 54
rect 220422 -960 220534 480
rect 221526 354 221638 480
rect 221844 474 221872 598
rect 222752 604 222804 610
rect 223744 598 223854 626
rect 224940 610 225092 626
rect 223854 575 223910 584
rect 223948 604 224000 610
rect 222752 546 222804 552
rect 224940 604 225104 610
rect 224940 598 225052 604
rect 223948 546 224000 552
rect 225052 546 225104 552
rect 225156 598 225368 626
rect 226044 620 226156 626
rect 231032 672 231084 678
rect 228730 640 228786 649
rect 226044 614 226208 620
rect 226044 598 226196 614
rect 226352 598 226564 626
rect 222764 480 222792 546
rect 223960 480 223988 546
rect 225156 480 225184 598
rect 225340 542 225368 598
rect 225328 536 225380 542
rect 221832 468 221884 474
rect 221832 410 221884 416
rect 221740 400 221792 406
rect 221526 348 221740 354
rect 221526 342 221792 348
rect 222476 400 222528 406
rect 222528 348 222640 354
rect 222476 342 222640 348
rect 221526 326 221780 342
rect 222488 326 222640 342
rect 221526 -960 221638 326
rect 222722 -960 222834 480
rect 223918 -960 224030 480
rect 225114 -960 225226 480
rect 225328 478 225380 484
rect 226352 480 226380 598
rect 226536 542 226564 598
rect 227272 598 227576 626
rect 226524 536 226576 542
rect 226310 -960 226422 480
rect 226524 478 226576 484
rect 227272 406 227300 598
rect 227548 480 227576 598
rect 230938 640 230994 649
rect 228730 575 228786 584
rect 229836 604 229888 610
rect 228744 480 228772 575
rect 230644 598 230938 626
rect 234620 672 234672 678
rect 231032 614 231084 620
rect 230938 575 230994 584
rect 229836 546 229888 552
rect 229652 536 229704 542
rect 229448 484 229652 490
rect 227260 400 227312 406
rect 227260 342 227312 348
rect 227148 202 227392 218
rect 227148 196 227404 202
rect 227148 190 227352 196
rect 227352 138 227404 144
rect 227506 -960 227618 480
rect 228548 128 228600 134
rect 228344 76 228548 82
rect 228344 70 228600 76
rect 228344 54 228588 70
rect 228702 -960 228814 480
rect 229448 478 229704 484
rect 229848 480 229876 546
rect 231044 480 231072 614
rect 231748 610 231900 626
rect 231748 604 231912 610
rect 231748 598 231860 604
rect 231860 546 231912 552
rect 232056 598 232268 626
rect 229448 462 229692 478
rect 229806 -960 229918 480
rect 231002 -960 231114 480
rect 232056 202 232084 598
rect 232240 480 232268 598
rect 233252 598 233464 626
rect 235448 672 235500 678
rect 234620 614 234672 620
rect 235152 620 235448 626
rect 237748 672 237800 678
rect 235152 614 235500 620
rect 235814 640 235870 649
rect 233148 536 233200 542
rect 232852 484 233148 490
rect 232044 196 232096 202
rect 232044 138 232096 144
rect 232198 -960 232310 480
rect 232852 478 233200 484
rect 232852 462 233188 478
rect 233252 134 233280 598
rect 233436 480 233464 598
rect 233240 128 233292 134
rect 233240 70 233292 76
rect 233394 -960 233506 480
rect 234048 474 234384 490
rect 234632 480 234660 614
rect 235152 598 235488 614
rect 237452 620 237748 626
rect 242900 672 242952 678
rect 238850 640 238906 649
rect 237452 614 237800 620
rect 235814 575 235870 584
rect 237012 604 237064 610
rect 235828 480 235856 575
rect 237452 598 237788 614
rect 238116 604 238168 610
rect 237012 546 237064 552
rect 238556 598 238850 626
rect 247960 672 248012 678
rect 242900 614 242952 620
rect 244094 640 244150 649
rect 238850 575 238906 584
rect 239312 604 239364 610
rect 238116 546 238168 552
rect 239312 546 239364 552
rect 240508 604 240560 610
rect 240508 546 240560 552
rect 241532 564 241744 592
rect 237024 480 237052 546
rect 238128 480 238156 546
rect 239324 480 239352 546
rect 234048 468 234396 474
rect 234048 462 234344 468
rect 234344 410 234396 416
rect 234590 -960 234702 480
rect 235786 -960 235898 480
rect 236552 128 236604 134
rect 236256 76 236552 82
rect 236256 70 236604 76
rect 236256 54 236592 70
rect 236982 -960 237094 480
rect 238086 -960 238198 480
rect 239282 -960 239394 480
rect 239660 474 239996 490
rect 240520 480 240548 546
rect 239660 468 240008 474
rect 239660 462 239956 468
rect 239956 410 240008 416
rect 240478 -960 240590 480
rect 241532 354 241560 564
rect 241716 480 241744 564
rect 242254 504 242310 513
rect 241440 326 241560 354
rect 241440 134 241468 326
rect 241428 128 241480 134
rect 240856 66 241192 82
rect 241428 70 241480 76
rect 240856 60 241204 66
rect 240856 54 241152 60
rect 241152 2 241204 8
rect 241674 -960 241786 480
rect 241960 462 242254 490
rect 242912 480 242940 614
rect 246468 598 246804 626
rect 247664 620 247960 626
rect 253480 672 253532 678
rect 249062 640 249118 649
rect 247664 614 248012 620
rect 247664 598 248000 614
rect 248768 598 249062 626
rect 244094 575 244150 584
rect 244108 480 244136 575
rect 244936 564 245240 592
rect 244556 536 244608 542
rect 244260 484 244556 490
rect 242254 439 242310 448
rect 242870 -960 242982 480
rect 243064 338 243400 354
rect 243064 332 243412 338
rect 243064 326 243360 332
rect 243360 274 243412 280
rect 244066 -960 244178 480
rect 244260 478 244608 484
rect 244260 462 244596 478
rect 244936 474 244964 564
rect 245212 480 245240 564
rect 244924 468 244976 474
rect 244924 410 244976 416
rect 245170 -960 245282 480
rect 245660 400 245712 406
rect 245364 348 245660 354
rect 245364 342 245712 348
rect 245364 326 245700 342
rect 246366 82 246478 480
rect 246776 474 246804 598
rect 252172 610 252324 626
rect 249062 575 249118 584
rect 249984 604 250036 610
rect 249984 546 250036 552
rect 251180 604 251232 610
rect 252172 604 252336 610
rect 252172 598 252284 604
rect 251180 546 251232 552
rect 252284 546 252336 552
rect 252388 598 252600 626
rect 255780 672 255832 678
rect 254674 640 254730 649
rect 253480 614 253532 620
rect 247314 504 247370 513
rect 246764 468 246816 474
rect 249996 480 250024 546
rect 250902 504 250958 513
rect 247314 439 247370 448
rect 246764 410 246816 416
rect 247328 218 247356 439
rect 247562 218 247674 480
rect 247328 190 247674 218
rect 246040 66 246478 82
rect 246028 60 246478 66
rect 246080 54 246478 60
rect 246028 2 246080 8
rect 246366 -960 246478 54
rect 247562 -960 247674 190
rect 248758 354 248870 480
rect 248758 338 249012 354
rect 249720 338 249872 354
rect 248758 332 249024 338
rect 248758 326 248972 332
rect 248758 -960 248870 326
rect 248972 274 249024 280
rect 249708 332 249872 338
rect 249760 326 249872 332
rect 249708 274 249760 280
rect 249954 -960 250066 480
rect 250958 462 251068 490
rect 251192 480 251220 546
rect 252388 480 252416 598
rect 250902 439 250958 448
rect 251150 -960 251262 480
rect 252346 -960 252458 480
rect 252572 474 252600 598
rect 253492 480 253520 614
rect 254472 610 254624 626
rect 254472 604 254636 610
rect 254472 598 254584 604
rect 254674 575 254730 584
rect 255226 640 255282 649
rect 255576 620 255780 626
rect 261760 672 261812 678
rect 255576 614 255832 620
rect 255870 640 255926 649
rect 255576 598 255820 614
rect 255226 575 255282 584
rect 255870 575 255926 584
rect 257066 640 257122 649
rect 257066 575 257122 584
rect 258092 598 258304 626
rect 262680 672 262732 678
rect 261760 614 261812 620
rect 262384 620 262680 626
rect 268844 672 268896 678
rect 267278 640 267334 649
rect 262384 614 262732 620
rect 254584 546 254636 552
rect 254688 480 254716 575
rect 252560 468 252612 474
rect 252560 410 252612 416
rect 253112 400 253164 406
rect 253164 348 253276 354
rect 253112 342 253276 348
rect 253124 326 253276 342
rect 253450 -960 253562 480
rect 254646 -960 254758 480
rect 255240 338 255268 575
rect 255884 480 255912 575
rect 257080 480 257108 575
rect 258092 542 258120 598
rect 258080 536 258132 542
rect 255228 332 255280 338
rect 255228 274 255280 280
rect 255842 -960 255954 480
rect 256772 338 256924 354
rect 256772 332 256936 338
rect 256772 326 256884 332
rect 256884 274 256936 280
rect 257038 -960 257150 480
rect 258080 478 258132 484
rect 258276 480 258304 598
rect 260656 604 260708 610
rect 259288 564 259500 592
rect 259288 490 259316 564
rect 257876 202 258028 218
rect 257876 196 258040 202
rect 257876 190 257988 196
rect 257988 138 258040 144
rect 258234 -960 258346 480
rect 259104 474 259316 490
rect 259472 480 259500 564
rect 260656 546 260708 552
rect 260472 536 260524 542
rect 260176 484 260472 490
rect 259092 468 259316 474
rect 259144 462 259316 468
rect 259092 410 259144 416
rect 259276 400 259328 406
rect 258980 348 259276 354
rect 258980 342 259328 348
rect 258980 326 259316 342
rect 259430 -960 259542 480
rect 260176 478 260524 484
rect 260668 480 260696 546
rect 261576 536 261628 542
rect 261280 484 261576 490
rect 260176 462 260512 478
rect 260626 -960 260738 480
rect 261280 478 261628 484
rect 261772 480 261800 614
rect 262384 598 262720 614
rect 266544 604 266596 610
rect 262784 564 262996 592
rect 261280 462 261616 478
rect 261730 -960 261842 480
rect 262784 338 262812 564
rect 262968 480 262996 564
rect 263980 564 264192 592
rect 262772 332 262824 338
rect 262772 274 262824 280
rect 262926 -960 263038 480
rect 263580 474 263732 490
rect 263580 468 263744 474
rect 263580 462 263692 468
rect 263692 410 263744 416
rect 263980 354 264008 564
rect 264164 480 264192 564
rect 265176 564 265388 592
rect 265176 490 265204 564
rect 263888 326 264008 354
rect 263888 202 263916 326
rect 263876 196 263928 202
rect 263876 138 263928 144
rect 264122 -960 264234 480
rect 264992 462 265204 490
rect 265360 480 265388 564
rect 266984 598 267278 626
rect 275836 672 275888 678
rect 273626 640 273682 649
rect 268844 614 268896 620
rect 267278 575 267334 584
rect 267740 604 267792 610
rect 266544 546 266596 552
rect 267740 546 267792 552
rect 266556 480 266584 546
rect 267752 480 267780 546
rect 268384 536 268436 542
rect 268088 484 268384 490
rect 264992 406 265020 462
rect 264980 400 265032 406
rect 264980 342 265032 348
rect 264888 264 264940 270
rect 264684 212 264888 218
rect 264684 206 264940 212
rect 264684 190 264928 206
rect 265318 -960 265430 480
rect 266084 128 266136 134
rect 265788 76 266084 82
rect 265788 70 266136 76
rect 265788 54 266124 70
rect 266514 -960 266626 480
rect 267710 -960 267822 480
rect 268088 478 268436 484
rect 268856 480 268884 614
rect 270040 604 270092 610
rect 270040 546 270092 552
rect 271064 598 271276 626
rect 271492 610 271828 626
rect 271492 604 271840 610
rect 271492 598 271788 604
rect 269486 504 269542 513
rect 268088 462 268424 478
rect 268814 -960 268926 480
rect 269192 462 269486 490
rect 270052 480 270080 546
rect 269486 439 269542 448
rect 270010 -960 270122 480
rect 270388 474 270724 490
rect 270388 468 270736 474
rect 270388 462 270684 468
rect 270684 410 270736 416
rect 271064 270 271092 598
rect 271248 480 271276 598
rect 271788 546 271840 552
rect 272260 564 272472 592
rect 275190 640 275246 649
rect 274896 598 275190 626
rect 273626 575 273682 584
rect 277492 672 277544 678
rect 275888 620 276000 626
rect 275836 614 276000 620
rect 275848 598 276000 614
rect 277196 620 277492 626
rect 284300 672 284352 678
rect 278594 640 278650 649
rect 277196 614 277544 620
rect 277196 598 277532 614
rect 278300 598 278594 626
rect 275190 575 275246 584
rect 281704 610 281856 626
rect 278594 575 278650 584
rect 279516 604 279568 610
rect 271052 264 271104 270
rect 271052 206 271104 212
rect 271206 -960 271318 480
rect 272260 354 272288 564
rect 272444 480 272472 564
rect 273640 480 273668 575
rect 279516 546 279568 552
rect 280712 604 280764 610
rect 281704 604 281868 610
rect 281704 598 281816 604
rect 280712 546 280764 552
rect 281816 546 281868 552
rect 281920 598 282132 626
rect 286600 672 286652 678
rect 284300 614 284352 620
rect 285402 640 285458 649
rect 274548 536 274600 542
rect 278504 536 278556 542
rect 272168 326 272288 354
rect 272168 134 272196 326
rect 272156 128 272208 134
rect 272156 70 272208 76
rect 272402 -960 272514 480
rect 272892 400 272944 406
rect 272596 348 272892 354
rect 272596 342 272944 348
rect 272596 326 272932 342
rect 273598 -960 273710 480
rect 274548 478 274600 484
rect 276202 504 276258 513
rect 274560 354 274588 478
rect 274794 354 274906 480
rect 274560 326 274906 354
rect 273792 202 274128 218
rect 273792 196 274140 202
rect 273792 190 274088 196
rect 274088 138 274140 144
rect 274794 -960 274906 326
rect 275990 218 276102 480
rect 276202 439 276258 448
rect 276756 468 276808 474
rect 276216 218 276244 439
rect 276756 410 276808 416
rect 276768 354 276796 410
rect 277094 354 277206 480
rect 276768 326 277206 354
rect 275990 190 276244 218
rect 275990 -960 276102 190
rect 277094 -960 277206 326
rect 278290 354 278402 480
rect 278504 478 278556 484
rect 279528 480 279556 546
rect 278516 354 278544 478
rect 278290 326 278544 354
rect 279252 338 279404 354
rect 279240 332 279404 338
rect 278290 -960 278402 326
rect 279292 326 279404 332
rect 279240 274 279292 280
rect 279486 -960 279598 480
rect 280448 474 280600 490
rect 280724 480 280752 546
rect 281920 480 281948 598
rect 282104 513 282132 598
rect 283104 604 283156 610
rect 283104 546 283156 552
rect 282090 504 282146 513
rect 280436 468 280600 474
rect 280488 462 280600 468
rect 280436 410 280488 416
rect 280682 -960 280794 480
rect 281878 -960 281990 480
rect 283116 480 283144 546
rect 284312 480 284340 614
rect 285402 575 285458 584
rect 285678 640 285734 649
rect 288992 672 289044 678
rect 286600 614 286652 620
rect 287794 640 287850 649
rect 285678 575 285734 584
rect 285218 504 285274 513
rect 282090 439 282146 448
rect 282920 264 282972 270
rect 282808 212 282920 218
rect 282808 206 282972 212
rect 282808 190 282960 206
rect 283074 -960 283186 480
rect 284004 202 284156 218
rect 284004 196 284168 202
rect 284004 190 284116 196
rect 284116 138 284168 144
rect 284270 -960 284382 480
rect 285108 462 285218 490
rect 285416 480 285444 575
rect 285218 439 285274 448
rect 285374 -960 285486 480
rect 285692 474 285720 575
rect 286612 480 286640 614
rect 288512 610 288848 626
rect 291108 672 291160 678
rect 288992 614 289044 620
rect 288512 604 288860 610
rect 288512 598 288808 604
rect 287794 575 287850 584
rect 285680 468 285732 474
rect 285680 410 285732 416
rect 286414 368 286470 377
rect 286304 326 286414 354
rect 286414 303 286470 312
rect 286570 -960 286682 480
rect 287408 474 287652 490
rect 287808 480 287836 575
rect 288808 546 288860 552
rect 289004 480 289032 614
rect 290016 598 290228 626
rect 290812 620 291108 626
rect 293408 672 293460 678
rect 292578 640 292634 649
rect 290812 614 291160 620
rect 290812 598 291148 614
rect 291212 598 291424 626
rect 287408 468 287664 474
rect 287408 462 287612 468
rect 287612 410 287664 416
rect 287766 -960 287878 480
rect 288962 -960 289074 480
rect 289708 338 289860 354
rect 289708 332 289872 338
rect 289708 326 289820 332
rect 289820 274 289872 280
rect 290016 270 290044 598
rect 290200 480 290228 598
rect 290004 264 290056 270
rect 290004 206 290056 212
rect 290158 -960 290270 480
rect 291212 202 291240 598
rect 291396 480 291424 598
rect 293112 620 293408 626
rect 298468 672 298520 678
rect 293866 640 293922 649
rect 293112 614 293460 620
rect 293112 598 293448 614
rect 293512 598 293724 626
rect 292578 575 292634 584
rect 292212 536 292264 542
rect 291916 484 292212 490
rect 291200 196 291252 202
rect 291200 138 291252 144
rect 291354 -960 291466 480
rect 291916 478 292264 484
rect 292592 480 292620 575
rect 291916 462 292252 478
rect 292550 -960 292662 480
rect 293406 368 293462 377
rect 293512 354 293540 598
rect 293696 480 293724 598
rect 293866 575 293922 584
rect 294878 640 294934 649
rect 295614 640 295670 649
rect 295320 598 295614 626
rect 294878 575 294934 584
rect 298468 614 298520 620
rect 300768 672 300820 678
rect 301320 672 301372 678
rect 300768 614 300820 620
rect 301024 620 301320 626
rect 307668 672 307720 678
rect 301024 614 301372 620
rect 303158 640 303214 649
rect 295614 575 295670 584
rect 296076 604 296128 610
rect 293462 326 293540 354
rect 293406 303 293462 312
rect 293654 -960 293766 480
rect 293880 474 293908 575
rect 294892 480 294920 575
rect 296076 546 296128 552
rect 297272 604 297324 610
rect 297272 546 297324 552
rect 296088 480 296116 546
rect 297284 480 297312 546
rect 298480 480 298508 614
rect 299664 604 299716 610
rect 299664 546 299716 552
rect 299676 480 299704 546
rect 300216 536 300268 542
rect 299920 484 300216 490
rect 293868 468 293920 474
rect 293868 410 293920 416
rect 294512 400 294564 406
rect 294216 348 294512 354
rect 294216 342 294564 348
rect 294216 326 294552 342
rect 294850 -960 294962 480
rect 296046 -960 296158 480
rect 296516 202 296852 218
rect 296516 196 296864 202
rect 296516 190 296812 196
rect 296812 138 296864 144
rect 297242 -960 297354 480
rect 297620 338 297956 354
rect 297620 332 297968 338
rect 297620 326 297916 332
rect 297916 274 297968 280
rect 298438 -960 298550 480
rect 299020 128 299072 134
rect 298724 76 299020 82
rect 298724 70 299072 76
rect 298724 54 299060 70
rect 299634 -960 299746 480
rect 299920 478 300268 484
rect 300780 480 300808 614
rect 301024 598 301360 614
rect 301964 604 302016 610
rect 305826 640 305882 649
rect 304428 598 304764 626
rect 305532 598 305826 626
rect 303158 575 303214 584
rect 301964 546 302016 552
rect 301976 480 302004 546
rect 303172 480 303200 575
rect 303802 504 303858 513
rect 299920 462 300256 478
rect 300738 -960 300850 480
rect 301934 -960 302046 480
rect 302424 264 302476 270
rect 302128 212 302424 218
rect 302128 206 302476 212
rect 302128 190 302464 206
rect 303130 -960 303242 480
rect 303324 474 303660 490
rect 303324 468 303672 474
rect 303324 462 303620 468
rect 303802 439 303858 448
rect 303620 410 303672 416
rect 303816 134 303844 439
rect 304326 218 304438 480
rect 304736 406 304764 598
rect 306728 598 307064 626
rect 309048 672 309100 678
rect 307720 620 307832 626
rect 307668 614 307832 620
rect 307680 598 307832 614
rect 307956 610 308076 626
rect 311348 672 311400 678
rect 309048 614 309100 620
rect 311236 620 311348 626
rect 315948 672 316000 678
rect 311236 614 311400 620
rect 313830 640 313886 649
rect 307956 604 308088 610
rect 307956 598 308036 604
rect 305826 575 305882 584
rect 306930 504 306986 513
rect 304724 400 304776 406
rect 304724 342 304776 348
rect 305522 354 305634 480
rect 304000 202 304438 218
rect 303988 196 304438 202
rect 304040 190 304438 196
rect 303988 138 304040 144
rect 303804 128 303856 134
rect 303804 70 303856 76
rect 304326 -960 304438 190
rect 305522 338 305776 354
rect 305522 332 305788 338
rect 305522 326 305736 332
rect 305522 -960 305634 326
rect 305736 274 305788 280
rect 306718 218 306830 480
rect 306930 439 306986 448
rect 306944 218 306972 439
rect 307036 338 307064 598
rect 307956 480 307984 598
rect 308036 546 308088 552
rect 308772 536 308824 542
rect 308824 484 308936 490
rect 307024 332 307076 338
rect 307024 274 307076 280
rect 306718 190 306972 218
rect 306718 -960 306830 190
rect 307914 -960 308026 480
rect 308772 478 308936 484
rect 309060 480 309088 614
rect 310244 604 310296 610
rect 311236 598 311388 614
rect 311440 604 311492 610
rect 310244 546 310296 552
rect 311440 546 311492 552
rect 312636 604 312688 610
rect 315836 620 315948 626
rect 318340 672 318392 678
rect 315836 614 316000 620
rect 315836 598 315988 614
rect 316052 598 316264 626
rect 318044 620 318340 626
rect 326804 672 326856 678
rect 318044 614 318392 620
rect 318522 640 318578 649
rect 313830 575 313886 584
rect 312636 546 312688 552
rect 309966 504 310022 513
rect 308784 462 308936 478
rect 309018 -960 309130 480
rect 310022 462 310132 490
rect 310256 480 310284 546
rect 311452 480 311480 546
rect 309966 439 310022 448
rect 310214 -960 310326 480
rect 311410 -960 311522 480
rect 312340 474 312492 490
rect 312648 480 312676 546
rect 313844 480 313872 575
rect 314856 564 315068 592
rect 312340 468 312504 474
rect 312340 462 312452 468
rect 312452 410 312504 416
rect 312606 -960 312718 480
rect 313536 338 313688 354
rect 313536 332 313700 338
rect 313536 326 313648 332
rect 313648 274 313700 280
rect 313802 -960 313914 480
rect 314856 406 314884 564
rect 315040 480 315068 564
rect 316052 542 316080 598
rect 316040 536 316092 542
rect 314844 400 314896 406
rect 314844 342 314896 348
rect 314640 66 314792 82
rect 314640 60 314804 66
rect 314640 54 314752 60
rect 314752 2 314804 8
rect 314998 -960 315110 480
rect 316040 478 316092 484
rect 316236 480 316264 598
rect 317328 604 317380 610
rect 318044 598 318380 614
rect 318522 575 318578 584
rect 318890 640 318946 649
rect 318890 575 318946 584
rect 319718 640 319774 649
rect 326048 610 326384 626
rect 327448 672 327500 678
rect 326804 614 326856 620
rect 327152 620 327448 626
rect 339776 672 339828 678
rect 334898 640 334954 649
rect 327152 614 327500 620
rect 324412 604 324464 610
rect 319718 575 319774 584
rect 317328 546 317380 552
rect 317144 536 317196 542
rect 316940 484 317144 490
rect 316194 -960 316306 480
rect 316940 478 317196 484
rect 317340 480 317368 546
rect 318536 480 318564 575
rect 316940 462 317184 478
rect 317298 -960 317410 480
rect 318494 -960 318606 480
rect 318904 406 318932 575
rect 319732 480 319760 575
rect 320744 564 320956 592
rect 318892 400 318944 406
rect 318892 342 318944 348
rect 319444 264 319496 270
rect 319240 212 319444 218
rect 319240 206 319496 212
rect 319240 190 319484 206
rect 319690 -960 319802 480
rect 320744 474 320772 564
rect 320928 480 320956 564
rect 321848 564 322152 592
rect 320732 468 320784 474
rect 320732 410 320784 416
rect 320344 202 320680 218
rect 320344 196 320692 202
rect 320344 190 320640 196
rect 320640 138 320692 144
rect 320886 -960 320998 480
rect 321848 474 321876 564
rect 322124 480 322152 564
rect 323136 564 323348 592
rect 321836 468 321888 474
rect 321836 410 321888 416
rect 321560 264 321612 270
rect 321448 212 321560 218
rect 321448 206 321612 212
rect 321448 190 321600 206
rect 322082 -960 322194 480
rect 322848 128 322900 134
rect 322644 76 322848 82
rect 323136 82 323164 564
rect 323320 480 323348 564
rect 324412 546 324464 552
rect 325608 604 325660 610
rect 326048 604 326396 610
rect 326048 598 326344 604
rect 325608 546 325660 552
rect 326344 546 326396 552
rect 324424 480 324452 546
rect 322644 70 322900 76
rect 322644 54 322888 70
rect 322952 66 323164 82
rect 322940 60 323164 66
rect 322992 54 323164 60
rect 322940 2 322992 8
rect 323278 -960 323390 480
rect 323748 66 324084 82
rect 323748 60 324096 66
rect 323748 54 324044 60
rect 324044 2 324096 8
rect 324382 -960 324494 480
rect 324852 474 325188 490
rect 325620 480 325648 546
rect 326816 480 326844 614
rect 327152 598 327488 614
rect 327828 598 328040 626
rect 324852 468 325200 474
rect 324852 462 325148 468
rect 325148 410 325200 416
rect 325578 -960 325690 480
rect 326774 -960 326886 480
rect 327828 406 327856 598
rect 328012 480 328040 598
rect 329024 598 329236 626
rect 327816 400 327868 406
rect 327816 342 327868 348
rect 327970 -960 328082 480
rect 328458 232 328514 241
rect 328256 190 328458 218
rect 329024 202 329052 598
rect 329208 480 329236 598
rect 330220 598 330432 626
rect 331660 598 331996 626
rect 330220 490 330248 598
rect 328458 167 328514 176
rect 329012 196 329064 202
rect 329012 138 329064 144
rect 329166 -960 329278 480
rect 330128 462 330248 490
rect 330404 480 330432 598
rect 330128 270 330156 462
rect 330116 264 330168 270
rect 329452 202 329788 218
rect 330116 206 330168 212
rect 329452 196 329800 202
rect 329452 190 329748 196
rect 329748 138 329800 144
rect 330362 -960 330474 480
rect 330556 474 330892 490
rect 330556 468 330904 474
rect 330556 462 330852 468
rect 330852 410 330904 416
rect 331220 128 331272 134
rect 331558 82 331670 480
rect 331968 134 331996 598
rect 332520 598 332732 626
rect 333960 598 334296 626
rect 331272 76 331670 82
rect 331220 70 331670 76
rect 331956 128 332008 134
rect 331956 70 332008 76
rect 331232 54 331670 70
rect 332520 66 332548 598
rect 332704 480 332732 598
rect 331558 -960 331670 54
rect 332508 60 332560 66
rect 332508 2 332560 8
rect 332662 -960 332774 480
rect 333612 400 333664 406
rect 333858 354 333970 480
rect 333664 348 333970 354
rect 333612 342 333970 348
rect 333624 326 333970 342
rect 334268 338 334296 598
rect 334954 598 335064 626
rect 335268 604 335320 610
rect 334898 575 334954 584
rect 336260 598 336596 626
rect 339664 620 339776 626
rect 343180 672 343232 678
rect 339664 614 339828 620
rect 335268 546 335320 552
rect 332856 66 333192 82
rect 332856 60 333204 66
rect 332856 54 333152 60
rect 333152 2 333204 8
rect 333858 -960 333970 326
rect 334256 332 334308 338
rect 334256 274 334308 280
rect 335054 218 335166 480
rect 335280 218 335308 546
rect 336464 536 336516 542
rect 335054 190 335308 218
rect 336250 354 336362 480
rect 336464 478 336516 484
rect 336476 354 336504 478
rect 336568 406 336596 598
rect 336648 604 336700 610
rect 336648 546 336700 552
rect 337476 604 337528 610
rect 337476 546 337528 552
rect 338672 604 338724 610
rect 339664 598 339816 614
rect 339868 604 339920 610
rect 338672 546 338724 552
rect 339868 546 339920 552
rect 340972 604 341024 610
rect 340972 546 341024 552
rect 342180 598 342392 626
rect 343068 620 343180 626
rect 352840 672 352892 678
rect 343068 614 343232 620
rect 344558 640 344614 649
rect 343068 598 343220 614
rect 336250 326 336504 354
rect 336556 400 336608 406
rect 336556 342 336608 348
rect 335054 -960 335166 190
rect 336250 -960 336362 326
rect 336660 241 336688 546
rect 337200 536 337252 542
rect 337252 484 337364 490
rect 337200 478 337364 484
rect 337488 480 337516 546
rect 338302 504 338358 513
rect 337212 462 337364 478
rect 336646 232 336702 241
rect 336646 167 336702 176
rect 337446 -960 337558 480
rect 338358 462 338468 490
rect 338684 480 338712 546
rect 339880 480 339908 546
rect 338302 439 338358 448
rect 338642 -960 338754 480
rect 339838 -960 339950 480
rect 340616 474 340768 490
rect 340984 480 341012 546
rect 342180 480 342208 598
rect 340604 468 340768 474
rect 340656 462 340768 468
rect 340604 410 340656 416
rect 340942 -960 341054 480
rect 341800 128 341852 134
rect 341852 76 341964 82
rect 341800 70 341964 76
rect 341812 54 341964 70
rect 342138 -960 342250 480
rect 342364 66 342392 598
rect 343376 564 343588 592
rect 344558 575 344614 584
rect 344742 640 344798 649
rect 344742 575 344798 584
rect 345754 640 345810 649
rect 350170 640 350226 649
rect 345754 575 345810 584
rect 346780 598 346992 626
rect 343376 480 343404 564
rect 343560 524 343588 564
rect 343560 496 343634 524
rect 343606 490 343634 496
rect 342352 60 342404 66
rect 342352 2 342404 8
rect 343334 -960 343446 480
rect 343606 462 343680 490
rect 344572 480 344600 575
rect 343652 338 343680 462
rect 343640 332 343692 338
rect 343640 274 343692 280
rect 344172 202 344416 218
rect 344172 196 344428 202
rect 344172 190 344376 196
rect 344376 138 344428 144
rect 344530 -960 344642 480
rect 344756 406 344784 575
rect 345768 480 345796 575
rect 346780 542 346808 598
rect 346768 536 346820 542
rect 344744 400 344796 406
rect 344744 342 344796 348
rect 345572 400 345624 406
rect 345572 342 345624 348
rect 345584 218 345612 342
rect 345368 190 345612 218
rect 345726 -960 345838 480
rect 346768 478 346820 484
rect 346964 480 346992 598
rect 347884 598 348096 626
rect 347688 536 347740 542
rect 347576 484 347688 490
rect 347884 513 347912 598
rect 346768 264 346820 270
rect 346472 212 346768 218
rect 346472 206 346820 212
rect 346472 190 346808 206
rect 346922 -960 347034 480
rect 347576 478 347740 484
rect 347870 504 347926 513
rect 347576 462 347728 478
rect 348068 480 348096 598
rect 349252 604 349304 610
rect 349876 598 350170 626
rect 352562 640 352618 649
rect 350170 575 350226 584
rect 350276 598 350488 626
rect 349252 546 349304 552
rect 348422 504 348478 513
rect 347870 439 347926 448
rect 348026 -960 348138 480
rect 349264 480 349292 546
rect 350276 513 350304 598
rect 350262 504 350318 513
rect 348422 439 348424 448
rect 348476 439 348478 448
rect 348424 410 348476 416
rect 348772 66 349108 82
rect 348772 60 349120 66
rect 348772 54 349068 60
rect 349068 2 349120 8
rect 349222 -960 349334 480
rect 350460 480 350488 598
rect 351472 598 351684 626
rect 350262 439 350318 448
rect 349434 232 349490 241
rect 349434 167 349490 176
rect 349448 134 349476 167
rect 349436 128 349488 134
rect 349436 70 349488 76
rect 350418 -960 350530 480
rect 350980 338 351316 354
rect 350980 332 351328 338
rect 350980 326 351276 332
rect 351276 274 351328 280
rect 351472 241 351500 598
rect 351656 480 351684 598
rect 359280 672 359332 678
rect 352840 614 352892 620
rect 354034 640 354090 649
rect 352562 575 352618 584
rect 352472 536 352524 542
rect 352176 484 352472 490
rect 351458 232 351514 241
rect 351458 167 351514 176
rect 351614 -960 351726 480
rect 352176 478 352524 484
rect 352176 462 352512 478
rect 352576 202 352604 575
rect 352852 480 352880 614
rect 354034 575 354090 584
rect 355060 598 355272 626
rect 352564 196 352616 202
rect 352564 138 352616 144
rect 352810 -960 352922 480
rect 353280 474 353616 490
rect 354048 480 354076 575
rect 354680 536 354732 542
rect 354384 484 354680 490
rect 353280 468 353628 474
rect 353280 462 353576 468
rect 353576 410 353628 416
rect 354006 -960 354118 480
rect 354384 478 354732 484
rect 354384 462 354720 478
rect 355060 406 355088 598
rect 355244 480 355272 598
rect 356072 598 356376 626
rect 355048 400 355100 406
rect 355048 342 355100 348
rect 355202 -960 355314 480
rect 356072 270 356100 598
rect 356348 480 356376 598
rect 357532 604 357584 610
rect 357532 546 357584 552
rect 358556 598 358768 626
rect 358984 620 359280 626
rect 360384 672 360436 678
rect 358984 614 359332 620
rect 359922 640 359978 649
rect 358984 598 359320 614
rect 357544 480 357572 546
rect 356060 264 356112 270
rect 355580 202 355916 218
rect 356060 206 356112 212
rect 355580 196 355928 202
rect 355580 190 355876 196
rect 355876 138 355928 144
rect 356306 -960 356418 480
rect 356980 400 357032 406
rect 356684 348 356980 354
rect 356684 342 357032 348
rect 356684 326 357020 342
rect 357502 -960 357614 480
rect 358556 354 358584 598
rect 358740 480 358768 598
rect 360088 620 360384 626
rect 363788 672 363840 678
rect 363786 640 363788 649
rect 366088 672 366140 678
rect 363840 640 363842 649
rect 360088 614 360436 620
rect 360088 598 360424 614
rect 361192 598 361528 626
rect 359922 575 359978 584
rect 359936 480 359964 575
rect 361500 542 361528 598
rect 361948 604 362000 610
rect 362388 598 362724 626
rect 363492 598 363736 626
rect 361948 546 362000 552
rect 361488 536 361540 542
rect 358464 326 358584 354
rect 358084 264 358136 270
rect 357788 212 358084 218
rect 357788 206 358136 212
rect 357788 190 358124 206
rect 358464 66 358492 326
rect 358452 60 358504 66
rect 358452 2 358504 8
rect 358698 -960 358810 480
rect 359894 -960 360006 480
rect 361090 354 361202 480
rect 361488 478 361540 484
rect 360856 338 361202 354
rect 360844 332 361202 338
rect 360896 326 361202 332
rect 361960 354 361988 546
rect 362286 354 362398 480
rect 361960 326 362398 354
rect 362696 338 362724 598
rect 363708 513 363736 598
rect 364596 598 364932 626
rect 365792 620 366088 626
rect 371608 672 371660 678
rect 365792 614 366140 620
rect 370594 640 370650 649
rect 365792 598 366128 614
rect 367008 604 367060 610
rect 363786 575 363842 584
rect 363694 504 363750 513
rect 360844 274 360896 280
rect 361090 -960 361202 326
rect 362286 -960 362398 326
rect 362684 332 362736 338
rect 362684 274 362736 280
rect 363482 82 363594 480
rect 363694 439 363750 448
rect 364586 354 364698 480
rect 364800 468 364852 474
rect 364800 410 364852 416
rect 364812 354 364840 410
rect 364586 326 364840 354
rect 363696 128 363748 134
rect 363482 76 363696 82
rect 363482 70 363748 76
rect 363482 54 363736 70
rect 363482 -960 363594 54
rect 364586 -960 364698 326
rect 364904 270 364932 598
rect 367008 546 367060 552
rect 368204 604 368256 610
rect 368204 546 368256 552
rect 369400 604 369452 610
rect 371496 620 371608 626
rect 373908 672 373960 678
rect 371496 614 371660 620
rect 373704 620 373908 626
rect 382372 672 382424 678
rect 373704 614 373960 620
rect 374090 640 374146 649
rect 371496 598 371648 614
rect 371700 604 371752 610
rect 370594 575 370650 584
rect 369400 546 369452 552
rect 367020 480 367048 546
rect 368216 480 368244 546
rect 369412 480 369440 546
rect 370608 480 370636 575
rect 373704 598 373948 614
rect 371700 546 371752 552
rect 372908 564 373120 592
rect 374090 575 374146 584
rect 374274 640 374330 649
rect 374274 575 374330 584
rect 375286 640 375342 649
rect 375286 575 375342 584
rect 375470 640 375526 649
rect 378874 640 378930 649
rect 375470 575 375526 584
rect 376484 604 376536 610
rect 371712 480 371740 546
rect 364982 368 365038 377
rect 364982 303 364984 312
rect 365036 303 365038 312
rect 364984 274 365036 280
rect 364892 264 364944 270
rect 364892 206 364944 212
rect 365782 218 365894 480
rect 365782 202 366036 218
rect 365782 196 366048 202
rect 365782 190 365996 196
rect 365782 -960 365894 190
rect 365996 138 366048 144
rect 366732 128 366784 134
rect 366784 76 366896 82
rect 366732 70 366896 76
rect 366744 54 366896 70
rect 366978 -960 367090 480
rect 367848 202 368000 218
rect 367836 196 368000 202
rect 367888 190 368000 196
rect 367836 138 367888 144
rect 368174 -960 368286 480
rect 369044 66 369196 82
rect 369032 60 369196 66
rect 369084 54 369196 60
rect 369032 2 369084 8
rect 369370 -960 369482 480
rect 370412 400 370464 406
rect 370300 348 370412 354
rect 370300 342 370464 348
rect 370300 326 370452 342
rect 370566 -960 370678 480
rect 371670 -960 371782 480
rect 372600 474 372752 490
rect 372908 480 372936 564
rect 372600 468 372764 474
rect 372600 462 372712 468
rect 372712 410 372764 416
rect 372866 -960 372978 480
rect 373092 377 373120 564
rect 374104 480 374132 575
rect 373078 368 373134 377
rect 373078 303 373134 312
rect 374062 -960 374174 480
rect 374288 270 374316 575
rect 374368 536 374420 542
rect 374366 504 374368 513
rect 374420 504 374422 513
rect 375300 480 375328 575
rect 374366 439 374422 448
rect 374276 264 374328 270
rect 375104 264 375156 270
rect 374276 206 374328 212
rect 374900 212 375104 218
rect 374900 206 375156 212
rect 374900 190 375144 206
rect 375258 -960 375370 480
rect 375484 202 375512 575
rect 376484 546 376536 552
rect 377508 564 377720 592
rect 378874 575 378930 584
rect 379058 640 379114 649
rect 381174 640 381230 649
rect 379408 610 379560 626
rect 379408 604 379572 610
rect 379408 598 379520 604
rect 379058 575 379114 584
rect 376496 480 376524 546
rect 377404 536 377456 542
rect 377108 484 377404 490
rect 377508 513 377536 564
rect 376004 338 376340 354
rect 376004 332 376352 338
rect 376004 326 376300 332
rect 376300 274 376352 280
rect 375472 196 375524 202
rect 375472 138 375524 144
rect 376454 -960 376566 480
rect 377108 478 377456 484
rect 377494 504 377550 513
rect 377108 462 377444 478
rect 377692 480 377720 564
rect 378888 480 378916 575
rect 377494 439 377550 448
rect 376758 96 376814 105
rect 376758 31 376760 40
rect 376812 31 376814 40
rect 376760 2 376812 8
rect 377650 -960 377762 480
rect 378304 66 378640 82
rect 378304 60 378652 66
rect 378304 54 378600 60
rect 378600 2 378652 8
rect 378846 -960 378958 480
rect 379072 406 379100 575
rect 379520 546 379572 552
rect 379808 564 380020 592
rect 383108 672 383160 678
rect 382372 614 382424 620
rect 382812 620 383108 626
rect 390284 672 390336 678
rect 382812 614 383160 620
rect 383566 640 383622 649
rect 381174 575 381230 584
rect 379610 504 379666 513
rect 379610 439 379612 448
rect 379664 439 379666 448
rect 379612 410 379664 416
rect 379060 400 379112 406
rect 379060 342 379112 348
rect 379808 105 379836 564
rect 379992 480 380020 564
rect 381188 480 381216 575
rect 382004 536 382056 542
rect 379794 96 379850 105
rect 379794 31 379850 40
rect 379950 -960 380062 480
rect 380512 202 380848 218
rect 380512 196 380860 202
rect 380512 190 380808 196
rect 380808 138 380860 144
rect 381146 -960 381258 480
rect 382004 478 382056 484
rect 382384 480 382412 614
rect 382812 598 383148 614
rect 383566 575 383622 584
rect 384592 598 384804 626
rect 383580 480 383608 575
rect 384210 504 384266 513
rect 381912 400 381964 406
rect 381708 348 381912 354
rect 381708 342 381964 348
rect 381708 326 381952 342
rect 382016 241 382044 478
rect 382002 232 382058 241
rect 382002 167 382058 176
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 383916 462 384210 490
rect 384210 439 384266 448
rect 384592 241 384620 598
rect 384776 480 384804 598
rect 385960 604 386012 610
rect 385960 546 386012 552
rect 386984 598 387196 626
rect 385972 480 386000 546
rect 384578 232 384634 241
rect 384578 167 384634 176
rect 384734 -960 384846 480
rect 385408 128 385460 134
rect 385112 76 385408 82
rect 385112 70 385460 76
rect 385112 54 385448 70
rect 385930 -960 386042 480
rect 386984 338 387012 598
rect 387168 480 387196 598
rect 388260 604 388312 610
rect 388260 546 388312 552
rect 389284 598 389496 626
rect 392216 672 392268 678
rect 391018 640 391074 649
rect 390284 614 390336 620
rect 388272 480 388300 546
rect 388812 536 388864 542
rect 388516 484 388812 490
rect 386972 332 387024 338
rect 386972 274 387024 280
rect 386512 264 386564 270
rect 386216 212 386512 218
rect 386216 206 386564 212
rect 386216 190 386552 206
rect 387126 -960 387238 480
rect 387320 338 387656 354
rect 387320 332 387668 338
rect 387320 326 387616 332
rect 387616 274 387668 280
rect 388230 -960 388342 480
rect 388516 478 388864 484
rect 388516 462 388852 478
rect 389284 218 389312 598
rect 389468 480 389496 598
rect 389192 190 389312 218
rect 389192 66 389220 190
rect 389180 60 389232 66
rect 389180 2 389232 8
rect 389426 -960 389538 480
rect 390296 354 390324 614
rect 390724 598 391018 626
rect 391920 620 392216 626
rect 394240 672 394292 678
rect 391920 614 392268 620
rect 391920 598 392256 614
rect 393024 610 393360 626
rect 395620 672 395672 678
rect 394240 614 394292 620
rect 395324 620 395620 626
rect 403072 672 403124 678
rect 402518 640 402574 649
rect 395324 614 395672 620
rect 393024 604 393372 610
rect 393024 598 393320 604
rect 391018 575 391074 584
rect 393320 546 393372 552
rect 390622 354 390734 480
rect 390296 326 390734 354
rect 389620 66 389956 82
rect 389620 60 389968 66
rect 389620 54 389916 60
rect 389916 2 389968 8
rect 390622 -960 390734 326
rect 391818 218 391930 480
rect 391584 202 391930 218
rect 391572 196 391930 202
rect 391624 190 391930 196
rect 391572 138 391624 144
rect 391818 -960 391930 190
rect 393014 354 393126 480
rect 393976 474 394128 490
rect 394252 480 394280 614
rect 395324 598 395660 614
rect 396552 598 396764 626
rect 395526 504 395582 513
rect 393964 468 394128 474
rect 394016 462 394128 468
rect 393964 410 394016 416
rect 393228 400 393280 406
rect 393014 348 393228 354
rect 393014 342 393280 348
rect 393014 326 393268 342
rect 393014 -960 393126 326
rect 394210 -960 394322 480
rect 395314 354 395426 480
rect 396552 480 396580 598
rect 395526 439 395582 448
rect 395540 354 395568 439
rect 395314 326 395568 354
rect 395314 -960 395426 326
rect 396276 202 396428 218
rect 396264 196 396428 202
rect 396316 190 396428 196
rect 396264 138 396316 144
rect 396510 -960 396622 480
rect 396736 354 396764 598
rect 397748 598 398052 626
rect 397748 480 397776 598
rect 397460 400 397512 406
rect 396736 326 396856 354
rect 397512 348 397624 354
rect 397460 342 397624 348
rect 397472 326 397624 342
rect 396828 134 396856 326
rect 396816 128 396868 134
rect 396816 70 396868 76
rect 397706 -960 397818 480
rect 398024 270 398052 598
rect 398944 598 399248 626
rect 398944 480 398972 598
rect 398012 264 398064 270
rect 398012 206 398064 212
rect 398564 264 398616 270
rect 398616 212 398728 218
rect 398564 206 398728 212
rect 398576 190 398728 206
rect 398902 -960 399014 480
rect 399220 338 399248 598
rect 400128 604 400180 610
rect 400128 546 400180 552
rect 401336 598 401548 626
rect 400140 480 400168 546
rect 399208 332 399260 338
rect 399208 274 399260 280
rect 399832 66 399984 82
rect 399832 60 399996 66
rect 399832 54 399944 60
rect 399944 2 399996 8
rect 400098 -960 400210 480
rect 401028 474 401180 490
rect 401336 480 401364 598
rect 401028 468 401192 474
rect 401028 462 401140 468
rect 401140 410 401192 416
rect 401294 -960 401406 480
rect 401520 338 401548 598
rect 402518 575 402574 584
rect 403070 640 403072 649
rect 403440 672 403492 678
rect 403124 640 403126 649
rect 403236 620 403440 626
rect 407212 672 407264 678
rect 403236 614 403492 620
rect 403622 640 403678 649
rect 403236 598 403480 614
rect 403070 575 403126 584
rect 405646 640 405702 649
rect 405384 610 405536 626
rect 403622 575 403678 584
rect 404820 604 404872 610
rect 402532 480 402560 575
rect 403636 480 403664 575
rect 404820 546 404872 552
rect 405372 604 405536 610
rect 405424 598 405536 604
rect 405646 575 405702 584
rect 405844 598 406056 626
rect 408132 672 408184 678
rect 407212 614 407264 620
rect 407836 620 408132 626
rect 415492 672 415544 678
rect 407836 614 408184 620
rect 408406 640 408462 649
rect 405372 546 405424 552
rect 404832 480 404860 546
rect 402132 338 402376 354
rect 401508 332 401560 338
rect 402132 332 402388 338
rect 402132 326 402336 332
rect 401508 274 401560 280
rect 402336 274 402388 280
rect 402490 -960 402602 480
rect 403594 -960 403706 480
rect 404636 128 404688 134
rect 404432 76 404636 82
rect 404432 70 404688 76
rect 404432 54 404676 70
rect 404790 -960 404902 480
rect 405660 202 405688 575
rect 405844 406 405872 598
rect 406028 480 406056 598
rect 407224 480 407252 614
rect 407836 598 408172 614
rect 409602 640 409658 649
rect 408940 610 409276 626
rect 408940 604 409288 610
rect 408940 598 409236 604
rect 408406 575 408462 584
rect 407488 536 407540 542
rect 407486 504 407488 513
rect 407540 504 407542 513
rect 405832 400 405884 406
rect 405832 342 405884 348
rect 405648 196 405700 202
rect 405648 138 405700 144
rect 405986 -960 406098 480
rect 406640 202 406976 218
rect 406640 196 406988 202
rect 406640 190 406936 196
rect 406936 138 406988 144
rect 407182 -960 407294 480
rect 408420 480 408448 575
rect 409602 575 409658 584
rect 410536 598 410840 626
rect 409236 546 409288 552
rect 409616 480 409644 575
rect 407486 439 407542 448
rect 408378 -960 408490 480
rect 409574 -960 409686 480
rect 410340 400 410392 406
rect 410044 348 410340 354
rect 410044 342 410392 348
rect 410044 326 410380 342
rect 410536 270 410564 598
rect 410812 480 410840 598
rect 411732 598 411944 626
rect 412344 610 412680 626
rect 412344 604 412692 610
rect 412344 598 412640 604
rect 410524 264 410576 270
rect 410524 206 410576 212
rect 410770 -960 410882 480
rect 411732 354 411760 598
rect 411916 480 411944 598
rect 412640 546 412692 552
rect 412928 598 413140 626
rect 411640 326 411760 354
rect 411536 264 411588 270
rect 411240 212 411536 218
rect 411240 206 411588 212
rect 411240 190 411576 206
rect 411640 66 411668 326
rect 411628 60 411680 66
rect 411628 2 411680 8
rect 411874 -960 411986 480
rect 412928 474 412956 598
rect 413112 480 413140 598
rect 414032 598 414336 626
rect 421012 672 421064 678
rect 421010 640 421012 649
rect 421104 672 421156 678
rect 421064 640 421066 649
rect 415492 614 415544 620
rect 413744 536 413796 542
rect 413448 484 413744 490
rect 412916 468 412968 474
rect 412916 410 412968 416
rect 413070 -960 413182 480
rect 413448 478 413796 484
rect 413448 462 413784 478
rect 414032 338 414060 598
rect 414308 480 414336 598
rect 415504 480 415532 614
rect 416516 598 416728 626
rect 416852 610 417188 626
rect 416852 604 417200 610
rect 416852 598 417148 604
rect 416516 490 416544 598
rect 414020 332 414072 338
rect 414020 274 414072 280
rect 414266 -960 414378 480
rect 414940 264 414992 270
rect 414644 212 414940 218
rect 414644 206 414992 212
rect 414644 190 414980 206
rect 415462 -960 415574 480
rect 415748 474 416176 490
rect 415748 468 416188 474
rect 415748 462 416136 468
rect 416136 410 416188 416
rect 416424 462 416544 490
rect 416700 480 416728 598
rect 417148 546 417200 552
rect 417884 604 417936 610
rect 417884 546 417936 552
rect 418620 604 418672 610
rect 418620 546 418672 552
rect 418816 598 419028 626
rect 420256 610 420592 626
rect 417896 480 417924 546
rect 418632 513 418660 546
rect 418618 504 418674 513
rect 416424 134 416452 462
rect 416412 128 416464 134
rect 416412 70 416464 76
rect 416658 -960 416770 480
rect 417854 -960 417966 480
rect 418618 439 418674 448
rect 418344 400 418396 406
rect 418048 348 418344 354
rect 418048 342 418396 348
rect 418048 326 418384 342
rect 418816 202 418844 598
rect 419000 480 419028 598
rect 419908 604 419960 610
rect 420256 604 420604 610
rect 420256 598 420552 604
rect 419908 546 419960 552
rect 421748 672 421800 678
rect 421104 614 421156 620
rect 421452 620 421748 626
rect 426072 672 426124 678
rect 423770 640 423826 649
rect 421452 614 421800 620
rect 421010 575 421066 584
rect 420552 546 420604 552
rect 418804 196 418856 202
rect 418804 138 418856 144
rect 418958 -960 419070 480
rect 419152 338 419488 354
rect 419152 332 419500 338
rect 419152 326 419448 332
rect 419448 274 419500 280
rect 419920 218 419948 546
rect 420154 218 420266 480
rect 421116 354 421144 614
rect 421452 598 421788 614
rect 422404 598 422556 626
rect 421350 354 421462 480
rect 421116 326 421462 354
rect 419920 190 420266 218
rect 420154 -960 420266 190
rect 421350 -960 421462 326
rect 422404 66 422432 598
rect 423770 575 423826 584
rect 424966 640 425022 649
rect 425960 620 426072 626
rect 426348 672 426400 678
rect 425960 614 426124 620
rect 426176 620 426348 626
rect 426176 614 426400 620
rect 426992 672 427044 678
rect 427268 672 427320 678
rect 427044 620 427156 626
rect 426992 614 427156 620
rect 427912 672 427964 678
rect 427268 614 427320 620
rect 427910 640 427912 649
rect 428372 672 428424 678
rect 427964 640 427966 649
rect 425960 598 426112 614
rect 426176 598 426388 614
rect 427004 598 427156 614
rect 424966 575 425022 584
rect 422760 536 422812 542
rect 422546 354 422658 480
rect 422760 478 422812 484
rect 423784 480 423812 575
rect 424980 480 425008 575
rect 426176 480 426204 598
rect 427280 480 427308 614
rect 428260 620 428372 626
rect 431868 672 431920 678
rect 428260 614 428424 620
rect 429658 640 429714 649
rect 428260 598 428412 614
rect 428464 604 428516 610
rect 427910 575 427966 584
rect 431038 640 431094 649
rect 429658 575 429714 584
rect 430684 598 430896 626
rect 428464 546 428516 552
rect 428476 480 428504 546
rect 429476 536 429528 542
rect 429364 484 429476 490
rect 422772 354 422800 478
rect 422546 326 422800 354
rect 422392 60 422444 66
rect 422392 2 422444 8
rect 422546 -960 422658 326
rect 423508 202 423660 218
rect 423496 196 423660 202
rect 423548 190 423660 196
rect 423496 138 423548 144
rect 423742 -960 423854 480
rect 424692 128 424744 134
rect 424744 76 424856 82
rect 424692 70 424856 76
rect 424704 54 424856 70
rect 424938 -960 425050 480
rect 426134 -960 426246 480
rect 427238 -960 427350 480
rect 428434 -960 428546 480
rect 429364 478 429528 484
rect 429672 480 429700 575
rect 429364 462 429516 478
rect 429630 -960 429742 480
rect 430408 474 430560 490
rect 430396 468 430560 474
rect 430448 462 430560 468
rect 430396 410 430448 416
rect 430684 406 430712 598
rect 430868 480 430896 598
rect 431664 620 431868 626
rect 434444 672 434496 678
rect 431664 614 431920 620
rect 432050 640 432106 649
rect 431664 598 431908 614
rect 431038 575 431094 584
rect 441528 672 441580 678
rect 434444 614 434496 620
rect 432050 575 432106 584
rect 433248 604 433300 610
rect 430672 400 430724 406
rect 430672 342 430724 348
rect 430826 -960 430938 480
rect 431052 338 431080 575
rect 432064 480 432092 575
rect 433248 546 433300 552
rect 433260 480 433288 546
rect 434456 480 434484 614
rect 435548 604 435600 610
rect 435548 546 435600 552
rect 436572 598 436784 626
rect 435364 536 435416 542
rect 435068 484 435364 490
rect 431040 332 431092 338
rect 431040 274 431092 280
rect 432022 -960 432134 480
rect 433064 400 433116 406
rect 432768 348 433064 354
rect 432768 342 433116 348
rect 432768 326 433104 342
rect 433218 -960 433330 480
rect 433964 338 434300 354
rect 433964 332 434312 338
rect 433964 326 434260 332
rect 434260 274 434312 280
rect 434414 -960 434526 480
rect 435068 478 435416 484
rect 435560 480 435588 546
rect 435068 462 435404 478
rect 435518 -960 435630 480
rect 436572 354 436600 598
rect 436756 480 436784 598
rect 437768 598 437980 626
rect 438472 610 438808 626
rect 440772 610 441108 626
rect 442172 672 442224 678
rect 441528 614 441580 620
rect 441876 620 442172 626
rect 443276 672 443328 678
rect 441876 614 442224 620
rect 442980 620 443276 626
rect 445024 672 445076 678
rect 442980 614 443328 620
rect 438472 604 438820 610
rect 438472 598 438768 604
rect 436480 326 436600 354
rect 436480 202 436508 326
rect 436468 196 436520 202
rect 436468 138 436520 144
rect 436172 66 436508 82
rect 436172 60 436520 66
rect 436172 54 436468 60
rect 436468 2 436520 8
rect 436714 -960 436826 480
rect 437368 202 437520 218
rect 437368 196 437532 202
rect 437368 190 437480 196
rect 437480 138 437532 144
rect 437768 134 437796 598
rect 437952 480 437980 598
rect 438768 546 438820 552
rect 439136 604 439188 610
rect 439136 546 439188 552
rect 440332 604 440384 610
rect 440772 604 441120 610
rect 440772 598 441068 604
rect 440332 546 440384 552
rect 441068 546 441120 552
rect 439148 480 439176 546
rect 440344 480 440372 546
rect 441540 480 441568 614
rect 441876 598 442212 614
rect 442632 604 442684 610
rect 442980 598 443316 614
rect 443656 598 443868 626
rect 444176 610 444512 626
rect 445576 672 445628 678
rect 445024 614 445076 620
rect 445280 620 445576 626
rect 452384 672 452436 678
rect 445280 614 445628 620
rect 444176 604 444524 610
rect 444176 598 444472 604
rect 442632 546 442684 552
rect 442644 480 442672 546
rect 437756 128 437808 134
rect 437756 70 437808 76
rect 437910 -960 438022 480
rect 439106 -960 439218 480
rect 439872 264 439924 270
rect 439576 212 439872 218
rect 439576 206 439924 212
rect 439576 190 439912 206
rect 440302 -960 440414 480
rect 441498 -960 441610 480
rect 442602 -960 442714 480
rect 443656 474 443684 598
rect 443840 480 443868 598
rect 444472 546 444524 552
rect 445036 480 445064 614
rect 445280 598 445616 614
rect 446048 598 446260 626
rect 443644 468 443696 474
rect 443644 410 443696 416
rect 443798 -960 443910 480
rect 444994 -960 445106 480
rect 446048 406 446076 598
rect 446232 480 446260 598
rect 447152 598 447456 626
rect 448684 598 449020 626
rect 446036 400 446088 406
rect 446036 342 446088 348
rect 446190 -960 446302 480
rect 446384 474 446720 490
rect 446384 468 446732 474
rect 446384 462 446680 468
rect 446680 410 446732 416
rect 447152 338 447180 598
rect 447428 480 447456 598
rect 448244 536 448296 542
rect 447140 332 447192 338
rect 447140 274 447192 280
rect 447386 -960 447498 480
rect 448244 478 448296 484
rect 447876 400 447928 406
rect 447580 348 447876 354
rect 447580 342 447928 348
rect 448256 354 448284 478
rect 448582 354 448694 480
rect 447580 326 447916 342
rect 448256 326 448694 354
rect 448992 338 449020 598
rect 449636 598 449788 626
rect 450984 598 451320 626
rect 452088 620 452384 626
rect 454500 672 454552 678
rect 452088 614 452436 620
rect 452088 598 452424 614
rect 453284 598 453528 626
rect 457076 672 457128 678
rect 456062 640 456118 649
rect 454500 614 454552 620
rect 449636 542 449664 598
rect 449624 536 449676 542
rect 449624 478 449676 484
rect 449866 496 450032 524
rect 449866 480 449894 496
rect 448582 -960 448694 326
rect 448980 332 449032 338
rect 448980 274 449032 280
rect 449778 190 449894 480
rect 449778 -960 449890 190
rect 450004 66 450032 496
rect 450882 218 450994 480
rect 450648 202 450994 218
rect 450636 196 450994 202
rect 450688 190 450994 196
rect 450636 138 450688 144
rect 449992 60 450044 66
rect 449992 2 450044 8
rect 450882 -960 450994 190
rect 451292 134 451320 598
rect 452292 536 452344 542
rect 453500 513 453528 598
rect 452078 354 452190 480
rect 452292 478 452344 484
rect 453486 504 453542 513
rect 452304 354 452332 478
rect 452078 326 452332 354
rect 451280 128 451332 134
rect 451280 70 451332 76
rect 452078 -960 452190 326
rect 453274 218 453386 480
rect 454512 480 454540 614
rect 455492 610 455644 626
rect 455492 604 455656 610
rect 455492 598 455604 604
rect 455604 546 455656 552
rect 455708 598 455920 626
rect 455708 480 455736 598
rect 455892 542 455920 598
rect 456062 575 456118 584
rect 456904 632 457076 660
rect 455880 536 455932 542
rect 453486 439 453542 448
rect 453488 264 453540 270
rect 453274 212 453488 218
rect 453274 206 453540 212
rect 453274 190 453528 206
rect 453274 -960 453386 190
rect 454236 66 454388 82
rect 454224 60 454388 66
rect 454276 54 454388 60
rect 454224 2 454276 8
rect 454470 -960 454582 480
rect 455666 -960 455778 480
rect 455880 478 455932 484
rect 456076 474 456104 575
rect 456904 480 456932 632
rect 457996 672 458048 678
rect 457076 614 457128 620
rect 457792 620 457996 626
rect 458180 672 458232 678
rect 457792 614 458048 620
rect 458100 620 458180 626
rect 458100 614 458232 620
rect 459192 672 459244 678
rect 460296 672 460348 678
rect 459192 614 459244 620
rect 460092 620 460296 626
rect 461952 672 462004 678
rect 460092 614 460348 620
rect 460386 640 460442 649
rect 457792 598 458036 614
rect 458100 598 458220 614
rect 458100 480 458128 598
rect 459204 480 459232 614
rect 460092 598 460336 614
rect 460386 575 460442 584
rect 460938 640 460994 649
rect 461504 610 461624 626
rect 464712 672 464764 678
rect 461952 614 462004 620
rect 462778 640 462834 649
rect 460938 575 460994 584
rect 461492 604 461624 610
rect 460400 480 460428 575
rect 456064 468 456116 474
rect 456064 410 456116 416
rect 456536 338 456688 354
rect 456524 332 456688 338
rect 456576 326 456688 332
rect 456524 274 456576 280
rect 456862 -960 456974 480
rect 458058 -960 458170 480
rect 458896 66 459048 82
rect 458896 60 459060 66
rect 458896 54 459008 60
rect 459008 2 459060 8
rect 459162 -960 459274 480
rect 460358 -960 460470 480
rect 460952 202 460980 575
rect 461544 598 461624 604
rect 461492 546 461544 552
rect 461196 474 461440 490
rect 461596 480 461624 598
rect 461768 604 461820 610
rect 461768 546 461820 552
rect 461780 513 461808 546
rect 461964 513 461992 614
rect 462778 575 462834 584
rect 463974 640 464030 649
rect 464600 620 464712 626
rect 464600 614 464764 620
rect 466276 672 466328 678
rect 472256 672 472308 678
rect 466276 614 466328 620
rect 464600 598 464752 614
rect 463974 575 464030 584
rect 461766 504 461822 513
rect 461196 468 461452 474
rect 461196 462 461400 468
rect 461400 410 461452 416
rect 460940 196 460992 202
rect 460940 138 460992 144
rect 461554 -960 461666 480
rect 461766 439 461822 448
rect 461950 504 462006 513
rect 462792 480 462820 575
rect 463988 480 464016 575
rect 465000 564 465212 592
rect 461950 439 462006 448
rect 462412 264 462464 270
rect 462300 212 462412 218
rect 462300 206 462464 212
rect 462300 190 462452 206
rect 462750 -960 462862 480
rect 463496 202 463648 218
rect 463496 196 463660 202
rect 463496 190 463608 196
rect 463608 138 463660 144
rect 463946 -960 464058 480
rect 465000 406 465028 564
rect 465184 480 465212 564
rect 464988 400 465040 406
rect 464988 342 465040 348
rect 465142 -960 465254 480
rect 465704 474 466040 490
rect 466288 480 466316 614
rect 468004 610 468340 626
rect 467472 604 467524 610
rect 468004 604 468352 610
rect 468004 598 468300 604
rect 467472 546 467524 552
rect 468300 546 468352 552
rect 468496 598 468708 626
rect 467484 480 467512 546
rect 468496 542 468524 598
rect 468484 536 468536 542
rect 465704 468 466052 474
rect 465704 462 466000 468
rect 466000 410 466052 416
rect 466246 -960 466358 480
rect 467196 400 467248 406
rect 466900 348 467196 354
rect 466900 342 467248 348
rect 466900 326 467236 342
rect 467442 -960 467554 480
rect 468484 478 468536 484
rect 468680 480 468708 598
rect 469692 598 469904 626
rect 469220 536 469272 542
rect 469108 484 469220 490
rect 469692 490 469720 598
rect 468638 -960 468750 480
rect 469108 478 469272 484
rect 469108 462 469260 478
rect 469600 462 469720 490
rect 469876 480 469904 598
rect 470888 598 471100 626
rect 472808 672 472860 678
rect 472256 614 472308 620
rect 472512 620 472808 626
rect 474556 672 474608 678
rect 472512 614 472860 620
rect 469600 134 469628 462
rect 469588 128 469640 134
rect 469588 70 469640 76
rect 469834 -960 469946 480
rect 470888 338 470916 598
rect 471072 480 471100 598
rect 472268 480 472296 614
rect 472512 598 472848 614
rect 473280 598 473492 626
rect 484032 672 484084 678
rect 480810 640 480866 649
rect 474556 614 474608 620
rect 470876 332 470928 338
rect 470876 274 470928 280
rect 470600 128 470652 134
rect 470304 76 470600 82
rect 470304 70 470652 76
rect 470304 54 470640 70
rect 471030 -960 471142 480
rect 471408 338 471744 354
rect 471408 332 471756 338
rect 471408 326 471704 332
rect 471704 274 471756 280
rect 472226 -960 472338 480
rect 473280 66 473308 598
rect 473464 480 473492 598
rect 474568 480 474596 614
rect 475752 604 475804 610
rect 478216 598 478552 626
rect 479168 610 479320 626
rect 475752 546 475804 552
rect 476776 564 476988 592
rect 475108 536 475160 542
rect 474812 484 475108 490
rect 473268 60 473320 66
rect 473268 2 473320 8
rect 473422 -960 473534 480
rect 473708 66 474044 82
rect 473708 60 474056 66
rect 473708 54 474004 60
rect 474004 2 474056 8
rect 474526 -960 474638 480
rect 474812 478 475160 484
rect 475764 480 475792 546
rect 476212 536 476264 542
rect 475916 484 476212 490
rect 474812 462 475148 478
rect 475722 -960 475834 480
rect 475916 478 476264 484
rect 475916 462 476252 478
rect 476776 270 476804 564
rect 476960 480 476988 564
rect 477406 504 477462 513
rect 476764 264 476816 270
rect 476764 206 476816 212
rect 476918 -960 477030 480
rect 477112 462 477406 490
rect 477406 439 477462 448
rect 478114 218 478226 480
rect 477880 202 478226 218
rect 478524 202 478552 598
rect 479156 604 479320 610
rect 479208 598 479320 604
rect 480516 610 480668 626
rect 480516 604 480680 610
rect 480516 598 480628 604
rect 479156 546 479208 552
rect 480810 575 480812 584
rect 480628 546 480680 552
rect 480864 575 480866 584
rect 481730 640 481786 649
rect 483570 640 483626 649
rect 481730 575 481786 584
rect 482664 598 482816 626
rect 480812 546 480864 552
rect 481456 536 481508 542
rect 481508 484 481620 490
rect 479310 218 479422 480
rect 480506 354 480618 480
rect 481456 478 481620 484
rect 481744 480 481772 575
rect 481468 462 481620 478
rect 480720 400 480772 406
rect 480506 348 480720 354
rect 480506 342 480772 348
rect 480506 326 480760 342
rect 479524 264 479576 270
rect 479310 212 479524 218
rect 479310 206 479576 212
rect 477868 196 478226 202
rect 477920 190 478226 196
rect 477868 138 477920 144
rect 478114 -960 478226 190
rect 478512 196 478564 202
rect 478512 138 478564 144
rect 479310 190 479564 206
rect 479310 -960 479422 190
rect 480506 -960 480618 326
rect 481702 -960 481814 480
rect 482664 270 482692 598
rect 485136 672 485188 678
rect 484032 614 484084 620
rect 485024 620 485136 626
rect 487436 672 487488 678
rect 485024 614 485188 620
rect 487324 620 487436 626
rect 487712 672 487764 678
rect 487324 614 487488 620
rect 487632 620 487712 626
rect 492680 672 492732 678
rect 487632 614 487764 620
rect 488814 640 488870 649
rect 483570 575 483626 584
rect 482652 264 482704 270
rect 482652 206 482704 212
rect 482806 82 482918 480
rect 482974 128 483026 134
rect 482806 76 482974 82
rect 482806 70 483026 76
rect 482806 54 483014 70
rect 483584 66 483612 575
rect 483756 536 483808 542
rect 483808 484 483920 490
rect 483756 478 483920 484
rect 484044 480 484072 614
rect 485024 598 485176 614
rect 485228 604 485280 610
rect 485228 546 485280 552
rect 486424 604 486476 610
rect 487324 598 487476 614
rect 487632 598 487752 614
rect 486424 546 486476 552
rect 485240 480 485268 546
rect 486436 480 486464 546
rect 487632 480 487660 598
rect 492310 640 492366 649
rect 488814 575 488870 584
rect 489920 604 489972 610
rect 488828 480 488856 575
rect 489920 546 489972 552
rect 490944 598 491156 626
rect 489736 536 489788 542
rect 489624 484 489736 490
rect 483768 462 483920 478
rect 483572 60 483624 66
rect 482806 -960 482918 54
rect 483572 2 483624 8
rect 484002 -960 484114 480
rect 485198 -960 485310 480
rect 486056 264 486108 270
rect 486108 212 486220 218
rect 486056 206 486220 212
rect 486068 190 486220 206
rect 486394 -960 486506 480
rect 487590 -960 487702 480
rect 488428 66 488580 82
rect 488428 60 488592 66
rect 488428 54 488540 60
rect 488540 2 488592 8
rect 488786 -960 488898 480
rect 489624 478 489788 484
rect 489932 480 489960 546
rect 489624 462 489776 478
rect 489890 -960 490002 480
rect 490944 406 490972 598
rect 491128 480 491156 598
rect 492678 640 492680 649
rect 493324 672 493376 678
rect 492732 640 492734 649
rect 492310 575 492366 584
rect 492588 604 492640 610
rect 490932 400 490984 406
rect 490932 342 490984 348
rect 490932 264 490984 270
rect 490728 212 490932 218
rect 490728 206 490984 212
rect 490728 190 490972 206
rect 491086 -960 491198 480
rect 491832 474 492168 490
rect 492324 480 492352 575
rect 493028 620 493324 626
rect 494428 672 494480 678
rect 493028 614 493376 620
rect 494132 620 494428 626
rect 505192 672 505244 678
rect 494132 614 494480 620
rect 495898 640 495954 649
rect 493028 598 493364 614
rect 493508 604 493560 610
rect 492678 575 492734 584
rect 492588 546 492640 552
rect 494132 598 494468 614
rect 494704 604 494756 610
rect 493508 546 493560 552
rect 498106 640 498162 649
rect 495898 575 495954 584
rect 497094 606 497150 615
rect 494704 546 494756 552
rect 492600 490 492628 546
rect 492678 504 492734 513
rect 491832 468 492180 474
rect 491832 462 492128 468
rect 492128 410 492180 416
rect 492282 -960 492394 480
rect 492600 462 492678 490
rect 493520 480 493548 546
rect 494716 480 494744 546
rect 495912 480 495940 575
rect 500590 640 500646 649
rect 498640 610 498976 626
rect 499836 610 500172 626
rect 498106 575 498108 584
rect 497094 541 497150 550
rect 498160 575 498162 584
rect 498200 604 498252 610
rect 498108 546 498160 552
rect 498640 604 498988 610
rect 498640 598 498936 604
rect 498200 546 498252 552
rect 498936 546 498988 552
rect 499396 604 499448 610
rect 499836 604 500184 610
rect 499836 598 500132 604
rect 499396 546 499448 552
rect 500590 575 500646 584
rect 501616 598 501828 626
rect 503240 610 503576 626
rect 505744 672 505796 678
rect 505192 614 505244 620
rect 505448 620 505744 626
rect 507860 672 507912 678
rect 505448 614 505796 620
rect 507748 620 507860 626
rect 517152 672 517204 678
rect 509882 640 509938 649
rect 507748 614 507912 620
rect 500132 546 500184 552
rect 497108 480 497136 541
rect 497832 536 497884 542
rect 497536 484 497832 490
rect 492678 439 492734 448
rect 493478 -960 493590 480
rect 494674 -960 494786 480
rect 495348 400 495400 406
rect 495236 348 495348 354
rect 495236 342 495400 348
rect 495236 326 495388 342
rect 495870 -960 495982 480
rect 496432 202 496768 218
rect 496432 196 496780 202
rect 496432 190 496728 196
rect 496728 138 496780 144
rect 497066 -960 497178 480
rect 497536 478 497884 484
rect 498212 480 498240 546
rect 499408 480 499436 546
rect 500604 480 500632 575
rect 497536 462 497872 478
rect 498170 -960 498282 480
rect 499366 -960 499478 480
rect 500562 -960 500674 480
rect 500940 474 501276 490
rect 500940 468 501288 474
rect 500940 462 501236 468
rect 501236 410 501288 416
rect 501616 338 501644 598
rect 501800 480 501828 598
rect 502984 604 503036 610
rect 503240 604 503588 610
rect 503240 598 503536 604
rect 502984 546 503036 552
rect 503536 546 503588 552
rect 504008 564 504220 592
rect 502996 480 503024 546
rect 501604 332 501656 338
rect 501604 274 501656 280
rect 501758 -960 501870 480
rect 502340 128 502392 134
rect 502044 76 502340 82
rect 502044 70 502392 76
rect 502044 54 502380 70
rect 502954 -960 503066 480
rect 504008 66 504036 564
rect 504192 480 504220 564
rect 504640 536 504692 542
rect 504344 484 504640 490
rect 503996 60 504048 66
rect 503996 2 504048 8
rect 504150 -960 504262 480
rect 504344 478 504692 484
rect 504344 462 504680 478
rect 505204 218 505232 614
rect 505448 598 505784 614
rect 507748 598 507900 614
rect 508944 598 509280 626
rect 506308 564 506520 592
rect 506308 490 506336 564
rect 505346 218 505458 480
rect 506216 462 506336 490
rect 506492 480 506520 564
rect 509252 542 509280 598
rect 512458 640 512514 649
rect 510048 598 510384 626
rect 509882 575 509938 584
rect 507308 536 507360 542
rect 506216 270 506244 462
rect 505204 190 505458 218
rect 506204 264 506256 270
rect 506204 206 506256 212
rect 505346 -960 505458 190
rect 506450 -960 506562 480
rect 507308 478 507360 484
rect 509240 536 509292 542
rect 507320 354 507348 478
rect 507646 354 507758 480
rect 506644 338 506980 354
rect 506644 332 506992 338
rect 506644 326 506940 332
rect 507320 326 507758 354
rect 506940 274 506992 280
rect 507646 -960 507758 326
rect 508596 264 508648 270
rect 508842 218 508954 480
rect 509240 478 509292 484
rect 508648 212 508954 218
rect 508596 206 508954 212
rect 508608 190 508954 206
rect 509896 202 509924 575
rect 510038 218 510150 480
rect 510356 474 510384 598
rect 511276 598 511580 626
rect 511000 474 511152 490
rect 511276 480 511304 598
rect 510344 468 510396 474
rect 510344 410 510396 416
rect 510988 468 511152 474
rect 511040 462 511152 468
rect 510988 410 511040 416
rect 510252 264 510304 270
rect 510038 212 510252 218
rect 510038 206 510304 212
rect 508842 -960 508954 190
rect 509884 196 509936 202
rect 509884 138 509936 144
rect 510038 190 510292 206
rect 510038 -960 510150 190
rect 511234 -960 511346 480
rect 511552 406 511580 598
rect 514666 640 514722 649
rect 512458 575 512514 584
rect 513576 598 513788 626
rect 514556 598 514666 626
rect 512184 536 512236 542
rect 512236 484 512348 490
rect 512184 478 512348 484
rect 512472 480 512500 575
rect 513576 480 513604 598
rect 513760 542 513788 598
rect 515402 640 515458 649
rect 514666 575 514722 584
rect 514772 598 514984 626
rect 513748 536 513800 542
rect 512196 462 512348 478
rect 511540 400 511592 406
rect 511540 342 511592 348
rect 512430 -960 512542 480
rect 513288 400 513340 406
rect 513340 348 513452 354
rect 513288 342 513452 348
rect 513300 326 513452 342
rect 513534 -960 513646 480
rect 513748 478 513800 484
rect 514772 480 514800 598
rect 514730 -960 514842 480
rect 514956 406 514984 598
rect 515402 575 515458 584
rect 515954 640 516010 649
rect 517152 614 517204 620
rect 518992 672 519044 678
rect 520740 672 520792 678
rect 519044 620 519156 626
rect 518992 614 519156 620
rect 515954 575 516010 584
rect 515416 406 515444 575
rect 515968 480 515996 575
rect 517164 480 517192 614
rect 519004 598 519156 614
rect 519280 610 519584 626
rect 520740 614 520792 620
rect 521844 672 521896 678
rect 521844 614 521896 620
rect 523040 672 523092 678
rect 523316 672 523368 678
rect 523040 614 523092 620
rect 523222 640 523278 649
rect 519268 604 519584 610
rect 518176 564 518388 592
rect 514944 400 514996 406
rect 514944 342 514996 348
rect 515404 400 515456 406
rect 515404 342 515456 348
rect 515600 66 515752 82
rect 515588 60 515752 66
rect 515640 54 515752 60
rect 515588 2 515640 8
rect 515926 -960 516038 480
rect 516856 338 517008 354
rect 516856 332 517020 338
rect 516856 326 516968 332
rect 516968 274 517020 280
rect 517122 -960 517234 480
rect 518176 218 518204 564
rect 518360 480 518388 564
rect 519320 598 519584 604
rect 519268 546 519320 552
rect 519556 480 519584 598
rect 520752 480 520780 614
rect 521856 480 521884 614
rect 523052 480 523080 614
rect 523960 672 524012 678
rect 523316 614 523368 620
rect 523664 620 523960 626
rect 526260 672 526312 678
rect 523664 614 524012 620
rect 525430 640 525486 649
rect 523222 575 523278 584
rect 518084 202 518204 218
rect 518072 196 518204 202
rect 518124 190 518204 196
rect 518072 138 518124 144
rect 518164 128 518216 134
rect 517960 76 518164 82
rect 517960 70 518216 76
rect 517960 54 518204 70
rect 518318 -960 518430 480
rect 519514 -960 519626 480
rect 520260 202 520412 218
rect 520260 196 520424 202
rect 520260 190 520372 196
rect 520372 138 520424 144
rect 520710 -960 520822 480
rect 521568 264 521620 270
rect 521364 212 521568 218
rect 521364 206 521620 212
rect 521364 190 521608 206
rect 521814 -960 521926 480
rect 522856 400 522908 406
rect 522560 348 522856 354
rect 522560 342 522908 348
rect 522560 326 522896 342
rect 523010 -960 523122 480
rect 523236 474 523264 575
rect 523328 513 523356 614
rect 523664 598 524000 614
rect 524236 604 524288 610
rect 525964 620 526260 626
rect 533068 672 533120 678
rect 527178 640 527234 649
rect 525964 614 526312 620
rect 525964 598 526300 614
rect 526628 604 526680 610
rect 525430 575 525486 584
rect 524236 546 524288 552
rect 523314 504 523370 513
rect 523224 468 523276 474
rect 524248 480 524276 546
rect 525064 536 525116 542
rect 524768 484 525064 490
rect 523314 439 523370 448
rect 523224 410 523276 416
rect 524206 -960 524318 480
rect 524768 478 525116 484
rect 525444 480 525472 575
rect 527068 598 527178 626
rect 527178 575 527234 584
rect 527652 598 527864 626
rect 526628 546 526680 552
rect 526640 480 526668 546
rect 527652 513 527680 598
rect 527638 504 527694 513
rect 524768 462 525104 478
rect 525402 -960 525514 480
rect 526598 -960 526710 480
rect 527836 480 527864 598
rect 529020 604 529072 610
rect 529020 546 529072 552
rect 530124 604 530176 610
rect 530124 546 530176 552
rect 531148 598 531360 626
rect 531576 610 531912 626
rect 531576 604 531924 610
rect 531576 598 531872 604
rect 528466 504 528522 513
rect 527638 439 527694 448
rect 527794 -960 527906 480
rect 528172 462 528466 490
rect 529032 480 529060 546
rect 530136 480 530164 546
rect 528466 439 528522 448
rect 528990 -960 529102 480
rect 529664 128 529716 134
rect 529368 76 529664 82
rect 529368 70 529716 76
rect 529368 54 529704 70
rect 530094 -960 530206 480
rect 530766 368 530822 377
rect 530472 326 530766 354
rect 530766 303 530822 312
rect 531148 241 531176 598
rect 531332 480 531360 598
rect 531872 546 531924 552
rect 532344 598 532556 626
rect 532772 620 533068 626
rect 535828 672 535880 678
rect 534170 640 534226 649
rect 532772 614 533120 620
rect 532772 598 533108 614
rect 533448 598 533752 626
rect 533876 598 534170 626
rect 531134 232 531190 241
rect 531134 167 531190 176
rect 531290 -960 531402 480
rect 532344 66 532372 598
rect 532528 480 532556 598
rect 532332 60 532384 66
rect 532332 2 532384 8
rect 532486 -960 532598 480
rect 533448 474 533476 598
rect 533724 480 533752 598
rect 534980 598 535316 626
rect 540980 672 541032 678
rect 540518 640 540574 649
rect 535828 614 535880 620
rect 534170 575 534226 584
rect 534170 504 534226 513
rect 533436 468 533488 474
rect 533436 410 533488 416
rect 533682 -960 533794 480
rect 534170 439 534172 448
rect 534224 439 534226 448
rect 534172 410 534224 416
rect 534878 354 534990 480
rect 534552 338 534990 354
rect 534540 332 534990 338
rect 534592 326 534990 332
rect 534540 274 534592 280
rect 534878 -960 534990 326
rect 535288 134 535316 598
rect 535840 218 535868 614
rect 536176 598 536512 626
rect 537280 598 537616 626
rect 538476 598 538812 626
rect 536484 513 536512 598
rect 536470 504 536526 513
rect 536074 218 536186 480
rect 536470 439 536526 448
rect 537178 218 537290 480
rect 535840 190 536186 218
rect 536944 202 537290 218
rect 537588 202 537616 598
rect 538036 264 538088 270
rect 538374 218 538486 480
rect 538784 270 538812 598
rect 539428 598 539580 626
rect 539428 338 539456 598
rect 540574 598 540684 626
rect 553768 672 553820 678
rect 540980 614 541032 620
rect 540796 604 540848 610
rect 540518 575 540574 584
rect 540796 546 540848 552
rect 540808 480 540836 546
rect 540992 513 541020 614
rect 542004 598 542216 626
rect 540978 504 541034 513
rect 539570 354 539682 480
rect 539784 400 539836 406
rect 539570 348 539784 354
rect 539570 342 539836 348
rect 539416 332 539468 338
rect 539416 274 539468 280
rect 539570 326 539824 342
rect 538088 212 538486 218
rect 538036 206 538486 212
rect 538772 264 538824 270
rect 538772 206 538824 212
rect 535276 128 535328 134
rect 535276 70 535328 76
rect 536074 -960 536186 190
rect 536932 196 537290 202
rect 536984 190 537290 196
rect 536932 138 536984 144
rect 537178 -960 537290 190
rect 537576 196 537628 202
rect 538048 190 538486 206
rect 537576 138 537628 144
rect 538374 -960 538486 190
rect 539570 -960 539682 326
rect 540766 -960 540878 480
rect 542004 480 542032 598
rect 540978 439 541034 448
rect 541714 232 541770 241
rect 541770 190 541880 218
rect 541714 167 541770 176
rect 541962 -960 542074 480
rect 542188 406 542216 598
rect 543200 598 543412 626
rect 542634 504 542690 513
rect 542634 439 542690 448
rect 542818 504 542874 513
rect 542874 462 542984 490
rect 543200 480 543228 598
rect 543384 542 543412 598
rect 544212 598 544424 626
rect 543372 536 543424 542
rect 542818 439 542874 448
rect 542648 406 542676 439
rect 542176 400 542228 406
rect 542176 342 542228 348
rect 542636 400 542688 406
rect 542636 342 542688 348
rect 543158 -960 543270 480
rect 543372 478 543424 484
rect 543462 504 543518 513
rect 543462 439 543518 448
rect 543476 202 543504 439
rect 544212 406 544240 598
rect 544396 480 544424 598
rect 545500 598 545712 626
rect 545500 480 545528 598
rect 544200 400 544252 406
rect 544200 342 544252 348
rect 544088 202 544240 218
rect 543464 196 543516 202
rect 544088 196 544252 202
rect 544088 190 544200 196
rect 543464 138 543516 144
rect 544200 138 544252 144
rect 544354 -960 544466 480
rect 545120 400 545172 406
rect 545172 348 545284 354
rect 545120 342 545284 348
rect 545132 326 545284 342
rect 545458 -960 545570 480
rect 545684 474 545712 598
rect 546512 598 546724 626
rect 550896 610 551232 626
rect 546224 536 546276 542
rect 546276 484 546388 490
rect 546224 478 546388 484
rect 545672 468 545724 474
rect 546236 462 546388 478
rect 545672 410 545724 416
rect 546512 66 546540 598
rect 546696 480 546724 598
rect 549076 604 549128 610
rect 547892 564 548104 592
rect 546500 60 546552 66
rect 546500 2 546552 8
rect 546654 -960 546766 480
rect 547492 474 547736 490
rect 547892 480 547920 564
rect 547492 468 547748 474
rect 547492 462 547696 468
rect 547696 410 547748 416
rect 547850 -960 547962 480
rect 548076 377 548104 564
rect 549076 546 549128 552
rect 550272 604 550324 610
rect 550896 604 551244 610
rect 550896 598 551192 604
rect 550272 546 550324 552
rect 551192 546 551244 552
rect 551296 598 551508 626
rect 553044 610 553196 626
rect 555792 672 555844 678
rect 553768 614 553820 620
rect 548892 536 548944 542
rect 548688 484 548892 490
rect 548688 478 548944 484
rect 549088 480 549116 546
rect 550088 536 550140 542
rect 549792 484 550088 490
rect 548688 462 548932 478
rect 548062 368 548118 377
rect 548062 303 548118 312
rect 549046 -960 549158 480
rect 549792 478 550140 484
rect 550284 480 550312 546
rect 551296 490 551324 598
rect 549792 462 550128 478
rect 550242 -960 550354 480
rect 551204 462 551324 490
rect 551480 480 551508 598
rect 552664 604 552716 610
rect 552664 546 552716 552
rect 553032 604 553196 610
rect 553084 598 553196 604
rect 553032 546 553084 552
rect 552676 480 552704 546
rect 553780 480 553808 614
rect 554792 598 555004 626
rect 555496 620 555792 626
rect 556896 672 556948 678
rect 555496 614 555844 620
rect 556600 620 556896 626
rect 558736 672 558788 678
rect 558550 640 558606 649
rect 556600 614 556948 620
rect 555496 598 555832 614
rect 556600 598 556936 614
rect 557184 598 557396 626
rect 554792 513 554820 598
rect 554778 504 554834 513
rect 551204 377 551232 462
rect 551190 368 551246 377
rect 551190 303 551246 312
rect 551438 -960 551550 480
rect 552092 66 552428 82
rect 552092 60 552440 66
rect 552092 54 552388 60
rect 552388 2 552440 8
rect 552634 -960 552746 480
rect 553738 -960 553850 480
rect 554976 480 555004 598
rect 555988 564 556200 592
rect 555988 490 556016 564
rect 554778 439 554834 448
rect 554300 202 554636 218
rect 554300 196 554648 202
rect 554300 190 554596 196
rect 554596 138 554648 144
rect 554934 -960 555046 480
rect 555896 462 556016 490
rect 556172 480 556200 564
rect 555896 270 555924 462
rect 555884 264 555936 270
rect 555884 206 555936 212
rect 556130 -960 556242 480
rect 557184 338 557212 598
rect 557368 480 557396 598
rect 562600 672 562652 678
rect 560850 640 560906 649
rect 558788 620 558900 626
rect 558736 614 558900 620
rect 558748 598 558900 614
rect 559576 598 559788 626
rect 558550 575 558606 584
rect 558564 480 558592 575
rect 557172 332 557224 338
rect 557172 274 557224 280
rect 557326 -960 557438 480
rect 558000 264 558052 270
rect 557704 212 558000 218
rect 557704 206 558052 212
rect 557704 190 558040 206
rect 558522 -960 558634 480
rect 559576 241 559604 598
rect 559760 480 559788 598
rect 560850 575 560906 584
rect 561784 598 562088 626
rect 562304 620 562600 626
rect 562304 614 562652 620
rect 562304 598 562640 614
rect 563072 598 563284 626
rect 560864 480 560892 575
rect 559562 232 559618 241
rect 559562 167 559618 176
rect 559718 -960 559830 480
rect 560004 338 560248 354
rect 560004 332 560260 338
rect 560004 326 560208 332
rect 560208 274 560260 280
rect 560822 -960 560934 480
rect 561784 406 561812 598
rect 562060 480 562088 598
rect 561772 400 561824 406
rect 561772 342 561824 348
rect 561404 128 561456 134
rect 561108 76 561404 82
rect 561108 70 561456 76
rect 561108 54 561444 70
rect 562018 -960 562130 480
rect 563072 474 563100 598
rect 563256 480 563284 598
rect 563060 468 563112 474
rect 563060 410 563112 416
rect 563214 -960 563326 480
rect 563808 270 563836 2858
rect 564452 2106 564480 701082
rect 565082 699816 565138 699825
rect 565082 699751 565138 699760
rect 565096 73166 565124 699751
rect 565360 699100 565412 699106
rect 565360 699042 565412 699048
rect 565174 698728 565230 698737
rect 565174 698663 565230 698672
rect 565188 126954 565216 698663
rect 565268 698488 565320 698494
rect 565268 698430 565320 698436
rect 565280 245614 565308 698430
rect 565372 511970 565400 699042
rect 566646 698592 566702 698601
rect 566646 698527 566702 698536
rect 566556 698352 566608 698358
rect 566462 698320 566518 698329
rect 566556 698294 566608 698300
rect 566462 698255 566518 698264
rect 565360 511964 565412 511970
rect 565360 511906 565412 511912
rect 565268 245608 565320 245614
rect 565268 245550 565320 245556
rect 565176 126948 565228 126954
rect 565176 126890 565228 126896
rect 565084 73160 565136 73166
rect 565084 73102 565136 73108
rect 566476 33114 566504 698255
rect 566568 167006 566596 698294
rect 566556 167000 566608 167006
rect 566556 166942 566608 166948
rect 566660 113150 566688 698527
rect 566740 698420 566792 698426
rect 566740 698362 566792 698368
rect 566752 206990 566780 698362
rect 566740 206984 566792 206990
rect 566740 206926 566792 206932
rect 566648 113144 566700 113150
rect 566648 113086 566700 113092
rect 566464 33108 566516 33114
rect 566464 33050 566516 33056
rect 569236 20670 569264 702063
rect 569314 698864 569370 698873
rect 569314 698799 569370 698808
rect 569328 153202 569356 698799
rect 569420 233238 569448 702374
rect 572168 701752 572220 701758
rect 572168 701694 572220 701700
rect 571982 700088 572038 700097
rect 571982 700023 572038 700032
rect 570602 699952 570658 699961
rect 570602 699887 570658 699896
rect 569592 699236 569644 699242
rect 569592 699178 569644 699184
rect 569500 698692 569552 698698
rect 569500 698634 569552 698640
rect 569512 299470 569540 698634
rect 569604 592006 569632 699178
rect 569592 592000 569644 592006
rect 569592 591942 569644 591948
rect 569500 299464 569552 299470
rect 569500 299406 569552 299412
rect 569408 233232 569460 233238
rect 569408 233174 569460 233180
rect 569316 153196 569368 153202
rect 569316 153138 569368 153144
rect 570616 60722 570644 699887
rect 570880 699780 570932 699786
rect 570880 699722 570932 699728
rect 570788 698828 570840 698834
rect 570788 698770 570840 698776
rect 570696 698556 570748 698562
rect 570696 698498 570748 698504
rect 570708 273222 570736 698498
rect 570800 485790 570828 698770
rect 570892 632058 570920 699722
rect 570880 632052 570932 632058
rect 570880 631994 570932 632000
rect 570788 485784 570840 485790
rect 570788 485726 570840 485732
rect 570696 273216 570748 273222
rect 570696 273158 570748 273164
rect 571996 100706 572024 700023
rect 572074 697912 572130 697921
rect 572074 697847 572130 697856
rect 572088 353258 572116 697847
rect 572180 431934 572208 701694
rect 573456 701616 573508 701622
rect 573456 701558 573508 701564
rect 573362 700224 573418 700233
rect 573362 700159 573418 700168
rect 572260 699372 572312 699378
rect 572260 699314 572312 699320
rect 572272 644434 572300 699314
rect 572260 644428 572312 644434
rect 572260 644370 572312 644376
rect 572168 431928 572220 431934
rect 572168 431870 572220 431876
rect 572076 353252 572128 353258
rect 572076 353194 572128 353200
rect 573376 139398 573404 700159
rect 573468 379506 573496 701558
rect 573548 699032 573600 699038
rect 573548 698974 573600 698980
rect 573560 538218 573588 698974
rect 573652 564398 573680 702918
rect 574836 701480 574888 701486
rect 574836 701422 574888 701428
rect 574744 697672 574796 697678
rect 574744 697614 574796 697620
rect 573640 564392 573692 564398
rect 573640 564334 573692 564340
rect 573548 538212 573600 538218
rect 573548 538154 573600 538160
rect 573456 379500 573508 379506
rect 573456 379442 573508 379448
rect 573364 139392 573416 139398
rect 573364 139334 573416 139340
rect 571984 100700 572036 100706
rect 571984 100642 572036 100648
rect 574756 86970 574784 697614
rect 574848 313274 574876 701422
rect 574928 698624 574980 698630
rect 574928 698566 574980 698572
rect 574940 325650 574968 698566
rect 575032 618254 575060 703054
rect 576124 702500 576176 702506
rect 576124 702442 576176 702448
rect 575020 618248 575072 618254
rect 575020 618190 575072 618196
rect 574928 325644 574980 325650
rect 574928 325586 574980 325592
rect 574836 313268 574888 313274
rect 574836 313210 574888 313216
rect 574744 86964 574796 86970
rect 574744 86906 574796 86912
rect 570604 60716 570656 60722
rect 570604 60658 570656 60664
rect 576136 46918 576164 702442
rect 576308 698896 576360 698902
rect 576308 698838 576360 698844
rect 576216 698760 576268 698766
rect 576216 698702 576268 698708
rect 576228 419490 576256 698702
rect 576320 471986 576348 698838
rect 576412 672042 576440 703190
rect 578976 702840 579028 702846
rect 578976 702782 579028 702788
rect 577596 701956 577648 701962
rect 577596 701898 577648 701904
rect 577504 701276 577556 701282
rect 577504 701218 577556 701224
rect 576400 672036 576452 672042
rect 576400 671978 576452 671984
rect 576308 471980 576360 471986
rect 576308 471922 576360 471928
rect 576216 419484 576268 419490
rect 576216 419426 576268 419432
rect 577516 259418 577544 701218
rect 577608 578202 577636 701898
rect 578884 701684 578936 701690
rect 578884 701626 578936 701632
rect 577688 699916 577740 699922
rect 577688 699858 577740 699864
rect 577700 684486 577728 699858
rect 577688 684480 577740 684486
rect 577688 684422 577740 684428
rect 577596 578196 577648 578202
rect 577596 578138 577648 578144
rect 578896 365129 578924 701626
rect 578988 404977 579016 702782
rect 580540 700800 580592 700806
rect 580540 700742 580592 700748
rect 580448 700664 580500 700670
rect 580448 700606 580500 700612
rect 580080 700596 580132 700602
rect 580080 700538 580132 700544
rect 580092 697241 580120 700538
rect 580356 699576 580408 699582
rect 580356 699518 580408 699524
rect 580262 699136 580318 699145
rect 580262 699071 580318 699080
rect 580078 697232 580134 697241
rect 580078 697167 580134 697176
rect 579620 672036 579672 672042
rect 579620 671978 579672 671984
rect 579632 670721 579660 671978
rect 579618 670712 579674 670721
rect 579618 670647 579674 670656
rect 580172 644428 580224 644434
rect 580172 644370 580224 644376
rect 580184 644065 580212 644370
rect 580170 644056 580226 644065
rect 580170 643991 580226 644000
rect 580172 632052 580224 632058
rect 580172 631994 580224 632000
rect 580184 630873 580212 631994
rect 580170 630864 580226 630873
rect 580170 630799 580226 630808
rect 580172 618248 580224 618254
rect 580172 618190 580224 618196
rect 580184 617545 580212 618190
rect 580170 617536 580226 617545
rect 580170 617471 580226 617480
rect 580172 592000 580224 592006
rect 580172 591942 580224 591948
rect 580184 591025 580212 591942
rect 580170 591016 580226 591025
rect 580170 590951 580226 590960
rect 580172 564392 580224 564398
rect 580170 564360 580172 564369
rect 580224 564360 580226 564369
rect 580170 564295 580226 564304
rect 580172 538212 580224 538218
rect 580172 538154 580224 538160
rect 580184 537849 580212 538154
rect 580170 537840 580226 537849
rect 580170 537775 580226 537784
rect 580172 511964 580224 511970
rect 580172 511906 580224 511912
rect 580184 511329 580212 511906
rect 580170 511320 580226 511329
rect 580170 511255 580226 511264
rect 579620 485784 579672 485790
rect 579620 485726 579672 485732
rect 579632 484673 579660 485726
rect 579618 484664 579674 484673
rect 579618 484599 579674 484608
rect 579804 471980 579856 471986
rect 579804 471922 579856 471928
rect 579816 471481 579844 471922
rect 579802 471472 579858 471481
rect 579802 471407 579858 471416
rect 579712 431928 579764 431934
rect 579712 431870 579764 431876
rect 579724 431633 579752 431870
rect 579710 431624 579766 431633
rect 579710 431559 579766 431568
rect 580172 419484 580224 419490
rect 580172 419426 580224 419432
rect 580184 418305 580212 419426
rect 580170 418296 580226 418305
rect 580170 418231 580226 418240
rect 578974 404968 579030 404977
rect 578974 404903 579030 404912
rect 579620 379500 579672 379506
rect 579620 379442 579672 379448
rect 579632 378457 579660 379442
rect 579618 378448 579674 378457
rect 579618 378383 579674 378392
rect 578882 365120 578938 365129
rect 578882 365055 578938 365064
rect 580172 353252 580224 353258
rect 580172 353194 580224 353200
rect 580184 351937 580212 353194
rect 580170 351928 580226 351937
rect 580170 351863 580226 351872
rect 580172 325644 580224 325650
rect 580172 325586 580224 325592
rect 580184 325281 580212 325586
rect 580170 325272 580226 325281
rect 580170 325207 580226 325216
rect 580172 313268 580224 313274
rect 580172 313210 580224 313216
rect 580184 312089 580212 313210
rect 580170 312080 580226 312089
rect 580170 312015 580226 312024
rect 580172 299464 580224 299470
rect 580172 299406 580224 299412
rect 580184 298761 580212 299406
rect 580170 298752 580226 298761
rect 580170 298687 580226 298696
rect 579620 273216 579672 273222
rect 579620 273158 579672 273164
rect 579632 272241 579660 273158
rect 579618 272232 579674 272241
rect 579618 272167 579674 272176
rect 577504 259412 577556 259418
rect 577504 259354 577556 259360
rect 580172 245608 580224 245614
rect 580170 245576 580172 245585
rect 580224 245576 580226 245585
rect 580170 245511 580226 245520
rect 579988 233232 580040 233238
rect 579988 233174 580040 233180
rect 580000 232393 580028 233174
rect 579986 232384 580042 232393
rect 579986 232319 580042 232328
rect 580172 206984 580224 206990
rect 580172 206926 580224 206932
rect 580184 205737 580212 206926
rect 580170 205728 580226 205737
rect 580170 205663 580226 205672
rect 580172 167000 580224 167006
rect 580172 166942 580224 166948
rect 580184 165889 580212 166942
rect 580170 165880 580226 165889
rect 580170 165815 580226 165824
rect 579804 153196 579856 153202
rect 579804 153138 579856 153144
rect 579816 152697 579844 153138
rect 579802 152688 579858 152697
rect 579802 152623 579858 152632
rect 580172 139392 580224 139398
rect 580170 139360 580172 139369
rect 580224 139360 580226 139369
rect 580170 139295 580226 139304
rect 580172 126948 580224 126954
rect 580172 126890 580224 126896
rect 580184 126041 580212 126890
rect 580170 126032 580226 126041
rect 580170 125967 580226 125976
rect 580172 113144 580224 113150
rect 580172 113086 580224 113092
rect 580184 112849 580212 113086
rect 580170 112840 580226 112849
rect 580170 112775 580226 112784
rect 580172 100700 580224 100706
rect 580172 100642 580224 100648
rect 580184 99521 580212 100642
rect 580170 99512 580226 99521
rect 580170 99447 580226 99456
rect 580172 86964 580224 86970
rect 580172 86906 580224 86912
rect 580184 86193 580212 86906
rect 580170 86184 580226 86193
rect 580170 86119 580226 86128
rect 579988 73160 580040 73166
rect 579988 73102 580040 73108
rect 580000 73001 580028 73102
rect 579986 72992 580042 73001
rect 579986 72927 580042 72936
rect 580172 60716 580224 60722
rect 580172 60658 580224 60664
rect 580184 59673 580212 60658
rect 580170 59664 580226 59673
rect 580170 59599 580226 59608
rect 576124 46912 576176 46918
rect 576124 46854 576176 46860
rect 580172 46912 580224 46918
rect 580172 46854 580224 46860
rect 580184 46345 580212 46854
rect 580170 46336 580226 46345
rect 580170 46271 580226 46280
rect 580170 33144 580226 33153
rect 580170 33079 580172 33088
rect 580224 33079 580226 33088
rect 580172 33050 580224 33056
rect 569224 20664 569276 20670
rect 569224 20606 569276 20612
rect 580172 20664 580224 20670
rect 580172 20606 580224 20612
rect 580184 19825 580212 20606
rect 580170 19816 580226 19825
rect 580170 19751 580226 19760
rect 580276 6633 580304 699071
rect 580368 179217 580396 699518
rect 580460 192545 580488 700606
rect 580552 219065 580580 700742
rect 580724 700732 580776 700738
rect 580724 700674 580776 700680
rect 580632 700528 580684 700534
rect 580632 700470 580684 700476
rect 580644 458153 580672 700470
rect 580736 524521 580764 700674
rect 580816 684480 580868 684486
rect 580816 684422 580868 684428
rect 580828 683913 580856 684422
rect 580814 683904 580870 683913
rect 580814 683839 580870 683848
rect 580816 578196 580868 578202
rect 580816 578138 580868 578144
rect 580828 577697 580856 578138
rect 580814 577688 580870 577697
rect 580814 577623 580870 577632
rect 580722 524512 580778 524521
rect 580722 524447 580778 524456
rect 580630 458144 580686 458153
rect 580630 458079 580686 458088
rect 580632 259412 580684 259418
rect 580632 259354 580684 259360
rect 580644 258913 580672 259354
rect 580630 258904 580686 258913
rect 580630 258839 580686 258848
rect 580538 219056 580594 219065
rect 580538 218991 580594 219000
rect 580446 192536 580502 192545
rect 580446 192471 580502 192480
rect 580354 179208 580410 179217
rect 580354 179143 580410 179152
rect 580262 6624 580318 6633
rect 580262 6559 580318 6568
rect 569132 3120 569184 3126
rect 569132 3062 569184 3068
rect 577412 3120 577464 3126
rect 577412 3062 577464 3068
rect 564440 2100 564492 2106
rect 564440 2042 564492 2048
rect 565820 1420 565872 1426
rect 565820 1362 565872 1368
rect 569040 1420 569092 1426
rect 569040 1362 569092 1368
rect 564440 1284 564492 1290
rect 564440 1226 564492 1232
rect 564452 480 564480 1226
rect 565832 882 565860 1362
rect 565820 876 565872 882
rect 565820 818 565872 824
rect 566832 808 566884 814
rect 566832 750 566884 756
rect 569052 762 569080 1362
rect 569144 1018 569172 3062
rect 573916 2984 573968 2990
rect 573916 2926 573968 2932
rect 571524 1216 571576 1222
rect 571524 1158 571576 1164
rect 569132 1012 569184 1018
rect 569132 954 569184 960
rect 570328 808 570380 814
rect 565464 598 565676 626
rect 565464 542 565492 598
rect 565452 536 565504 542
rect 563796 264 563848 270
rect 563796 206 563848 212
rect 564410 -960 564522 480
rect 565452 478 565504 484
rect 565648 480 565676 598
rect 566844 480 566872 750
rect 569052 734 569172 762
rect 570328 750 570380 756
rect 568028 604 568080 610
rect 568028 546 568080 552
rect 568040 480 568068 546
rect 569144 480 569172 734
rect 570340 480 570368 750
rect 571536 480 571564 1158
rect 572732 598 572944 626
rect 572732 480 572760 598
rect 565606 -960 565718 480
rect 566802 -960 566914 480
rect 567998 -960 568110 480
rect 569102 -960 569214 480
rect 570298 -960 570410 480
rect 571494 -960 571606 480
rect 572690 -960 572802 480
rect 572916 202 572944 598
rect 573928 480 573956 2926
rect 575480 2916 575532 2922
rect 575480 2858 575532 2864
rect 575112 740 575164 746
rect 575112 682 575164 688
rect 575124 480 575152 682
rect 575492 678 575520 2858
rect 576308 2848 576360 2854
rect 576308 2790 576360 2796
rect 575480 672 575532 678
rect 575480 614 575532 620
rect 576320 480 576348 2790
rect 577424 480 577452 3062
rect 583392 3052 583444 3058
rect 583392 2994 583444 3000
rect 582196 2916 582248 2922
rect 582196 2858 582248 2864
rect 578436 598 578648 626
rect 578436 490 578464 598
rect 572904 196 572956 202
rect 572904 138 572956 144
rect 573886 -960 573998 480
rect 575082 -960 575194 480
rect 576278 -960 576390 480
rect 577382 -960 577494 480
rect 578344 462 578464 490
rect 578620 480 578648 598
rect 580828 598 581040 626
rect 578344 338 578372 462
rect 578332 332 578384 338
rect 578332 274 578384 280
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580828 354 580856 598
rect 581012 480 581040 598
rect 582208 480 582236 2858
rect 583404 480 583432 2994
rect 580736 326 580856 354
rect 580736 134 580764 326
rect 580724 128 580776 134
rect 580724 70 580776 76
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 294 701392 350 701448
rect 386 697584 442 697640
rect 1490 684256 1546 684312
rect 1582 632032 1638 632088
rect 938 606056 994 606112
rect 1674 579944 1730 580000
rect 846 553832 902 553888
rect 1858 698128 1914 698184
rect 1766 527856 1822 527912
rect 754 501744 810 501800
rect 1858 475632 1914 475688
rect 2134 701256 2190 701312
rect 1950 449520 2006 449576
rect 662 358400 718 358456
rect 570 345344 626 345400
rect 570 241032 626 241088
rect 570 214920 626 214976
rect 570 201864 626 201920
rect 202 163376 258 163432
rect 110 111152 166 111208
rect 18 71848 74 71904
rect 2318 701528 2374 701584
rect 2226 267144 2282 267200
rect 2502 697720 2558 697776
rect 4066 700576 4122 700632
rect 3146 700440 3202 700496
rect 2686 697992 2742 698048
rect 3054 697856 3110 697912
rect 2962 671200 3018 671256
rect 3054 566888 3110 566944
rect 2778 514836 2780 514856
rect 2780 514836 2832 514856
rect 2832 514836 2834 514856
rect 2778 514800 2834 514836
rect 3146 462576 3202 462632
rect 2686 423544 2742 423600
rect 3238 410488 3294 410544
rect 3514 698400 3570 698456
rect 3330 397432 3386 397488
rect 2594 371320 2650 371376
rect 2502 319232 2558 319288
rect 2410 306176 2466 306232
rect 2318 188808 2374 188864
rect 2134 97552 2190 97608
rect 2042 32408 2098 32464
rect 3882 700304 3938 700360
rect 3790 698944 3846 699000
rect 4250 658144 4306 658200
rect 4066 619112 4122 619168
rect 3974 293120 4030 293176
rect 6642 701664 6698 701720
rect 16302 702072 16358 702128
rect 70122 701936 70178 701992
rect 60416 700168 60472 700224
rect 46018 700032 46074 700088
rect 31206 699896 31262 699952
rect 26146 699760 26202 699816
rect 266358 701800 266414 701856
rect 260838 701664 260894 701720
rect 286690 701120 286746 701176
rect 295338 701120 295394 701176
rect 326066 701936 326122 701992
rect 326250 701936 326306 701992
rect 384302 700576 384358 700632
rect 399022 701936 399078 701992
rect 428462 700440 428518 700496
rect 497278 701528 497334 701584
rect 502338 701392 502394 701448
rect 526718 701800 526774 701856
rect 516966 700304 517022 700360
rect 531686 701256 531742 701312
rect 546498 701664 546554 701720
rect 569222 702072 569278 702128
rect 561126 701936 561182 701992
rect 453946 699508 454002 699544
rect 453946 699488 453948 699508
rect 453948 699488 454000 699508
rect 454000 699488 454002 699508
rect 11610 699352 11666 699408
rect 41050 699352 41106 699408
rect 50894 699352 50950 699408
rect 55770 699352 55826 699408
rect 124586 699352 124642 699408
rect 326250 699352 326306 699408
rect 418710 699352 418766 699408
rect 433430 699352 433486 699408
rect 462870 699352 462926 699408
rect 492586 699352 492642 699408
rect 511998 699352 512054 699408
rect 541530 699352 541586 699408
rect 4066 254088 4122 254144
rect 3882 149776 3938 149832
rect 3790 136720 3846 136776
rect 3698 84632 3754 84688
rect 3606 58520 3662 58576
rect 3514 45464 3570 45520
rect 3422 19352 3478 19408
rect 2962 6432 3018 6488
rect 4066 584 4122 640
rect 7838 584 7894 640
rect 9954 584 10010 640
rect 13726 584 13782 640
rect 26514 584 26570 640
rect 28722 604 28778 640
rect 28722 584 28724 604
rect 28724 584 28776 604
rect 28776 584 28778 604
rect 27894 448 27950 504
rect 30286 584 30342 640
rect 31298 584 31354 640
rect 33598 584 33654 640
rect 32218 312 32274 368
rect 33874 448 33930 504
rect 35990 584 36046 640
rect 34978 312 35034 368
rect 36174 448 36230 504
rect 38474 584 38530 640
rect 52550 584 52606 640
rect 53562 448 53618 504
rect 54206 584 54262 640
rect 56046 584 56102 640
rect 55310 448 55366 504
rect 57610 584 57666 640
rect 58438 584 58494 640
rect 57426 448 57482 504
rect 59818 584 59874 640
rect 60830 584 60886 640
rect 58806 448 58862 504
rect 59450 448 59506 504
rect 62118 584 62174 640
rect 61106 448 61162 504
rect 142066 584 142122 640
rect 143446 584 143502 640
rect 144734 584 144790 640
rect 145746 584 145802 640
rect 143722 448 143778 504
rect 147126 584 147182 640
rect 148966 584 149022 640
rect 147770 448 147826 504
rect 149334 448 149390 504
rect 150622 584 150678 640
rect 151818 584 151874 640
rect 150254 448 150310 504
rect 164790 584 164846 640
rect 167366 584 167422 640
rect 169482 584 169538 640
rect 168194 312 168250 368
rect 171966 584 172022 640
rect 172978 584 173034 640
rect 170954 312 171010 368
rect 171690 312 171746 368
rect 173898 448 173954 504
rect 175462 584 175518 640
rect 176382 584 176438 640
rect 173990 312 174046 368
rect 175186 312 175242 368
rect 176842 448 176898 504
rect 177486 448 177542 504
rect 179050 584 179106 640
rect 180246 584 180302 640
rect 177670 312 177726 368
rect 178682 312 178738 368
rect 182086 584 182142 640
rect 184938 584 184994 640
rect 181258 312 181314 368
rect 186594 448 186650 504
rect 192298 584 192354 640
rect 188802 312 188858 368
rect 189906 448 189962 504
rect 192206 312 192262 368
rect 194046 448 194102 504
rect 195610 584 195666 640
rect 197910 584 197966 640
rect 200026 584 200082 640
rect 196622 312 196678 368
rect 197726 40 197782 96
rect 198922 448 198978 504
rect 200118 312 200174 368
rect 201314 448 201370 504
rect 203890 584 203946 640
rect 204166 604 204222 640
rect 204166 584 204168 604
rect 204168 584 204220 604
rect 204220 584 204222 604
rect 202510 312 202566 368
rect 202418 176 202474 232
rect 201682 40 201738 96
rect 204902 448 204958 504
rect 207386 584 207442 640
rect 208214 584 208270 640
rect 208398 584 208454 640
rect 204810 312 204866 368
rect 206006 448 206062 504
rect 206926 448 206982 504
rect 209318 584 209374 640
rect 208766 312 208822 368
rect 210790 448 210846 504
rect 213366 584 213422 640
rect 216126 584 216182 640
rect 220450 584 220506 640
rect 223854 584 223910 640
rect 228730 584 228786 640
rect 230938 584 230994 640
rect 235814 584 235870 640
rect 238850 584 238906 640
rect 242254 448 242310 504
rect 244094 584 244150 640
rect 249062 584 249118 640
rect 247314 448 247370 504
rect 250902 448 250958 504
rect 254674 584 254730 640
rect 255226 584 255282 640
rect 255870 584 255926 640
rect 257066 584 257122 640
rect 267278 584 267334 640
rect 269486 448 269542 504
rect 273626 584 273682 640
rect 275190 584 275246 640
rect 278594 584 278650 640
rect 276202 448 276258 504
rect 282090 448 282146 504
rect 285402 584 285458 640
rect 285678 584 285734 640
rect 285218 448 285274 504
rect 287794 584 287850 640
rect 286414 312 286470 368
rect 292578 584 292634 640
rect 293406 312 293462 368
rect 293866 584 293922 640
rect 294878 584 294934 640
rect 295614 584 295670 640
rect 303158 584 303214 640
rect 303802 448 303858 504
rect 305826 584 305882 640
rect 306930 448 306986 504
rect 313830 584 313886 640
rect 309966 448 310022 504
rect 318522 584 318578 640
rect 318890 584 318946 640
rect 319718 584 319774 640
rect 328458 176 328514 232
rect 334898 584 334954 640
rect 336646 176 336702 232
rect 338302 448 338358 504
rect 344558 584 344614 640
rect 344742 584 344798 640
rect 345754 584 345810 640
rect 347870 448 347926 504
rect 350170 584 350226 640
rect 348422 468 348478 504
rect 348422 448 348424 468
rect 348424 448 348476 468
rect 348476 448 348478 468
rect 350262 448 350318 504
rect 349434 176 349490 232
rect 352562 584 352618 640
rect 351458 176 351514 232
rect 354034 584 354090 640
rect 359922 584 359978 640
rect 363786 620 363788 640
rect 363788 620 363840 640
rect 363840 620 363842 640
rect 363786 584 363842 620
rect 363694 448 363750 504
rect 370594 584 370650 640
rect 374090 584 374146 640
rect 374274 584 374330 640
rect 375286 584 375342 640
rect 375470 584 375526 640
rect 364982 332 365038 368
rect 364982 312 364984 332
rect 364984 312 365036 332
rect 365036 312 365038 332
rect 373078 312 373134 368
rect 374366 484 374368 504
rect 374368 484 374420 504
rect 374420 484 374422 504
rect 374366 448 374422 484
rect 378874 584 378930 640
rect 379058 584 379114 640
rect 377494 448 377550 504
rect 376758 60 376814 96
rect 376758 40 376760 60
rect 376760 40 376812 60
rect 376812 40 376814 60
rect 381174 584 381230 640
rect 379610 468 379666 504
rect 379610 448 379612 468
rect 379612 448 379664 468
rect 379664 448 379666 468
rect 379794 40 379850 96
rect 383566 584 383622 640
rect 382002 176 382058 232
rect 384210 448 384266 504
rect 384578 176 384634 232
rect 391018 584 391074 640
rect 395526 448 395582 504
rect 402518 584 402574 640
rect 403070 620 403072 640
rect 403072 620 403124 640
rect 403124 620 403126 640
rect 403070 584 403126 620
rect 403622 584 403678 640
rect 405646 584 405702 640
rect 408406 584 408462 640
rect 407486 484 407488 504
rect 407488 484 407540 504
rect 407540 484 407542 504
rect 407486 448 407542 484
rect 409602 584 409658 640
rect 421010 620 421012 640
rect 421012 620 421064 640
rect 421064 620 421066 640
rect 418618 448 418674 504
rect 421010 584 421066 620
rect 423770 584 423826 640
rect 424966 584 425022 640
rect 427910 620 427912 640
rect 427912 620 427964 640
rect 427964 620 427966 640
rect 427910 584 427966 620
rect 429658 584 429714 640
rect 431038 584 431094 640
rect 432050 584 432106 640
rect 453486 448 453542 504
rect 456062 584 456118 640
rect 460386 584 460442 640
rect 460938 584 460994 640
rect 462778 584 462834 640
rect 463974 584 464030 640
rect 461766 448 461822 504
rect 461950 448 462006 504
rect 477406 448 477462 504
rect 480810 604 480866 640
rect 480810 584 480812 604
rect 480812 584 480864 604
rect 480864 584 480866 604
rect 481730 584 481786 640
rect 483570 584 483626 640
rect 488814 584 488870 640
rect 492310 584 492366 640
rect 492678 620 492680 640
rect 492680 620 492732 640
rect 492732 620 492734 640
rect 492678 584 492734 620
rect 495898 584 495954 640
rect 492678 448 492734 504
rect 497094 550 497150 606
rect 498106 604 498162 640
rect 498106 584 498108 604
rect 498108 584 498160 604
rect 498160 584 498162 604
rect 500590 584 500646 640
rect 509882 584 509938 640
rect 512458 584 512514 640
rect 514666 584 514722 640
rect 515402 584 515458 640
rect 515954 584 516010 640
rect 523222 584 523278 640
rect 525430 584 525486 640
rect 523314 448 523370 504
rect 527178 584 527234 640
rect 527638 448 527694 504
rect 528466 448 528522 504
rect 530766 312 530822 368
rect 531134 176 531190 232
rect 534170 584 534226 640
rect 534170 468 534226 504
rect 534170 448 534172 468
rect 534172 448 534224 468
rect 534224 448 534226 468
rect 536470 448 536526 504
rect 540518 584 540574 640
rect 540978 448 541034 504
rect 541714 176 541770 232
rect 542634 448 542690 504
rect 542818 448 542874 504
rect 543462 448 543518 504
rect 548062 312 548118 368
rect 551190 312 551246 368
rect 554778 448 554834 504
rect 558550 584 558606 640
rect 560850 584 560906 640
rect 559562 176 559618 232
rect 565082 699760 565138 699816
rect 565174 698672 565230 698728
rect 566646 698536 566702 698592
rect 566462 698264 566518 698320
rect 569314 698808 569370 698864
rect 571982 700032 572038 700088
rect 570602 699896 570658 699952
rect 572074 697856 572130 697912
rect 573362 700168 573418 700224
rect 580262 699080 580318 699136
rect 580078 697176 580134 697232
rect 579618 670656 579674 670712
rect 580170 644000 580226 644056
rect 580170 630808 580226 630864
rect 580170 617480 580226 617536
rect 580170 590960 580226 591016
rect 580170 564340 580172 564360
rect 580172 564340 580224 564360
rect 580224 564340 580226 564360
rect 580170 564304 580226 564340
rect 580170 537784 580226 537840
rect 580170 511264 580226 511320
rect 579618 484608 579674 484664
rect 579802 471416 579858 471472
rect 579710 431568 579766 431624
rect 580170 418240 580226 418296
rect 578974 404912 579030 404968
rect 579618 378392 579674 378448
rect 578882 365064 578938 365120
rect 580170 351872 580226 351928
rect 580170 325216 580226 325272
rect 580170 312024 580226 312080
rect 580170 298696 580226 298752
rect 579618 272176 579674 272232
rect 580170 245556 580172 245576
rect 580172 245556 580224 245576
rect 580224 245556 580226 245576
rect 580170 245520 580226 245556
rect 579986 232328 580042 232384
rect 580170 205672 580226 205728
rect 580170 165824 580226 165880
rect 579802 152632 579858 152688
rect 580170 139340 580172 139360
rect 580172 139340 580224 139360
rect 580224 139340 580226 139360
rect 580170 139304 580226 139340
rect 580170 125976 580226 126032
rect 580170 112784 580226 112840
rect 580170 99456 580226 99512
rect 580170 86128 580226 86184
rect 579986 72936 580042 72992
rect 580170 59608 580226 59664
rect 580170 46280 580226 46336
rect 580170 33108 580226 33144
rect 580170 33088 580172 33108
rect 580172 33088 580224 33108
rect 580224 33088 580226 33108
rect 580170 19760 580226 19816
rect 580814 683848 580870 683904
rect 580814 577632 580870 577688
rect 580722 524456 580778 524512
rect 580630 458088 580686 458144
rect 580630 258848 580686 258904
rect 580538 219000 580594 219056
rect 580446 192480 580502 192536
rect 580354 179152 580410 179208
rect 580262 6568 580318 6624
<< metal3 >>
rect 16297 702130 16363 702133
rect 569217 702130 569283 702133
rect 16297 702128 569283 702130
rect 16297 702072 16302 702128
rect 16358 702072 569222 702128
rect 569278 702072 569283 702128
rect 16297 702070 569283 702072
rect 16297 702067 16363 702070
rect 569217 702067 569283 702070
rect 70117 701994 70183 701997
rect 326061 701994 326127 701997
rect 70117 701992 326127 701994
rect 70117 701936 70122 701992
rect 70178 701936 326066 701992
rect 326122 701936 326127 701992
rect 70117 701934 326127 701936
rect 70117 701931 70183 701934
rect 326061 701931 326127 701934
rect 326245 701994 326311 701997
rect 399017 701994 399083 701997
rect 326245 701992 399083 701994
rect 326245 701936 326250 701992
rect 326306 701936 399022 701992
rect 399078 701936 399083 701992
rect 326245 701934 399083 701936
rect 326245 701931 326311 701934
rect 399017 701931 399083 701934
rect 453982 701932 453988 701996
rect 454052 701994 454058 701996
rect 561121 701994 561187 701997
rect 454052 701992 561187 701994
rect 454052 701936 561126 701992
rect 561182 701936 561187 701992
rect 454052 701934 561187 701936
rect 454052 701932 454058 701934
rect 561121 701931 561187 701934
rect 266353 701858 266419 701861
rect 526713 701858 526779 701861
rect 266353 701856 526779 701858
rect 266353 701800 266358 701856
rect 266414 701800 526718 701856
rect 526774 701800 526779 701856
rect 266353 701798 526779 701800
rect 266353 701795 266419 701798
rect 526713 701795 526779 701798
rect 6637 701722 6703 701725
rect 259126 701722 259132 701724
rect 6637 701720 259132 701722
rect 6637 701664 6642 701720
rect 6698 701664 259132 701720
rect 6637 701662 259132 701664
rect 6637 701659 6703 701662
rect 259126 701660 259132 701662
rect 259196 701660 259202 701724
rect 260833 701722 260899 701725
rect 546493 701722 546559 701725
rect 260833 701720 546559 701722
rect 260833 701664 260838 701720
rect 260894 701664 546498 701720
rect 546554 701664 546559 701720
rect 260833 701662 546559 701664
rect 260833 701659 260899 701662
rect 546493 701659 546559 701662
rect 2313 701586 2379 701589
rect 497273 701586 497339 701589
rect 2313 701584 497339 701586
rect 2313 701528 2318 701584
rect 2374 701528 497278 701584
rect 497334 701528 497339 701584
rect 2313 701526 497339 701528
rect 2313 701523 2379 701526
rect 497273 701523 497339 701526
rect 289 701450 355 701453
rect 502333 701450 502399 701453
rect 289 701448 502399 701450
rect 289 701392 294 701448
rect 350 701392 502338 701448
rect 502394 701392 502399 701448
rect 289 701390 502399 701392
rect 289 701387 355 701390
rect 502333 701387 502399 701390
rect 2129 701314 2195 701317
rect 531681 701314 531747 701317
rect 2129 701312 531747 701314
rect 2129 701256 2134 701312
rect 2190 701256 531686 701312
rect 531742 701256 531747 701312
rect 2129 701254 531747 701256
rect 2129 701251 2195 701254
rect 531681 701251 531747 701254
rect 286685 701178 286751 701181
rect 295333 701178 295399 701181
rect 286685 701176 295399 701178
rect 286685 701120 286690 701176
rect 286746 701120 295338 701176
rect 295394 701120 295399 701176
rect 286685 701118 295399 701120
rect 286685 701115 286751 701118
rect 295333 701115 295399 701118
rect 4061 700634 4127 700637
rect 384297 700634 384363 700637
rect 4061 700632 384363 700634
rect 4061 700576 4066 700632
rect 4122 700576 384302 700632
rect 384358 700576 384363 700632
rect 4061 700574 384363 700576
rect 4061 700571 4127 700574
rect 384297 700571 384363 700574
rect 3141 700498 3207 700501
rect 428457 700498 428523 700501
rect 3141 700496 428523 700498
rect 3141 700440 3146 700496
rect 3202 700440 428462 700496
rect 428518 700440 428523 700496
rect 3141 700438 428523 700440
rect 3141 700435 3207 700438
rect 428457 700435 428523 700438
rect 3877 700362 3943 700365
rect 516961 700362 517027 700365
rect 3877 700360 517027 700362
rect 3877 700304 3882 700360
rect 3938 700304 516966 700360
rect 517022 700304 517027 700360
rect 3877 700302 517027 700304
rect 3877 700299 3943 700302
rect 516961 700299 517027 700302
rect 60411 700226 60477 700229
rect 573357 700226 573423 700229
rect 60411 700224 573423 700226
rect 60411 700168 60416 700224
rect 60472 700168 573362 700224
rect 573418 700168 573423 700224
rect 60411 700166 573423 700168
rect 60411 700163 60477 700166
rect 573357 700163 573423 700166
rect 46013 700090 46079 700093
rect 571977 700090 572043 700093
rect 46013 700088 572043 700090
rect 46013 700032 46018 700088
rect 46074 700032 571982 700088
rect 572038 700032 572043 700088
rect 46013 700030 572043 700032
rect 46013 700027 46079 700030
rect 571977 700027 572043 700030
rect 31201 699954 31267 699957
rect 570597 699954 570663 699957
rect 31201 699952 570663 699954
rect 31201 699896 31206 699952
rect 31262 699896 570602 699952
rect 570658 699896 570663 699952
rect 31201 699894 570663 699896
rect 31201 699891 31267 699894
rect 570597 699891 570663 699894
rect 26141 699818 26207 699821
rect 565077 699818 565143 699821
rect 26141 699816 565143 699818
rect 26141 699760 26146 699816
rect 26202 699760 565082 699816
rect 565138 699760 565143 699816
rect 26141 699758 565143 699760
rect 26141 699755 26207 699758
rect 565077 699755 565143 699758
rect 453941 699548 454007 699549
rect 453941 699546 453988 699548
rect 453896 699544 453988 699546
rect 453896 699488 453946 699544
rect 453896 699486 453988 699488
rect 453941 699484 453988 699486
rect 454052 699484 454058 699548
rect 453941 699483 454007 699484
rect 11605 699410 11671 699413
rect 13854 699410 13860 699412
rect 11605 699408 13860 699410
rect 11605 699352 11610 699408
rect 11666 699352 13860 699408
rect 11605 699350 13860 699352
rect 11605 699347 11671 699350
rect 13854 699348 13860 699350
rect 13924 699348 13930 699412
rect 41045 699410 41111 699413
rect 43110 699410 43116 699412
rect 41045 699408 43116 699410
rect 41045 699352 41050 699408
rect 41106 699352 43116 699408
rect 41045 699350 43116 699352
rect 41045 699347 41111 699350
rect 43110 699348 43116 699350
rect 43180 699348 43186 699412
rect 50889 699410 50955 699413
rect 52862 699410 52868 699412
rect 50889 699408 52868 699410
rect 50889 699352 50894 699408
rect 50950 699352 52868 699408
rect 50889 699350 52868 699352
rect 50889 699347 50955 699350
rect 52862 699348 52868 699350
rect 52932 699348 52938 699412
rect 55765 699410 55831 699413
rect 124581 699412 124647 699413
rect 60222 699410 60228 699412
rect 55765 699408 60228 699410
rect 55765 699352 55770 699408
rect 55826 699352 60228 699408
rect 55765 699350 60228 699352
rect 55765 699347 55831 699350
rect 60222 699348 60228 699350
rect 60292 699348 60298 699412
rect 124581 699408 124628 699412
rect 124692 699410 124698 699412
rect 326245 699410 326311 699413
rect 418705 699412 418771 699413
rect 433425 699412 433491 699413
rect 462865 699412 462931 699413
rect 418654 699410 418660 699412
rect 124581 699352 124586 699408
rect 124581 699348 124628 699352
rect 124692 699350 124738 699410
rect 251130 699350 260850 699410
rect 124692 699348 124698 699350
rect 124581 699347 124647 699348
rect 124438 699076 124444 699140
rect 124508 699138 124514 699140
rect 251130 699138 251190 699350
rect 260790 699274 260850 699350
rect 325650 699408 326311 699410
rect 325650 699352 326250 699408
rect 326306 699352 326311 699408
rect 325650 699350 326311 699352
rect 418614 699350 418660 699410
rect 418724 699408 418771 699412
rect 433374 699410 433380 699412
rect 418766 699352 418771 699408
rect 325650 699274 325710 699350
rect 326245 699347 326311 699350
rect 418654 699348 418660 699350
rect 418724 699348 418771 699352
rect 433334 699350 433380 699410
rect 433444 699408 433491 699412
rect 462814 699410 462820 699412
rect 433486 699352 433491 699408
rect 433374 699348 433380 699350
rect 433444 699348 433491 699352
rect 462774 699350 462820 699410
rect 462884 699408 462931 699412
rect 462926 699352 462931 699408
rect 462814 699348 462820 699350
rect 462884 699348 462931 699352
rect 418705 699347 418771 699348
rect 433425 699347 433491 699348
rect 462865 699347 462931 699348
rect 492581 699412 492647 699413
rect 492581 699408 492628 699412
rect 492692 699410 492698 699412
rect 492581 699352 492586 699408
rect 492581 699348 492628 699352
rect 492692 699350 492738 699410
rect 492692 699348 492698 699350
rect 510654 699348 510660 699412
rect 510724 699410 510730 699412
rect 511993 699410 512059 699413
rect 510724 699408 512059 699410
rect 510724 699352 511998 699408
rect 512054 699352 512059 699408
rect 510724 699350 512059 699352
rect 510724 699348 510730 699350
rect 492581 699347 492647 699348
rect 511993 699347 512059 699350
rect 539910 699348 539916 699412
rect 539980 699410 539986 699412
rect 541525 699410 541591 699413
rect 539980 699408 541591 699410
rect 539980 699352 541530 699408
rect 541586 699352 541591 699408
rect 539980 699350 541591 699352
rect 539980 699348 539986 699350
rect 541525 699347 541591 699350
rect 260790 699214 325710 699274
rect 124508 699078 251190 699138
rect 124508 699076 124514 699078
rect 259126 699076 259132 699140
rect 259196 699138 259202 699140
rect 580257 699138 580323 699141
rect 259196 699136 580323 699138
rect 259196 699080 580262 699136
rect 580318 699080 580323 699136
rect 259196 699078 580323 699080
rect 259196 699076 259202 699078
rect 580257 699075 580323 699078
rect 3785 699002 3851 699005
rect 510654 699002 510660 699004
rect 3785 699000 510660 699002
rect 3785 698944 3790 699000
rect 3846 698944 510660 699000
rect 3785 698942 510660 698944
rect 3785 698939 3851 698942
rect 510654 698940 510660 698942
rect 510724 698940 510730 699004
rect 60222 698804 60228 698868
rect 60292 698866 60298 698868
rect 569309 698866 569375 698869
rect 60292 698864 569375 698866
rect 60292 698808 569314 698864
rect 569370 698808 569375 698864
rect 60292 698806 569375 698808
rect 60292 698804 60298 698806
rect 569309 698803 569375 698806
rect 52862 698668 52868 698732
rect 52932 698730 52938 698732
rect 565169 698730 565235 698733
rect 52932 698728 565235 698730
rect 52932 698672 565174 698728
rect 565230 698672 565235 698728
rect 52932 698670 565235 698672
rect 52932 698668 52938 698670
rect 565169 698667 565235 698670
rect 43110 698532 43116 698596
rect 43180 698594 43186 698596
rect 566641 698594 566707 698597
rect 43180 698592 566707 698594
rect 43180 698536 566646 698592
rect 566702 698536 566707 698592
rect 43180 698534 566707 698536
rect 43180 698532 43186 698534
rect 566641 698531 566707 698534
rect 3509 698458 3575 698461
rect 539910 698458 539916 698460
rect 3509 698456 539916 698458
rect 3509 698400 3514 698456
rect 3570 698400 539916 698456
rect 3509 698398 539916 698400
rect 3509 698395 3575 698398
rect 539910 698396 539916 698398
rect 539980 698396 539986 698460
rect 13854 698260 13860 698324
rect 13924 698322 13930 698324
rect 566457 698322 566523 698325
rect 13924 698320 566523 698322
rect 13924 698264 566462 698320
rect 566518 698264 566523 698320
rect 13924 698262 566523 698264
rect 13924 698260 13930 698262
rect 566457 698259 566523 698262
rect 1853 698186 1919 698189
rect 418654 698186 418660 698188
rect 1853 698184 418660 698186
rect 1853 698128 1858 698184
rect 1914 698128 418660 698184
rect 1853 698126 418660 698128
rect 1853 698123 1919 698126
rect 418654 698124 418660 698126
rect 418724 698124 418730 698188
rect 2681 698050 2747 698053
rect 433374 698050 433380 698052
rect 2681 698048 433380 698050
rect 2681 697992 2686 698048
rect 2742 697992 433380 698048
rect 2681 697990 433380 697992
rect 2681 697987 2747 697990
rect 433374 697988 433380 697990
rect 433444 697988 433450 698052
rect 3049 697914 3115 697917
rect 124438 697914 124444 697916
rect 3049 697912 124444 697914
rect 3049 697856 3054 697912
rect 3110 697856 124444 697912
rect 3049 697854 124444 697856
rect 3049 697851 3115 697854
rect 124438 697852 124444 697854
rect 124508 697852 124514 697916
rect 124622 697852 124628 697916
rect 124692 697914 124698 697916
rect 572069 697914 572135 697917
rect 124692 697912 572135 697914
rect 124692 697856 572074 697912
rect 572130 697856 572135 697912
rect 124692 697854 572135 697856
rect 124692 697852 124698 697854
rect 572069 697851 572135 697854
rect 2497 697778 2563 697781
rect 462814 697778 462820 697780
rect 2497 697776 462820 697778
rect 2497 697720 2502 697776
rect 2558 697720 462820 697776
rect 2497 697718 462820 697720
rect 2497 697715 2563 697718
rect 462814 697716 462820 697718
rect 462884 697716 462890 697780
rect 381 697642 447 697645
rect 492622 697642 492628 697644
rect 381 697640 492628 697642
rect 381 697584 386 697640
rect 442 697584 492628 697640
rect 381 697582 492628 697584
rect 381 697579 447 697582
rect 492622 697580 492628 697582
rect 492692 697580 492698 697644
rect -960 697220 480 697460
rect 580073 697234 580139 697237
rect 583520 697234 584960 697324
rect 580073 697232 584960 697234
rect 580073 697176 580078 697232
rect 580134 697176 584960 697232
rect 580073 697174 584960 697176
rect 580073 697171 580139 697174
rect 583520 697084 584960 697174
rect -960 684314 480 684404
rect 1485 684314 1551 684317
rect -960 684312 1551 684314
rect -960 684256 1490 684312
rect 1546 684256 1551 684312
rect -960 684254 1551 684256
rect -960 684164 480 684254
rect 1485 684251 1551 684254
rect 580809 683906 580875 683909
rect 583520 683906 584960 683996
rect 580809 683904 584960 683906
rect 580809 683848 580814 683904
rect 580870 683848 584960 683904
rect 580809 683846 584960 683848
rect 580809 683843 580875 683846
rect 583520 683756 584960 683846
rect -960 671258 480 671348
rect 2957 671258 3023 671261
rect -960 671256 3023 671258
rect -960 671200 2962 671256
rect 3018 671200 3023 671256
rect -960 671198 3023 671200
rect -960 671108 480 671198
rect 2957 671195 3023 671198
rect 579613 670714 579679 670717
rect 583520 670714 584960 670804
rect 579613 670712 584960 670714
rect 579613 670656 579618 670712
rect 579674 670656 584960 670712
rect 579613 670654 584960 670656
rect 579613 670651 579679 670654
rect 583520 670564 584960 670654
rect -960 658202 480 658292
rect 4245 658202 4311 658205
rect -960 658200 4311 658202
rect -960 658144 4250 658200
rect 4306 658144 4311 658200
rect -960 658142 4311 658144
rect -960 658052 480 658142
rect 4245 658139 4311 658142
rect 583520 657236 584960 657476
rect -960 644996 480 645236
rect 580165 644058 580231 644061
rect 583520 644058 584960 644148
rect 580165 644056 584960 644058
rect 580165 644000 580170 644056
rect 580226 644000 584960 644056
rect 580165 643998 584960 644000
rect 580165 643995 580231 643998
rect 583520 643908 584960 643998
rect -960 632090 480 632180
rect 1577 632090 1643 632093
rect -960 632088 1643 632090
rect -960 632032 1582 632088
rect 1638 632032 1643 632088
rect -960 632030 1643 632032
rect -960 631940 480 632030
rect 1577 632027 1643 632030
rect 580165 630866 580231 630869
rect 583520 630866 584960 630956
rect 580165 630864 584960 630866
rect 580165 630808 580170 630864
rect 580226 630808 584960 630864
rect 580165 630806 584960 630808
rect 580165 630803 580231 630806
rect 583520 630716 584960 630806
rect -960 619170 480 619260
rect 4061 619170 4127 619173
rect -960 619168 4127 619170
rect -960 619112 4066 619168
rect 4122 619112 4127 619168
rect -960 619110 4127 619112
rect -960 619020 480 619110
rect 4061 619107 4127 619110
rect 580165 617538 580231 617541
rect 583520 617538 584960 617628
rect 580165 617536 584960 617538
rect 580165 617480 580170 617536
rect 580226 617480 584960 617536
rect 580165 617478 584960 617480
rect 580165 617475 580231 617478
rect 583520 617388 584960 617478
rect -960 606114 480 606204
rect 933 606114 999 606117
rect -960 606112 999 606114
rect -960 606056 938 606112
rect 994 606056 999 606112
rect -960 606054 999 606056
rect -960 605964 480 606054
rect 933 606051 999 606054
rect 583520 604060 584960 604300
rect -960 592908 480 593148
rect 580165 591018 580231 591021
rect 583520 591018 584960 591108
rect 580165 591016 584960 591018
rect 580165 590960 580170 591016
rect 580226 590960 584960 591016
rect 580165 590958 584960 590960
rect 580165 590955 580231 590958
rect 583520 590868 584960 590958
rect -960 580002 480 580092
rect 1669 580002 1735 580005
rect -960 580000 1735 580002
rect -960 579944 1674 580000
rect 1730 579944 1735 580000
rect -960 579942 1735 579944
rect -960 579852 480 579942
rect 1669 579939 1735 579942
rect 580809 577690 580875 577693
rect 583520 577690 584960 577780
rect 580809 577688 584960 577690
rect 580809 577632 580814 577688
rect 580870 577632 584960 577688
rect 580809 577630 584960 577632
rect 580809 577627 580875 577630
rect 583520 577540 584960 577630
rect -960 566946 480 567036
rect 3049 566946 3115 566949
rect -960 566944 3115 566946
rect -960 566888 3054 566944
rect 3110 566888 3115 566944
rect -960 566886 3115 566888
rect -960 566796 480 566886
rect 3049 566883 3115 566886
rect 580165 564362 580231 564365
rect 583520 564362 584960 564452
rect 580165 564360 584960 564362
rect 580165 564304 580170 564360
rect 580226 564304 584960 564360
rect 580165 564302 584960 564304
rect 580165 564299 580231 564302
rect 583520 564212 584960 564302
rect -960 553890 480 553980
rect 841 553890 907 553893
rect -960 553888 907 553890
rect -960 553832 846 553888
rect 902 553832 907 553888
rect -960 553830 907 553832
rect -960 553740 480 553830
rect 841 553827 907 553830
rect 583520 551020 584960 551260
rect -960 540684 480 540924
rect 580165 537842 580231 537845
rect 583520 537842 584960 537932
rect 580165 537840 584960 537842
rect 580165 537784 580170 537840
rect 580226 537784 584960 537840
rect 580165 537782 584960 537784
rect 580165 537779 580231 537782
rect 583520 537692 584960 537782
rect -960 527914 480 528004
rect 1761 527914 1827 527917
rect -960 527912 1827 527914
rect -960 527856 1766 527912
rect 1822 527856 1827 527912
rect -960 527854 1827 527856
rect -960 527764 480 527854
rect 1761 527851 1827 527854
rect 580717 524514 580783 524517
rect 583520 524514 584960 524604
rect 580717 524512 584960 524514
rect 580717 524456 580722 524512
rect 580778 524456 584960 524512
rect 580717 524454 584960 524456
rect 580717 524451 580783 524454
rect 583520 524364 584960 524454
rect -960 514858 480 514948
rect 2773 514858 2839 514861
rect -960 514856 2839 514858
rect -960 514800 2778 514856
rect 2834 514800 2839 514856
rect -960 514798 2839 514800
rect -960 514708 480 514798
rect 2773 514795 2839 514798
rect 580165 511322 580231 511325
rect 583520 511322 584960 511412
rect 580165 511320 584960 511322
rect 580165 511264 580170 511320
rect 580226 511264 584960 511320
rect 580165 511262 584960 511264
rect 580165 511259 580231 511262
rect 583520 511172 584960 511262
rect -960 501802 480 501892
rect 749 501802 815 501805
rect -960 501800 815 501802
rect -960 501744 754 501800
rect 810 501744 815 501800
rect -960 501742 815 501744
rect -960 501652 480 501742
rect 749 501739 815 501742
rect 583520 497844 584960 498084
rect -960 488596 480 488836
rect 579613 484666 579679 484669
rect 583520 484666 584960 484756
rect 579613 484664 584960 484666
rect 579613 484608 579618 484664
rect 579674 484608 584960 484664
rect 579613 484606 584960 484608
rect 579613 484603 579679 484606
rect 583520 484516 584960 484606
rect -960 475690 480 475780
rect 1853 475690 1919 475693
rect -960 475688 1919 475690
rect -960 475632 1858 475688
rect 1914 475632 1919 475688
rect -960 475630 1919 475632
rect -960 475540 480 475630
rect 1853 475627 1919 475630
rect 579797 471474 579863 471477
rect 583520 471474 584960 471564
rect 579797 471472 584960 471474
rect 579797 471416 579802 471472
rect 579858 471416 584960 471472
rect 579797 471414 584960 471416
rect 579797 471411 579863 471414
rect 583520 471324 584960 471414
rect -960 462634 480 462724
rect 3141 462634 3207 462637
rect -960 462632 3207 462634
rect -960 462576 3146 462632
rect 3202 462576 3207 462632
rect -960 462574 3207 462576
rect -960 462484 480 462574
rect 3141 462571 3207 462574
rect 580625 458146 580691 458149
rect 583520 458146 584960 458236
rect 580625 458144 584960 458146
rect 580625 458088 580630 458144
rect 580686 458088 584960 458144
rect 580625 458086 584960 458088
rect 580625 458083 580691 458086
rect 583520 457996 584960 458086
rect -960 449578 480 449668
rect 1945 449578 2011 449581
rect -960 449576 2011 449578
rect -960 449520 1950 449576
rect 2006 449520 2011 449576
rect -960 449518 2011 449520
rect -960 449428 480 449518
rect 1945 449515 2011 449518
rect 583520 444668 584960 444908
rect -960 436508 480 436748
rect 579705 431626 579771 431629
rect 583520 431626 584960 431716
rect 579705 431624 584960 431626
rect 579705 431568 579710 431624
rect 579766 431568 584960 431624
rect 579705 431566 584960 431568
rect 579705 431563 579771 431566
rect 583520 431476 584960 431566
rect -960 423602 480 423692
rect 2681 423602 2747 423605
rect -960 423600 2747 423602
rect -960 423544 2686 423600
rect 2742 423544 2747 423600
rect -960 423542 2747 423544
rect -960 423452 480 423542
rect 2681 423539 2747 423542
rect 580165 418298 580231 418301
rect 583520 418298 584960 418388
rect 580165 418296 584960 418298
rect 580165 418240 580170 418296
rect 580226 418240 584960 418296
rect 580165 418238 584960 418240
rect 580165 418235 580231 418238
rect 583520 418148 584960 418238
rect -960 410546 480 410636
rect 3233 410546 3299 410549
rect -960 410544 3299 410546
rect -960 410488 3238 410544
rect 3294 410488 3299 410544
rect -960 410486 3299 410488
rect -960 410396 480 410486
rect 3233 410483 3299 410486
rect 578969 404970 579035 404973
rect 583520 404970 584960 405060
rect 578969 404968 584960 404970
rect 578969 404912 578974 404968
rect 579030 404912 584960 404968
rect 578969 404910 584960 404912
rect 578969 404907 579035 404910
rect 583520 404820 584960 404910
rect -960 397490 480 397580
rect 3325 397490 3391 397493
rect -960 397488 3391 397490
rect -960 397432 3330 397488
rect 3386 397432 3391 397488
rect -960 397430 3391 397432
rect -960 397340 480 397430
rect 3325 397427 3391 397430
rect 583520 391628 584960 391868
rect -960 384284 480 384524
rect 579613 378450 579679 378453
rect 583520 378450 584960 378540
rect 579613 378448 584960 378450
rect 579613 378392 579618 378448
rect 579674 378392 584960 378448
rect 579613 378390 584960 378392
rect 579613 378387 579679 378390
rect 583520 378300 584960 378390
rect -960 371378 480 371468
rect 2589 371378 2655 371381
rect -960 371376 2655 371378
rect -960 371320 2594 371376
rect 2650 371320 2655 371376
rect -960 371318 2655 371320
rect -960 371228 480 371318
rect 2589 371315 2655 371318
rect 578877 365122 578943 365125
rect 583520 365122 584960 365212
rect 578877 365120 584960 365122
rect 578877 365064 578882 365120
rect 578938 365064 584960 365120
rect 578877 365062 584960 365064
rect 578877 365059 578943 365062
rect 583520 364972 584960 365062
rect -960 358458 480 358548
rect 657 358458 723 358461
rect -960 358456 723 358458
rect -960 358400 662 358456
rect 718 358400 723 358456
rect -960 358398 723 358400
rect -960 358308 480 358398
rect 657 358395 723 358398
rect 580165 351930 580231 351933
rect 583520 351930 584960 352020
rect 580165 351928 584960 351930
rect 580165 351872 580170 351928
rect 580226 351872 584960 351928
rect 580165 351870 584960 351872
rect 580165 351867 580231 351870
rect 583520 351780 584960 351870
rect -960 345402 480 345492
rect 565 345402 631 345405
rect -960 345400 631 345402
rect -960 345344 570 345400
rect 626 345344 631 345400
rect -960 345342 631 345344
rect -960 345252 480 345342
rect 565 345339 631 345342
rect 583520 338452 584960 338692
rect -960 332196 480 332436
rect 580165 325274 580231 325277
rect 583520 325274 584960 325364
rect 580165 325272 584960 325274
rect 580165 325216 580170 325272
rect 580226 325216 584960 325272
rect 580165 325214 584960 325216
rect 580165 325211 580231 325214
rect 583520 325124 584960 325214
rect -960 319290 480 319380
rect 2497 319290 2563 319293
rect -960 319288 2563 319290
rect -960 319232 2502 319288
rect 2558 319232 2563 319288
rect -960 319230 2563 319232
rect -960 319140 480 319230
rect 2497 319227 2563 319230
rect 580165 312082 580231 312085
rect 583520 312082 584960 312172
rect 580165 312080 584960 312082
rect 580165 312024 580170 312080
rect 580226 312024 584960 312080
rect 580165 312022 584960 312024
rect 580165 312019 580231 312022
rect 583520 311932 584960 312022
rect -960 306234 480 306324
rect 2405 306234 2471 306237
rect -960 306232 2471 306234
rect -960 306176 2410 306232
rect 2466 306176 2471 306232
rect -960 306174 2471 306176
rect -960 306084 480 306174
rect 2405 306171 2471 306174
rect 580165 298754 580231 298757
rect 583520 298754 584960 298844
rect 580165 298752 584960 298754
rect 580165 298696 580170 298752
rect 580226 298696 584960 298752
rect 580165 298694 584960 298696
rect 580165 298691 580231 298694
rect 583520 298604 584960 298694
rect -960 293178 480 293268
rect 3969 293178 4035 293181
rect -960 293176 4035 293178
rect -960 293120 3974 293176
rect 4030 293120 4035 293176
rect -960 293118 4035 293120
rect -960 293028 480 293118
rect 3969 293115 4035 293118
rect 583520 285276 584960 285516
rect -960 279972 480 280212
rect 579613 272234 579679 272237
rect 583520 272234 584960 272324
rect 579613 272232 584960 272234
rect 579613 272176 579618 272232
rect 579674 272176 584960 272232
rect 579613 272174 584960 272176
rect 579613 272171 579679 272174
rect 583520 272084 584960 272174
rect -960 267202 480 267292
rect 2221 267202 2287 267205
rect -960 267200 2287 267202
rect -960 267144 2226 267200
rect 2282 267144 2287 267200
rect -960 267142 2287 267144
rect -960 267052 480 267142
rect 2221 267139 2287 267142
rect 580625 258906 580691 258909
rect 583520 258906 584960 258996
rect 580625 258904 584960 258906
rect 580625 258848 580630 258904
rect 580686 258848 584960 258904
rect 580625 258846 584960 258848
rect 580625 258843 580691 258846
rect 583520 258756 584960 258846
rect -960 254146 480 254236
rect 4061 254146 4127 254149
rect -960 254144 4127 254146
rect -960 254088 4066 254144
rect 4122 254088 4127 254144
rect -960 254086 4127 254088
rect -960 253996 480 254086
rect 4061 254083 4127 254086
rect 580165 245578 580231 245581
rect 583520 245578 584960 245668
rect 580165 245576 584960 245578
rect 580165 245520 580170 245576
rect 580226 245520 584960 245576
rect 580165 245518 584960 245520
rect 580165 245515 580231 245518
rect 583520 245428 584960 245518
rect -960 241090 480 241180
rect 565 241090 631 241093
rect -960 241088 631 241090
rect -960 241032 570 241088
rect 626 241032 631 241088
rect -960 241030 631 241032
rect -960 240940 480 241030
rect 565 241027 631 241030
rect 579981 232386 580047 232389
rect 583520 232386 584960 232476
rect 579981 232384 584960 232386
rect 579981 232328 579986 232384
rect 580042 232328 584960 232384
rect 579981 232326 584960 232328
rect 579981 232323 580047 232326
rect 583520 232236 584960 232326
rect -960 227884 480 228124
rect 580533 219058 580599 219061
rect 583520 219058 584960 219148
rect 580533 219056 584960 219058
rect 580533 219000 580538 219056
rect 580594 219000 584960 219056
rect 580533 218998 584960 219000
rect 580533 218995 580599 218998
rect 583520 218908 584960 218998
rect -960 214978 480 215068
rect 565 214978 631 214981
rect -960 214976 631 214978
rect -960 214920 570 214976
rect 626 214920 631 214976
rect -960 214918 631 214920
rect -960 214828 480 214918
rect 565 214915 631 214918
rect 580165 205730 580231 205733
rect 583520 205730 584960 205820
rect 580165 205728 584960 205730
rect 580165 205672 580170 205728
rect 580226 205672 584960 205728
rect 580165 205670 584960 205672
rect 580165 205667 580231 205670
rect 583520 205580 584960 205670
rect -960 201922 480 202012
rect 565 201922 631 201925
rect -960 201920 631 201922
rect -960 201864 570 201920
rect 626 201864 631 201920
rect -960 201862 631 201864
rect -960 201772 480 201862
rect 565 201859 631 201862
rect 580441 192538 580507 192541
rect 583520 192538 584960 192628
rect 580441 192536 584960 192538
rect 580441 192480 580446 192536
rect 580502 192480 584960 192536
rect 580441 192478 584960 192480
rect 580441 192475 580507 192478
rect 583520 192388 584960 192478
rect -960 188866 480 188956
rect 2313 188866 2379 188869
rect -960 188864 2379 188866
rect -960 188808 2318 188864
rect 2374 188808 2379 188864
rect -960 188806 2379 188808
rect -960 188716 480 188806
rect 2313 188803 2379 188806
rect 580349 179210 580415 179213
rect 583520 179210 584960 179300
rect 580349 179208 584960 179210
rect 580349 179152 580354 179208
rect 580410 179152 584960 179208
rect 580349 179150 584960 179152
rect 580349 179147 580415 179150
rect 583520 179060 584960 179150
rect -960 175796 480 176036
rect 580165 165882 580231 165885
rect 583520 165882 584960 165972
rect 580165 165880 584960 165882
rect 580165 165824 580170 165880
rect 580226 165824 584960 165880
rect 580165 165822 584960 165824
rect 580165 165819 580231 165822
rect 583520 165732 584960 165822
rect 197 163434 263 163437
rect 197 163432 306 163434
rect 197 163376 202 163432
rect 258 163376 306 163432
rect 197 163371 306 163376
rect 246 163026 306 163371
rect 246 162980 674 163026
rect -960 162966 674 162980
rect -960 162890 480 162966
rect 614 162890 674 162966
rect -960 162830 674 162890
rect -960 162740 480 162830
rect 579797 152690 579863 152693
rect 583520 152690 584960 152780
rect 579797 152688 584960 152690
rect 579797 152632 579802 152688
rect 579858 152632 584960 152688
rect 579797 152630 584960 152632
rect 579797 152627 579863 152630
rect 583520 152540 584960 152630
rect -960 149834 480 149924
rect 3877 149834 3943 149837
rect -960 149832 3943 149834
rect -960 149776 3882 149832
rect 3938 149776 3943 149832
rect -960 149774 3943 149776
rect -960 149684 480 149774
rect 3877 149771 3943 149774
rect 580165 139362 580231 139365
rect 583520 139362 584960 139452
rect 580165 139360 584960 139362
rect 580165 139304 580170 139360
rect 580226 139304 584960 139360
rect 580165 139302 584960 139304
rect 580165 139299 580231 139302
rect 583520 139212 584960 139302
rect -960 136778 480 136868
rect 3785 136778 3851 136781
rect -960 136776 3851 136778
rect -960 136720 3790 136776
rect 3846 136720 3851 136776
rect -960 136718 3851 136720
rect -960 136628 480 136718
rect 3785 136715 3851 136718
rect 580165 126034 580231 126037
rect 583520 126034 584960 126124
rect 580165 126032 584960 126034
rect 580165 125976 580170 126032
rect 580226 125976 584960 126032
rect 580165 125974 584960 125976
rect 580165 125971 580231 125974
rect 583520 125884 584960 125974
rect -960 123572 480 123812
rect 580165 112842 580231 112845
rect 583520 112842 584960 112932
rect 580165 112840 584960 112842
rect 580165 112784 580170 112840
rect 580226 112784 584960 112840
rect 580165 112782 584960 112784
rect 580165 112779 580231 112782
rect 583520 112692 584960 112782
rect 105 111210 171 111213
rect 105 111208 306 111210
rect 105 111152 110 111208
rect 166 111152 306 111208
rect 105 111150 306 111152
rect 105 111147 171 111150
rect 246 110802 306 111150
rect 246 110756 674 110802
rect -960 110742 674 110756
rect -960 110666 480 110742
rect 614 110666 674 110742
rect -960 110606 674 110666
rect -960 110516 480 110606
rect 580165 99514 580231 99517
rect 583520 99514 584960 99604
rect 580165 99512 584960 99514
rect 580165 99456 580170 99512
rect 580226 99456 584960 99512
rect 580165 99454 584960 99456
rect 580165 99451 580231 99454
rect 583520 99364 584960 99454
rect -960 97610 480 97700
rect 2129 97610 2195 97613
rect -960 97608 2195 97610
rect -960 97552 2134 97608
rect 2190 97552 2195 97608
rect -960 97550 2195 97552
rect -960 97460 480 97550
rect 2129 97547 2195 97550
rect 580165 86186 580231 86189
rect 583520 86186 584960 86276
rect 580165 86184 584960 86186
rect 580165 86128 580170 86184
rect 580226 86128 584960 86184
rect 580165 86126 584960 86128
rect 580165 86123 580231 86126
rect 583520 86036 584960 86126
rect -960 84690 480 84780
rect 3693 84690 3759 84693
rect -960 84688 3759 84690
rect -960 84632 3698 84688
rect 3754 84632 3759 84688
rect -960 84630 3759 84632
rect -960 84540 480 84630
rect 3693 84627 3759 84630
rect 579981 72994 580047 72997
rect 583520 72994 584960 73084
rect 579981 72992 584960 72994
rect 579981 72936 579986 72992
rect 580042 72936 584960 72992
rect 579981 72934 584960 72936
rect 579981 72931 580047 72934
rect 583520 72844 584960 72934
rect 13 71906 79 71909
rect 13 71904 122 71906
rect 13 71848 18 71904
rect 74 71848 122 71904
rect 13 71843 122 71848
rect 62 71770 122 71843
rect 62 71724 674 71770
rect -960 71710 674 71724
rect -960 71634 480 71710
rect 614 71634 674 71710
rect -960 71574 674 71634
rect -960 71484 480 71574
rect 580165 59666 580231 59669
rect 583520 59666 584960 59756
rect 580165 59664 584960 59666
rect 580165 59608 580170 59664
rect 580226 59608 584960 59664
rect 580165 59606 584960 59608
rect 580165 59603 580231 59606
rect 583520 59516 584960 59606
rect -960 58578 480 58668
rect 3601 58578 3667 58581
rect -960 58576 3667 58578
rect -960 58520 3606 58576
rect 3662 58520 3667 58576
rect -960 58518 3667 58520
rect -960 58428 480 58518
rect 3601 58515 3667 58518
rect 580165 46338 580231 46341
rect 583520 46338 584960 46428
rect 580165 46336 584960 46338
rect 580165 46280 580170 46336
rect 580226 46280 584960 46336
rect 580165 46278 584960 46280
rect 580165 46275 580231 46278
rect 583520 46188 584960 46278
rect -960 45522 480 45612
rect 3509 45522 3575 45525
rect -960 45520 3575 45522
rect -960 45464 3514 45520
rect 3570 45464 3575 45520
rect -960 45462 3575 45464
rect -960 45372 480 45462
rect 3509 45459 3575 45462
rect 580165 33146 580231 33149
rect 583520 33146 584960 33236
rect 580165 33144 584960 33146
rect 580165 33088 580170 33144
rect 580226 33088 584960 33144
rect 580165 33086 584960 33088
rect 580165 33083 580231 33086
rect 583520 32996 584960 33086
rect -960 32466 480 32556
rect 2037 32466 2103 32469
rect -960 32464 2103 32466
rect -960 32408 2042 32464
rect 2098 32408 2103 32464
rect -960 32406 2103 32408
rect -960 32316 480 32406
rect 2037 32403 2103 32406
rect 580165 19818 580231 19821
rect 583520 19818 584960 19908
rect 580165 19816 584960 19818
rect 580165 19760 580170 19816
rect 580226 19760 584960 19816
rect 580165 19758 584960 19760
rect 580165 19755 580231 19758
rect 583520 19668 584960 19758
rect -960 19410 480 19500
rect 3417 19410 3483 19413
rect -960 19408 3483 19410
rect -960 19352 3422 19408
rect 3478 19352 3483 19408
rect -960 19350 3483 19352
rect -960 19260 480 19350
rect 3417 19347 3483 19350
rect 580257 6626 580323 6629
rect 583520 6626 584960 6716
rect 580257 6624 584960 6626
rect -960 6490 480 6580
rect 580257 6568 580262 6624
rect 580318 6568 584960 6624
rect 580257 6566 584960 6568
rect 580257 6563 580323 6566
rect 2957 6490 3023 6493
rect -960 6488 3023 6490
rect -960 6432 2962 6488
rect 3018 6432 3023 6488
rect 583520 6476 584960 6566
rect -960 6430 3023 6432
rect -960 6340 480 6430
rect 2957 6427 3023 6430
rect 531078 1458 531084 1460
rect 514710 1398 531084 1458
rect 514710 645 514770 1398
rect 531078 1396 531084 1398
rect 531148 1396 531154 1460
rect 542854 1124 542860 1188
rect 542924 1186 542930 1188
rect 542924 1126 553410 1186
rect 542924 1124 542930 1126
rect 542486 914 542492 916
rect 532006 854 542492 914
rect 4061 642 4127 645
rect 7833 642 7899 645
rect 4061 640 7899 642
rect 4061 584 4066 640
rect 4122 584 7838 640
rect 7894 584 7899 640
rect 4061 582 7899 584
rect 4061 579 4127 582
rect 7833 579 7899 582
rect 9949 642 10015 645
rect 13721 642 13787 645
rect 9949 640 13787 642
rect 9949 584 9954 640
rect 10010 584 13726 640
rect 13782 584 13787 640
rect 9949 582 13787 584
rect 9949 579 10015 582
rect 13721 579 13787 582
rect 26509 642 26575 645
rect 28717 642 28783 645
rect 30281 642 30347 645
rect 26509 640 28783 642
rect 26509 584 26514 640
rect 26570 584 28722 640
rect 28778 584 28783 640
rect 26509 582 28783 584
rect 26509 579 26575 582
rect 28717 579 28783 582
rect 29134 640 30347 642
rect 29134 584 30286 640
rect 30342 584 30347 640
rect 29134 582 30347 584
rect 27889 506 27955 509
rect 29134 506 29194 582
rect 30281 579 30347 582
rect 31293 642 31359 645
rect 33593 642 33659 645
rect 35985 642 36051 645
rect 38469 642 38535 645
rect 31293 640 31770 642
rect 31293 584 31298 640
rect 31354 584 31770 640
rect 31293 582 31770 584
rect 31293 579 31359 582
rect 27889 504 29194 506
rect 27889 448 27894 504
rect 27950 448 29194 504
rect 27889 446 29194 448
rect 31710 506 31770 582
rect 33593 640 34530 642
rect 33593 584 33598 640
rect 33654 584 34530 640
rect 33593 582 34530 584
rect 33593 579 33659 582
rect 33869 506 33935 509
rect 31710 504 33935 506
rect 31710 448 33874 504
rect 33930 448 33935 504
rect 31710 446 33935 448
rect 34470 506 34530 582
rect 35985 640 38535 642
rect 35985 584 35990 640
rect 36046 584 38474 640
rect 38530 584 38535 640
rect 35985 582 38535 584
rect 35985 579 36051 582
rect 38469 579 38535 582
rect 52545 642 52611 645
rect 54201 642 54267 645
rect 52545 640 54267 642
rect 52545 584 52550 640
rect 52606 584 54206 640
rect 54262 584 54267 640
rect 52545 582 54267 584
rect 52545 579 52611 582
rect 54201 579 54267 582
rect 56041 642 56107 645
rect 57605 642 57671 645
rect 56041 640 57671 642
rect 56041 584 56046 640
rect 56102 584 57610 640
rect 57666 584 57671 640
rect 56041 582 57671 584
rect 56041 579 56107 582
rect 57605 579 57671 582
rect 58433 642 58499 645
rect 59813 642 59879 645
rect 58433 640 59879 642
rect 58433 584 58438 640
rect 58494 584 59818 640
rect 59874 584 59879 640
rect 58433 582 59879 584
rect 58433 579 58499 582
rect 59813 579 59879 582
rect 60825 642 60891 645
rect 62113 642 62179 645
rect 60825 640 62179 642
rect 60825 584 60830 640
rect 60886 584 62118 640
rect 62174 584 62179 640
rect 60825 582 62179 584
rect 60825 579 60891 582
rect 62113 579 62179 582
rect 142061 642 142127 645
rect 143441 642 143507 645
rect 144729 642 144795 645
rect 142061 640 142170 642
rect 142061 584 142066 640
rect 142122 584 142170 640
rect 142061 579 142170 584
rect 143441 640 144795 642
rect 143441 584 143446 640
rect 143502 584 144734 640
rect 144790 584 144795 640
rect 143441 582 144795 584
rect 143441 579 143507 582
rect 144729 579 144795 582
rect 145741 642 145807 645
rect 147121 642 147187 645
rect 145741 640 147187 642
rect 145741 584 145746 640
rect 145802 584 147126 640
rect 147182 584 147187 640
rect 145741 582 147187 584
rect 145741 579 145807 582
rect 147121 579 147187 582
rect 148961 642 149027 645
rect 150617 642 150683 645
rect 151813 642 151879 645
rect 148961 640 150683 642
rect 148961 584 148966 640
rect 149022 584 150622 640
rect 150678 584 150683 640
rect 148961 582 150683 584
rect 148961 579 149027 582
rect 150617 579 150683 582
rect 151678 640 151879 642
rect 151678 584 151818 640
rect 151874 584 151879 640
rect 151678 582 151879 584
rect 36169 506 36235 509
rect 34470 504 36235 506
rect 34470 448 36174 504
rect 36230 448 36235 504
rect 34470 446 36235 448
rect 27889 443 27955 446
rect 33869 443 33935 446
rect 36169 443 36235 446
rect 53557 506 53623 509
rect 55305 506 55371 509
rect 53557 504 55371 506
rect 53557 448 53562 504
rect 53618 448 55310 504
rect 55366 448 55371 504
rect 53557 446 55371 448
rect 53557 443 53623 446
rect 55305 443 55371 446
rect 57421 506 57487 509
rect 58801 506 58867 509
rect 57421 504 58867 506
rect 57421 448 57426 504
rect 57482 448 58806 504
rect 58862 448 58867 504
rect 57421 446 58867 448
rect 57421 443 57487 446
rect 58801 443 58867 446
rect 59445 506 59511 509
rect 61101 506 61167 509
rect 59445 504 61167 506
rect 59445 448 59450 504
rect 59506 448 61106 504
rect 61162 448 61167 504
rect 59445 446 61167 448
rect 142110 506 142170 579
rect 143717 506 143783 509
rect 142110 504 143783 506
rect 142110 448 143722 504
rect 143778 448 143783 504
rect 142110 446 143783 448
rect 59445 443 59511 446
rect 61101 443 61167 446
rect 143717 443 143783 446
rect 147765 506 147831 509
rect 149329 506 149395 509
rect 147765 504 149395 506
rect 147765 448 147770 504
rect 147826 448 149334 504
rect 149390 448 149395 504
rect 147765 446 149395 448
rect 147765 443 147831 446
rect 149329 443 149395 446
rect 150249 506 150315 509
rect 151678 506 151738 582
rect 151813 579 151879 582
rect 164785 642 164851 645
rect 167361 642 167427 645
rect 164785 640 167427 642
rect 164785 584 164790 640
rect 164846 584 167366 640
rect 167422 584 167427 640
rect 164785 582 167427 584
rect 164785 579 164851 582
rect 167361 579 167427 582
rect 169477 642 169543 645
rect 171961 642 172027 645
rect 169477 640 172027 642
rect 169477 584 169482 640
rect 169538 584 171966 640
rect 172022 584 172027 640
rect 169477 582 172027 584
rect 169477 579 169543 582
rect 171961 579 172027 582
rect 172973 642 173039 645
rect 175457 642 175523 645
rect 172973 640 175523 642
rect 172973 584 172978 640
rect 173034 584 175462 640
rect 175518 584 175523 640
rect 172973 582 175523 584
rect 172973 579 173039 582
rect 175457 579 175523 582
rect 176377 642 176443 645
rect 179045 642 179111 645
rect 180241 642 180307 645
rect 176377 640 179111 642
rect 176377 584 176382 640
rect 176438 584 179050 640
rect 179106 584 179111 640
rect 176377 582 179111 584
rect 176377 579 176443 582
rect 179045 579 179111 582
rect 179370 640 180307 642
rect 179370 584 180246 640
rect 180302 584 180307 640
rect 179370 582 180307 584
rect 150249 504 151738 506
rect 150249 448 150254 504
rect 150310 448 151738 504
rect 150249 446 151738 448
rect 173893 506 173959 509
rect 176837 506 176903 509
rect 173893 504 176903 506
rect 173893 448 173898 504
rect 173954 448 176842 504
rect 176898 448 176903 504
rect 173893 446 176903 448
rect 150249 443 150315 446
rect 173893 443 173959 446
rect 176837 443 176903 446
rect 177481 506 177547 509
rect 179370 506 179430 582
rect 180241 579 180307 582
rect 182081 642 182147 645
rect 184933 642 184999 645
rect 182081 640 184999 642
rect 182081 584 182086 640
rect 182142 584 184938 640
rect 184994 584 184999 640
rect 182081 582 184999 584
rect 182081 579 182147 582
rect 184933 579 184999 582
rect 192293 642 192359 645
rect 195605 642 195671 645
rect 197905 642 197971 645
rect 192293 640 195671 642
rect 192293 584 192298 640
rect 192354 584 195610 640
rect 195666 584 195671 640
rect 192293 582 195671 584
rect 192293 579 192359 582
rect 195605 579 195671 582
rect 197310 640 197971 642
rect 197310 584 197910 640
rect 197966 584 197971 640
rect 197310 582 197971 584
rect 177481 504 179430 506
rect 177481 448 177486 504
rect 177542 448 179430 504
rect 177481 446 179430 448
rect 186589 506 186655 509
rect 189901 506 189967 509
rect 186589 504 189967 506
rect 186589 448 186594 504
rect 186650 448 189906 504
rect 189962 448 189967 504
rect 186589 446 189967 448
rect 177481 443 177547 446
rect 186589 443 186655 446
rect 189901 443 189967 446
rect 194041 506 194107 509
rect 197310 506 197370 582
rect 197905 579 197971 582
rect 200021 642 200087 645
rect 203885 642 203951 645
rect 200021 640 203951 642
rect 200021 584 200026 640
rect 200082 584 203890 640
rect 203946 584 203951 640
rect 200021 582 203951 584
rect 200021 579 200087 582
rect 203885 579 203951 582
rect 204161 642 204227 645
rect 207381 642 207447 645
rect 204161 640 207447 642
rect 204161 584 204166 640
rect 204222 584 207386 640
rect 207442 584 207447 640
rect 204161 582 207447 584
rect 204161 579 204227 582
rect 207381 579 207447 582
rect 208209 642 208275 645
rect 208393 642 208459 645
rect 208209 640 208459 642
rect 208209 584 208214 640
rect 208270 584 208398 640
rect 208454 584 208459 640
rect 208209 582 208459 584
rect 208209 579 208275 582
rect 208393 579 208459 582
rect 209313 642 209379 645
rect 213361 642 213427 645
rect 209313 640 213427 642
rect 209313 584 209318 640
rect 209374 584 213366 640
rect 213422 584 213427 640
rect 209313 582 213427 584
rect 209313 579 209379 582
rect 213361 579 213427 582
rect 216121 642 216187 645
rect 220445 642 220511 645
rect 216121 640 220511 642
rect 216121 584 216126 640
rect 216182 584 220450 640
rect 220506 584 220511 640
rect 216121 582 220511 584
rect 216121 579 216187 582
rect 220445 579 220511 582
rect 223849 642 223915 645
rect 228725 642 228791 645
rect 223849 640 228791 642
rect 223849 584 223854 640
rect 223910 584 228730 640
rect 228786 584 228791 640
rect 223849 582 228791 584
rect 223849 579 223915 582
rect 228725 579 228791 582
rect 230933 642 230999 645
rect 235809 642 235875 645
rect 230933 640 235875 642
rect 230933 584 230938 640
rect 230994 584 235814 640
rect 235870 584 235875 640
rect 230933 582 235875 584
rect 230933 579 230999 582
rect 235809 579 235875 582
rect 238845 642 238911 645
rect 244089 642 244155 645
rect 238845 640 244155 642
rect 238845 584 238850 640
rect 238906 584 244094 640
rect 244150 584 244155 640
rect 238845 582 244155 584
rect 238845 579 238911 582
rect 244089 579 244155 582
rect 249057 642 249123 645
rect 254669 642 254735 645
rect 249057 640 254735 642
rect 249057 584 249062 640
rect 249118 584 254674 640
rect 254730 584 254735 640
rect 249057 582 254735 584
rect 249057 579 249123 582
rect 254669 579 254735 582
rect 255221 642 255287 645
rect 255865 642 255931 645
rect 257061 642 257127 645
rect 255221 640 255931 642
rect 255221 584 255226 640
rect 255282 584 255870 640
rect 255926 584 255931 640
rect 255221 582 255931 584
rect 255221 579 255287 582
rect 255865 579 255931 582
rect 256650 640 257127 642
rect 256650 584 257066 640
rect 257122 584 257127 640
rect 256650 582 257127 584
rect 194041 504 197370 506
rect 194041 448 194046 504
rect 194102 448 197370 504
rect 194041 446 197370 448
rect 198917 506 198983 509
rect 201309 506 201375 509
rect 204897 506 204963 509
rect 198917 504 200866 506
rect 198917 448 198922 504
rect 198978 448 200866 504
rect 198917 446 200866 448
rect 194041 443 194107 446
rect 198917 443 198983 446
rect 32213 370 32279 373
rect 34973 370 35039 373
rect 32213 368 35039 370
rect 32213 312 32218 368
rect 32274 312 34978 368
rect 35034 312 35039 368
rect 32213 310 35039 312
rect 32213 307 32279 310
rect 34973 307 35039 310
rect 168189 370 168255 373
rect 170949 370 171015 373
rect 168189 368 171015 370
rect 168189 312 168194 368
rect 168250 312 170954 368
rect 171010 312 171015 368
rect 168189 310 171015 312
rect 168189 307 168255 310
rect 170949 307 171015 310
rect 171685 370 171751 373
rect 173985 370 174051 373
rect 171685 368 174051 370
rect 171685 312 171690 368
rect 171746 312 173990 368
rect 174046 312 174051 368
rect 171685 310 174051 312
rect 171685 307 171751 310
rect 173985 307 174051 310
rect 175181 370 175247 373
rect 177665 370 177731 373
rect 175181 368 177731 370
rect 175181 312 175186 368
rect 175242 312 177670 368
rect 177726 312 177731 368
rect 175181 310 177731 312
rect 175181 307 175247 310
rect 177665 307 177731 310
rect 178677 370 178743 373
rect 181253 370 181319 373
rect 178677 368 181319 370
rect 178677 312 178682 368
rect 178738 312 181258 368
rect 181314 312 181319 368
rect 178677 310 181319 312
rect 178677 307 178743 310
rect 181253 307 181319 310
rect 188797 370 188863 373
rect 192201 370 192267 373
rect 188797 368 192267 370
rect 188797 312 188802 368
rect 188858 312 192206 368
rect 192262 312 192267 368
rect 188797 310 192267 312
rect 188797 307 188863 310
rect 192201 307 192267 310
rect 196617 370 196683 373
rect 200113 370 200179 373
rect 196617 368 200179 370
rect 196617 312 196622 368
rect 196678 312 200118 368
rect 200174 312 200179 368
rect 196617 310 200179 312
rect 200806 370 200866 446
rect 201309 504 204963 506
rect 201309 448 201314 504
rect 201370 448 204902 504
rect 204958 448 204963 504
rect 201309 446 204963 448
rect 201309 443 201375 446
rect 204897 443 204963 446
rect 205582 444 205588 508
rect 205652 506 205658 508
rect 206001 506 206067 509
rect 205652 504 206067 506
rect 205652 448 206006 504
rect 206062 448 206067 504
rect 205652 446 206067 448
rect 205652 444 205658 446
rect 206001 443 206067 446
rect 206921 506 206987 509
rect 210785 506 210851 509
rect 206921 504 210851 506
rect 206921 448 206926 504
rect 206982 448 210790 504
rect 210846 448 210851 504
rect 206921 446 210851 448
rect 206921 443 206987 446
rect 210785 443 210851 446
rect 242249 506 242315 509
rect 247309 506 247375 509
rect 242249 504 247375 506
rect 242249 448 242254 504
rect 242310 448 247314 504
rect 247370 448 247375 504
rect 242249 446 247375 448
rect 242249 443 242315 446
rect 247309 443 247375 446
rect 250897 506 250963 509
rect 256650 506 256710 582
rect 257061 579 257127 582
rect 267273 642 267339 645
rect 273621 642 273687 645
rect 267273 640 273687 642
rect 267273 584 267278 640
rect 267334 584 273626 640
rect 273682 584 273687 640
rect 267273 582 273687 584
rect 267273 579 267339 582
rect 273621 579 273687 582
rect 275185 642 275251 645
rect 278589 642 278655 645
rect 285397 642 285463 645
rect 275185 640 278146 642
rect 275185 584 275190 640
rect 275246 584 278146 640
rect 275185 582 278146 584
rect 275185 579 275251 582
rect 250897 504 256710 506
rect 250897 448 250902 504
rect 250958 448 256710 504
rect 250897 446 256710 448
rect 269481 506 269547 509
rect 276197 506 276263 509
rect 269481 504 276263 506
rect 269481 448 269486 504
rect 269542 448 276202 504
rect 276258 448 276263 504
rect 269481 446 276263 448
rect 278086 506 278146 582
rect 278589 640 285463 642
rect 278589 584 278594 640
rect 278650 584 285402 640
rect 285458 584 285463 640
rect 278589 582 285463 584
rect 278589 579 278655 582
rect 285397 579 285463 582
rect 285673 642 285739 645
rect 287789 642 287855 645
rect 292573 642 292639 645
rect 285673 640 287855 642
rect 285673 584 285678 640
rect 285734 584 287794 640
rect 287850 584 287855 640
rect 285673 582 287855 584
rect 285673 579 285739 582
rect 287789 579 287855 582
rect 288758 640 292639 642
rect 288758 584 292578 640
rect 292634 584 292639 640
rect 288758 582 292639 584
rect 282085 506 282151 509
rect 278086 504 282151 506
rect 278086 448 282090 504
rect 282146 448 282151 504
rect 278086 446 282151 448
rect 250897 443 250963 446
rect 269481 443 269547 446
rect 276197 443 276263 446
rect 282085 443 282151 446
rect 285213 506 285279 509
rect 288758 506 288818 582
rect 292573 579 292639 582
rect 293861 642 293927 645
rect 294873 642 294939 645
rect 293861 640 294939 642
rect 293861 584 293866 640
rect 293922 584 294878 640
rect 294934 584 294939 640
rect 293861 582 294939 584
rect 293861 579 293927 582
rect 294873 579 294939 582
rect 295609 642 295675 645
rect 303153 642 303219 645
rect 295609 640 303219 642
rect 295609 584 295614 640
rect 295670 584 303158 640
rect 303214 584 303219 640
rect 295609 582 303219 584
rect 295609 579 295675 582
rect 303153 579 303219 582
rect 305821 642 305887 645
rect 313825 642 313891 645
rect 318517 642 318583 645
rect 305821 640 313891 642
rect 305821 584 305826 640
rect 305882 584 313830 640
rect 313886 584 313891 640
rect 305821 582 313891 584
rect 305821 579 305887 582
rect 313825 579 313891 582
rect 318382 640 318583 642
rect 318382 584 318522 640
rect 318578 584 318583 640
rect 318382 582 318583 584
rect 285213 504 288818 506
rect 285213 448 285218 504
rect 285274 448 288818 504
rect 285213 446 288818 448
rect 303797 506 303863 509
rect 306925 506 306991 509
rect 303797 504 306991 506
rect 303797 448 303802 504
rect 303858 448 306930 504
rect 306986 448 306991 504
rect 303797 446 306991 448
rect 285213 443 285279 446
rect 303797 443 303863 446
rect 306925 443 306991 446
rect 309961 506 310027 509
rect 318382 506 318442 582
rect 318517 579 318583 582
rect 318885 642 318951 645
rect 319713 642 319779 645
rect 318885 640 319779 642
rect 318885 584 318890 640
rect 318946 584 319718 640
rect 319774 584 319779 640
rect 318885 582 319779 584
rect 318885 579 318951 582
rect 319713 579 319779 582
rect 334893 642 334959 645
rect 344553 642 344619 645
rect 334893 640 344619 642
rect 334893 584 334898 640
rect 334954 584 344558 640
rect 344614 584 344619 640
rect 334893 582 344619 584
rect 334893 579 334959 582
rect 344553 579 344619 582
rect 344737 642 344803 645
rect 345749 642 345815 645
rect 344737 640 345815 642
rect 344737 584 344742 640
rect 344798 584 345754 640
rect 345810 584 345815 640
rect 344737 582 345815 584
rect 344737 579 344803 582
rect 345749 579 345815 582
rect 350165 642 350231 645
rect 352557 642 352623 645
rect 354029 642 354095 645
rect 359917 642 359983 645
rect 350165 640 350550 642
rect 350165 584 350170 640
rect 350226 584 350550 640
rect 350165 582 350550 584
rect 350165 579 350231 582
rect 309961 504 318442 506
rect 309961 448 309966 504
rect 310022 448 318442 504
rect 309961 446 318442 448
rect 338297 506 338363 509
rect 347865 506 347931 509
rect 338297 504 347931 506
rect 338297 448 338302 504
rect 338358 448 347870 504
rect 347926 448 347931 504
rect 338297 446 347931 448
rect 309961 443 310027 446
rect 338297 443 338363 446
rect 347865 443 347931 446
rect 348417 506 348483 509
rect 350257 506 350323 509
rect 348417 504 350323 506
rect 348417 448 348422 504
rect 348478 448 350262 504
rect 350318 448 350323 504
rect 348417 446 350323 448
rect 350490 506 350550 582
rect 352557 640 354095 642
rect 352557 584 352562 640
rect 352618 584 354034 640
rect 354090 584 354095 640
rect 352557 582 354095 584
rect 352557 579 352623 582
rect 354029 579 354095 582
rect 356010 640 359983 642
rect 356010 584 359922 640
rect 359978 584 359983 640
rect 356010 582 359983 584
rect 356010 506 356070 582
rect 359917 579 359983 582
rect 363781 642 363847 645
rect 370589 642 370655 645
rect 374085 642 374151 645
rect 363781 640 370655 642
rect 363781 584 363786 640
rect 363842 584 370594 640
rect 370650 584 370655 640
rect 363781 582 370655 584
rect 363781 579 363847 582
rect 370589 579 370655 582
rect 372570 640 374151 642
rect 372570 584 374090 640
rect 374146 584 374151 640
rect 372570 582 374151 584
rect 350490 446 356070 506
rect 363689 506 363755 509
rect 372570 506 372630 582
rect 374085 579 374151 582
rect 374269 642 374335 645
rect 375281 642 375347 645
rect 374269 640 375347 642
rect 374269 584 374274 640
rect 374330 584 375286 640
rect 375342 584 375347 640
rect 374269 582 375347 584
rect 374269 579 374335 582
rect 375281 579 375347 582
rect 375465 642 375531 645
rect 378869 642 378935 645
rect 375465 640 378935 642
rect 375465 584 375470 640
rect 375526 584 378874 640
rect 378930 584 378935 640
rect 375465 582 378935 584
rect 375465 579 375531 582
rect 378869 579 378935 582
rect 379053 642 379119 645
rect 381169 642 381235 645
rect 383561 642 383627 645
rect 379053 640 381235 642
rect 379053 584 379058 640
rect 379114 584 381174 640
rect 381230 584 381235 640
rect 379053 582 381235 584
rect 379053 579 379119 582
rect 381169 579 381235 582
rect 382230 640 383627 642
rect 382230 584 383566 640
rect 383622 584 383627 640
rect 382230 582 383627 584
rect 363689 504 372630 506
rect 363689 448 363694 504
rect 363750 448 372630 504
rect 363689 446 372630 448
rect 374361 506 374427 509
rect 377489 506 377555 509
rect 374361 504 377555 506
rect 374361 448 374366 504
rect 374422 448 377494 504
rect 377550 448 377555 504
rect 374361 446 377555 448
rect 348417 443 348483 446
rect 350257 443 350323 446
rect 363689 443 363755 446
rect 374361 443 374427 446
rect 377489 443 377555 446
rect 379605 506 379671 509
rect 382230 506 382290 582
rect 383561 579 383627 582
rect 391013 642 391079 645
rect 402513 642 402579 645
rect 391013 640 402579 642
rect 391013 584 391018 640
rect 391074 584 402518 640
rect 402574 584 402579 640
rect 391013 582 402579 584
rect 391013 579 391079 582
rect 402513 579 402579 582
rect 403065 642 403131 645
rect 403617 642 403683 645
rect 403065 640 403683 642
rect 403065 584 403070 640
rect 403126 584 403622 640
rect 403678 584 403683 640
rect 403065 582 403683 584
rect 403065 579 403131 582
rect 403617 579 403683 582
rect 405641 642 405707 645
rect 408401 642 408467 645
rect 409597 642 409663 645
rect 405641 640 408467 642
rect 405641 584 405646 640
rect 405702 584 408406 640
rect 408462 584 408467 640
rect 405641 582 408467 584
rect 405641 579 405707 582
rect 408401 579 408467 582
rect 409462 640 409663 642
rect 409462 584 409602 640
rect 409658 584 409663 640
rect 409462 582 409663 584
rect 379605 504 382290 506
rect 379605 448 379610 504
rect 379666 448 382290 504
rect 379605 446 382290 448
rect 384205 506 384271 509
rect 395521 506 395587 509
rect 384205 504 395587 506
rect 384205 448 384210 504
rect 384266 448 395526 504
rect 395582 448 395587 504
rect 384205 446 395587 448
rect 379605 443 379671 446
rect 384205 443 384271 446
rect 395521 443 395587 446
rect 407481 506 407547 509
rect 409462 506 409522 582
rect 409597 579 409663 582
rect 421005 642 421071 645
rect 423765 642 423831 645
rect 424961 642 425027 645
rect 421005 640 423831 642
rect 421005 584 421010 640
rect 421066 584 423770 640
rect 423826 584 423831 640
rect 421005 582 423831 584
rect 421005 579 421071 582
rect 423765 579 423831 582
rect 424918 640 425027 642
rect 424918 584 424966 640
rect 425022 584 425027 640
rect 424918 579 425027 584
rect 427905 642 427971 645
rect 429653 642 429719 645
rect 427905 640 429719 642
rect 427905 584 427910 640
rect 427966 584 429658 640
rect 429714 584 429719 640
rect 427905 582 429719 584
rect 427905 579 427971 582
rect 429653 579 429719 582
rect 431033 642 431099 645
rect 432045 642 432111 645
rect 431033 640 432111 642
rect 431033 584 431038 640
rect 431094 584 432050 640
rect 432106 584 432111 640
rect 431033 582 432111 584
rect 431033 579 431099 582
rect 432045 579 432111 582
rect 456057 642 456123 645
rect 460381 642 460447 645
rect 456057 640 460447 642
rect 456057 584 456062 640
rect 456118 584 460386 640
rect 460442 584 460447 640
rect 456057 582 460447 584
rect 456057 579 456123 582
rect 460381 579 460447 582
rect 460933 642 460999 645
rect 462773 642 462839 645
rect 463969 642 464035 645
rect 460933 640 462839 642
rect 460933 584 460938 640
rect 460994 584 462778 640
rect 462834 584 462839 640
rect 460933 582 462839 584
rect 460933 579 460999 582
rect 462773 579 462839 582
rect 463926 640 464035 642
rect 463926 584 463974 640
rect 464030 584 464035 640
rect 463926 579 464035 584
rect 480805 642 480871 645
rect 481725 642 481791 645
rect 480805 640 481791 642
rect 480805 584 480810 640
rect 480866 584 481730 640
rect 481786 584 481791 640
rect 480805 582 481791 584
rect 480805 579 480871 582
rect 481725 579 481791 582
rect 483565 642 483631 645
rect 488809 642 488875 645
rect 492305 642 492371 645
rect 483565 640 488875 642
rect 483565 584 483570 640
rect 483626 584 488814 640
rect 488870 584 488875 640
rect 483565 582 488875 584
rect 483565 579 483631 582
rect 488809 579 488875 582
rect 488950 640 492371 642
rect 488950 584 492310 640
rect 492366 584 492371 640
rect 488950 582 492371 584
rect 407481 504 409522 506
rect 407481 448 407486 504
rect 407542 448 409522 504
rect 407481 446 409522 448
rect 418613 506 418679 509
rect 424918 506 424978 579
rect 418613 504 424978 506
rect 418613 448 418618 504
rect 418674 448 424978 504
rect 418613 446 424978 448
rect 453481 506 453547 509
rect 461761 506 461827 509
rect 453481 504 461827 506
rect 453481 448 453486 504
rect 453542 448 461766 504
rect 461822 448 461827 504
rect 453481 446 461827 448
rect 407481 443 407547 446
rect 418613 443 418679 446
rect 453481 443 453547 446
rect 461761 443 461827 446
rect 461945 506 462011 509
rect 463926 506 463986 579
rect 461945 504 463986 506
rect 461945 448 461950 504
rect 462006 448 463986 504
rect 461945 446 463986 448
rect 477401 506 477467 509
rect 488950 506 489010 582
rect 492305 579 492371 582
rect 492673 642 492739 645
rect 495893 642 495959 645
rect 492673 640 495959 642
rect 492673 584 492678 640
rect 492734 584 495898 640
rect 495954 584 495959 640
rect 498101 642 498167 645
rect 500585 642 500651 645
rect 498101 640 500651 642
rect 497089 608 497155 611
rect 492673 582 495959 584
rect 492673 579 492739 582
rect 495893 579 495959 582
rect 497046 606 497155 608
rect 497046 550 497094 606
rect 497150 550 497155 606
rect 498101 584 498106 640
rect 498162 584 500590 640
rect 500646 584 500651 640
rect 498101 582 500651 584
rect 498101 579 498167 582
rect 500585 579 500651 582
rect 509877 642 509943 645
rect 512453 642 512519 645
rect 509877 640 512519 642
rect 509877 584 509882 640
rect 509938 584 512458 640
rect 512514 584 512519 640
rect 509877 582 512519 584
rect 509877 579 509943 582
rect 512453 579 512519 582
rect 514661 640 514770 645
rect 514661 584 514666 640
rect 514722 584 514770 640
rect 514661 582 514770 584
rect 515397 642 515463 645
rect 515949 642 516015 645
rect 515397 640 516015 642
rect 515397 584 515402 640
rect 515458 584 515954 640
rect 516010 584 516015 640
rect 515397 582 516015 584
rect 514661 579 514727 582
rect 515397 579 515463 582
rect 515949 579 516015 582
rect 523217 642 523283 645
rect 525425 642 525491 645
rect 523217 640 525491 642
rect 523217 584 523222 640
rect 523278 584 525430 640
rect 525486 584 525491 640
rect 523217 582 525491 584
rect 523217 579 523283 582
rect 525425 579 525491 582
rect 527173 642 527239 645
rect 532006 642 532066 854
rect 542486 852 542492 854
rect 542556 852 542562 916
rect 551134 778 551140 780
rect 535410 718 551140 778
rect 527173 640 532066 642
rect 527173 584 527178 640
rect 527234 584 532066 640
rect 527173 582 532066 584
rect 534165 642 534231 645
rect 535410 642 535470 718
rect 551134 716 551140 718
rect 551204 716 551210 780
rect 553350 778 553410 1126
rect 553350 718 560770 778
rect 534165 640 535470 642
rect 534165 584 534170 640
rect 534226 584 535470 640
rect 534165 582 535470 584
rect 540513 642 540579 645
rect 558545 642 558611 645
rect 540513 640 558611 642
rect 540513 584 540518 640
rect 540574 584 558550 640
rect 558606 584 558611 640
rect 540513 582 558611 584
rect 560710 642 560770 718
rect 560845 642 560911 645
rect 560710 640 560911 642
rect 560710 584 560850 640
rect 560906 584 560911 640
rect 560710 582 560911 584
rect 527173 579 527239 582
rect 534165 579 534231 582
rect 540513 579 540579 582
rect 558545 579 558611 582
rect 560845 579 560911 582
rect 497046 545 497155 550
rect 477401 504 489010 506
rect 477401 448 477406 504
rect 477462 448 489010 504
rect 477401 446 489010 448
rect 492673 506 492739 509
rect 497046 506 497106 545
rect 492673 504 497106 506
rect 492673 448 492678 504
rect 492734 448 497106 504
rect 492673 446 497106 448
rect 523309 506 523375 509
rect 527633 506 527699 509
rect 523309 504 527699 506
rect 523309 448 523314 504
rect 523370 448 527638 504
rect 527694 448 527699 504
rect 523309 446 527699 448
rect 461945 443 462011 446
rect 477401 443 477467 446
rect 492673 443 492739 446
rect 523309 443 523375 446
rect 527633 443 527699 446
rect 528461 506 528527 509
rect 534165 506 534231 509
rect 528461 504 534231 506
rect 528461 448 528466 504
rect 528522 448 534170 504
rect 534226 448 534231 504
rect 528461 446 534231 448
rect 528461 443 528527 446
rect 534165 443 534231 446
rect 536465 506 536531 509
rect 540973 506 541039 509
rect 536465 504 541039 506
rect 536465 448 536470 504
rect 536526 448 540978 504
rect 541034 448 541039 504
rect 536465 446 541039 448
rect 536465 443 536531 446
rect 540973 443 541039 446
rect 542486 444 542492 508
rect 542556 506 542562 508
rect 542629 506 542695 509
rect 542813 508 542879 509
rect 542813 506 542860 508
rect 542556 504 542695 506
rect 542556 448 542634 504
rect 542690 448 542695 504
rect 542556 446 542695 448
rect 542768 504 542860 506
rect 542768 448 542818 504
rect 542768 446 542860 448
rect 542556 444 542562 446
rect 542629 443 542695 446
rect 542813 444 542860 446
rect 542924 444 542930 508
rect 543457 506 543523 509
rect 554773 506 554839 509
rect 543457 504 554839 506
rect 543457 448 543462 504
rect 543518 448 554778 504
rect 554834 448 554839 504
rect 543457 446 554839 448
rect 542813 443 542879 444
rect 543457 443 543523 446
rect 554773 443 554839 446
rect 202505 370 202571 373
rect 200806 368 202571 370
rect 200806 312 202510 368
rect 202566 312 202571 368
rect 200806 310 202571 312
rect 196617 307 196683 310
rect 200113 307 200179 310
rect 202505 307 202571 310
rect 204805 370 204871 373
rect 208761 370 208827 373
rect 204805 368 208827 370
rect 204805 312 204810 368
rect 204866 312 208766 368
rect 208822 312 208827 368
rect 204805 310 208827 312
rect 204805 307 204871 310
rect 208761 307 208827 310
rect 286409 370 286475 373
rect 293401 370 293467 373
rect 286409 368 293467 370
rect 286409 312 286414 368
rect 286470 312 293406 368
rect 293462 312 293467 368
rect 286409 310 293467 312
rect 286409 307 286475 310
rect 293401 307 293467 310
rect 364977 370 365043 373
rect 373073 370 373139 373
rect 364977 368 373139 370
rect 364977 312 364982 368
rect 365038 312 373078 368
rect 373134 312 373139 368
rect 364977 310 373139 312
rect 364977 307 365043 310
rect 373073 307 373139 310
rect 530761 370 530827 373
rect 548057 370 548123 373
rect 551185 372 551251 373
rect 530761 368 548123 370
rect 530761 312 530766 368
rect 530822 312 548062 368
rect 548118 312 548123 368
rect 530761 310 548123 312
rect 530761 307 530827 310
rect 548057 307 548123 310
rect 551134 308 551140 372
rect 551204 370 551251 372
rect 551204 368 551296 370
rect 551246 312 551296 368
rect 551204 310 551296 312
rect 551204 308 551251 310
rect 551185 307 551251 308
rect 202413 234 202479 237
rect 205582 234 205588 236
rect 202413 232 205588 234
rect 202413 176 202418 232
rect 202474 176 205588 232
rect 202413 174 205588 176
rect 202413 171 202479 174
rect 205582 172 205588 174
rect 205652 172 205658 236
rect 328453 234 328519 237
rect 336641 234 336707 237
rect 328453 232 336707 234
rect 328453 176 328458 232
rect 328514 176 336646 232
rect 336702 176 336707 232
rect 328453 174 336707 176
rect 328453 171 328519 174
rect 336641 171 336707 174
rect 349429 234 349495 237
rect 351453 234 351519 237
rect 349429 232 351519 234
rect 349429 176 349434 232
rect 349490 176 351458 232
rect 351514 176 351519 232
rect 349429 174 351519 176
rect 349429 171 349495 174
rect 351453 171 351519 174
rect 381997 234 382063 237
rect 384573 234 384639 237
rect 531129 236 531195 237
rect 381997 232 384639 234
rect 381997 176 382002 232
rect 382058 176 384578 232
rect 384634 176 384639 232
rect 381997 174 384639 176
rect 381997 171 382063 174
rect 384573 171 384639 174
rect 531078 172 531084 236
rect 531148 234 531195 236
rect 541709 234 541775 237
rect 559557 234 559623 237
rect 531148 232 531240 234
rect 531190 176 531240 232
rect 531148 174 531240 176
rect 541709 232 559623 234
rect 541709 176 541714 232
rect 541770 176 559562 232
rect 559618 176 559623 232
rect 541709 174 559623 176
rect 531148 172 531195 174
rect 531129 171 531195 172
rect 541709 171 541775 174
rect 559557 171 559623 174
rect 197721 98 197787 101
rect 201677 98 201743 101
rect 197721 96 201743 98
rect 197721 40 197726 96
rect 197782 40 201682 96
rect 201738 40 201743 96
rect 197721 38 201743 40
rect 197721 35 197787 38
rect 201677 35 201743 38
rect 376753 98 376819 101
rect 379789 98 379855 101
rect 376753 96 379855 98
rect 376753 40 376758 96
rect 376814 40 379794 96
rect 379850 40 379855 96
rect 376753 38 379855 40
rect 376753 35 376819 38
rect 379789 35 379855 38
<< via3 >>
rect 453988 701932 454052 701996
rect 259132 701660 259196 701724
rect 453988 699544 454052 699548
rect 453988 699488 454002 699544
rect 454002 699488 454052 699544
rect 453988 699484 454052 699488
rect 13860 699348 13924 699412
rect 43116 699348 43180 699412
rect 52868 699348 52932 699412
rect 60228 699348 60292 699412
rect 124628 699408 124692 699412
rect 124628 699352 124642 699408
rect 124642 699352 124692 699408
rect 124628 699348 124692 699352
rect 124444 699076 124508 699140
rect 418660 699408 418724 699412
rect 418660 699352 418710 699408
rect 418710 699352 418724 699408
rect 418660 699348 418724 699352
rect 433380 699408 433444 699412
rect 433380 699352 433430 699408
rect 433430 699352 433444 699408
rect 433380 699348 433444 699352
rect 462820 699408 462884 699412
rect 462820 699352 462870 699408
rect 462870 699352 462884 699408
rect 462820 699348 462884 699352
rect 492628 699408 492692 699412
rect 492628 699352 492642 699408
rect 492642 699352 492692 699408
rect 492628 699348 492692 699352
rect 510660 699348 510724 699412
rect 539916 699348 539980 699412
rect 259132 699076 259196 699140
rect 510660 698940 510724 699004
rect 60228 698804 60292 698868
rect 52868 698668 52932 698732
rect 43116 698532 43180 698596
rect 539916 698396 539980 698460
rect 13860 698260 13924 698324
rect 418660 698124 418724 698188
rect 433380 697988 433444 698052
rect 124444 697852 124508 697916
rect 124628 697852 124692 697916
rect 462820 697716 462884 697780
rect 492628 697580 492692 697644
rect 531084 1396 531148 1460
rect 542860 1124 542924 1188
rect 205588 444 205652 508
rect 542492 852 542556 916
rect 551140 716 551204 780
rect 542492 444 542556 508
rect 542860 504 542924 508
rect 542860 448 542874 504
rect 542874 448 542924 504
rect 542860 444 542924 448
rect 551140 368 551204 372
rect 551140 312 551190 368
rect 551190 312 551204 368
rect 551140 308 551204 312
rect 205588 172 205652 236
rect 531084 232 531148 236
rect 531084 176 531134 232
rect 531134 176 531148 232
rect 531084 172 531148 176
<< metal4 >>
rect -8726 711558 -8106 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 -8106 711558
rect -8726 711238 -8106 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 -8106 711238
rect -8726 680614 -8106 711002
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 -8106 680614
rect -8726 680294 -8106 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 -8106 680294
rect -8726 644614 -8106 680058
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 -8106 644614
rect -8726 644294 -8106 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 -8106 644294
rect -8726 608614 -8106 644058
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 -8106 608614
rect -8726 608294 -8106 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 -8106 608294
rect -8726 572614 -8106 608058
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 -8106 572614
rect -8726 572294 -8106 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 -8106 572294
rect -8726 536614 -8106 572058
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 -8106 536614
rect -8726 536294 -8106 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 -8106 536294
rect -8726 500614 -8106 536058
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 -8106 500614
rect -8726 500294 -8106 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 -8106 500294
rect -8726 464614 -8106 500058
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 -8106 464614
rect -8726 464294 -8106 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 -8106 464294
rect -8726 428614 -8106 464058
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 -8106 428614
rect -8726 428294 -8106 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 -8106 428294
rect -8726 392614 -8106 428058
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 -8106 392614
rect -8726 392294 -8106 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 -8106 392294
rect -8726 356614 -8106 392058
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 -8106 356614
rect -8726 356294 -8106 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 -8106 356294
rect -8726 320614 -8106 356058
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 -8106 320614
rect -8726 320294 -8106 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 -8106 320294
rect -8726 284614 -8106 320058
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 -8106 284614
rect -8726 284294 -8106 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 -8106 284294
rect -8726 248614 -8106 284058
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 -8106 248614
rect -8726 248294 -8106 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 -8106 248294
rect -8726 212614 -8106 248058
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 -8106 212614
rect -8726 212294 -8106 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 -8106 212294
rect -8726 176614 -8106 212058
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 -8106 176614
rect -8726 176294 -8106 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 -8106 176294
rect -8726 140614 -8106 176058
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 -8106 140614
rect -8726 140294 -8106 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 -8106 140294
rect -8726 104614 -8106 140058
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 -8106 104614
rect -8726 104294 -8106 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 -8106 104294
rect -8726 68614 -8106 104058
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 -8106 68614
rect -8726 68294 -8106 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 -8106 68294
rect -8726 32614 -8106 68058
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 -8106 32614
rect -8726 32294 -8106 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 -8106 32294
rect -8726 -7066 -8106 32058
rect -7766 710598 -7146 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 -7146 710598
rect -7766 710278 -7146 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 -7146 710278
rect -7766 698614 -7146 710042
rect 12954 710598 13574 711590
rect 12954 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 13574 710598
rect 12954 710278 13574 710362
rect 12954 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 13574 710278
rect -7766 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 -7146 698614
rect -7766 698294 -7146 698378
rect -7766 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 -7146 698294
rect -7766 662614 -7146 698058
rect -7766 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 -7146 662614
rect -7766 662294 -7146 662378
rect -7766 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 -7146 662294
rect -7766 626614 -7146 662058
rect -7766 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 -7146 626614
rect -7766 626294 -7146 626378
rect -7766 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 -7146 626294
rect -7766 590614 -7146 626058
rect -7766 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 -7146 590614
rect -7766 590294 -7146 590378
rect -7766 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 -7146 590294
rect -7766 554614 -7146 590058
rect -7766 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 -7146 554614
rect -7766 554294 -7146 554378
rect -7766 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 -7146 554294
rect -7766 518614 -7146 554058
rect -7766 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 -7146 518614
rect -7766 518294 -7146 518378
rect -7766 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 -7146 518294
rect -7766 482614 -7146 518058
rect -7766 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 -7146 482614
rect -7766 482294 -7146 482378
rect -7766 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 -7146 482294
rect -7766 446614 -7146 482058
rect -7766 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 -7146 446614
rect -7766 446294 -7146 446378
rect -7766 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 -7146 446294
rect -7766 410614 -7146 446058
rect -7766 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 -7146 410614
rect -7766 410294 -7146 410378
rect -7766 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 -7146 410294
rect -7766 374614 -7146 410058
rect -7766 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 -7146 374614
rect -7766 374294 -7146 374378
rect -7766 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 -7146 374294
rect -7766 338614 -7146 374058
rect -7766 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 -7146 338614
rect -7766 338294 -7146 338378
rect -7766 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 -7146 338294
rect -7766 302614 -7146 338058
rect -7766 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 -7146 302614
rect -7766 302294 -7146 302378
rect -7766 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 -7146 302294
rect -7766 266614 -7146 302058
rect -7766 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 -7146 266614
rect -7766 266294 -7146 266378
rect -7766 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 -7146 266294
rect -7766 230614 -7146 266058
rect -7766 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 -7146 230614
rect -7766 230294 -7146 230378
rect -7766 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 -7146 230294
rect -7766 194614 -7146 230058
rect -7766 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 -7146 194614
rect -7766 194294 -7146 194378
rect -7766 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 -7146 194294
rect -7766 158614 -7146 194058
rect -7766 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 -7146 158614
rect -7766 158294 -7146 158378
rect -7766 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 -7146 158294
rect -7766 122614 -7146 158058
rect -7766 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 -7146 122614
rect -7766 122294 -7146 122378
rect -7766 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 -7146 122294
rect -7766 86614 -7146 122058
rect -7766 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 -7146 86614
rect -7766 86294 -7146 86378
rect -7766 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 -7146 86294
rect -7766 50614 -7146 86058
rect -7766 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 -7146 50614
rect -7766 50294 -7146 50378
rect -7766 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 -7146 50294
rect -7766 14614 -7146 50058
rect -7766 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 -7146 14614
rect -7766 14294 -7146 14378
rect -7766 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 -7146 14294
rect -7766 -6106 -7146 14058
rect -6806 709638 -6186 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 -6186 709638
rect -6806 709318 -6186 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 -6186 709318
rect -6806 676894 -6186 709082
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 -6186 676894
rect -6806 676574 -6186 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 -6186 676574
rect -6806 640894 -6186 676338
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 -6186 640894
rect -6806 640574 -6186 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 -6186 640574
rect -6806 604894 -6186 640338
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 -6186 604894
rect -6806 604574 -6186 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 -6186 604574
rect -6806 568894 -6186 604338
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 -6186 568894
rect -6806 568574 -6186 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 -6186 568574
rect -6806 532894 -6186 568338
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 -6186 532894
rect -6806 532574 -6186 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 -6186 532574
rect -6806 496894 -6186 532338
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 -6186 496894
rect -6806 496574 -6186 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 -6186 496574
rect -6806 460894 -6186 496338
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 -6186 460894
rect -6806 460574 -6186 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 -6186 460574
rect -6806 424894 -6186 460338
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 -6186 424894
rect -6806 424574 -6186 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 -6186 424574
rect -6806 388894 -6186 424338
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 -6186 388894
rect -6806 388574 -6186 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 -6186 388574
rect -6806 352894 -6186 388338
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 -6186 352894
rect -6806 352574 -6186 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 -6186 352574
rect -6806 316894 -6186 352338
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 -6186 316894
rect -6806 316574 -6186 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 -6186 316574
rect -6806 280894 -6186 316338
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 -6186 280894
rect -6806 280574 -6186 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 -6186 280574
rect -6806 244894 -6186 280338
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 -6186 244894
rect -6806 244574 -6186 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 -6186 244574
rect -6806 208894 -6186 244338
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 -6186 208894
rect -6806 208574 -6186 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 -6186 208574
rect -6806 172894 -6186 208338
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 -6186 172894
rect -6806 172574 -6186 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 -6186 172574
rect -6806 136894 -6186 172338
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 -6186 136894
rect -6806 136574 -6186 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 -6186 136574
rect -6806 100894 -6186 136338
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 -6186 100894
rect -6806 100574 -6186 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 -6186 100574
rect -6806 64894 -6186 100338
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 -6186 64894
rect -6806 64574 -6186 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 -6186 64574
rect -6806 28894 -6186 64338
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 -6186 28894
rect -6806 28574 -6186 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 -6186 28574
rect -6806 -5146 -6186 28338
rect -5846 708678 -5226 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 -5226 708678
rect -5846 708358 -5226 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 -5226 708358
rect -5846 694894 -5226 708122
rect 9234 708678 9854 709670
rect 9234 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 9854 708678
rect 9234 708358 9854 708442
rect 9234 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 9854 708358
rect -5846 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 -5226 694894
rect -5846 694574 -5226 694658
rect -5846 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 -5226 694574
rect -5846 658894 -5226 694338
rect -5846 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 -5226 658894
rect -5846 658574 -5226 658658
rect -5846 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 -5226 658574
rect -5846 622894 -5226 658338
rect -5846 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 -5226 622894
rect -5846 622574 -5226 622658
rect -5846 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 -5226 622574
rect -5846 586894 -5226 622338
rect -5846 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 -5226 586894
rect -5846 586574 -5226 586658
rect -5846 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 -5226 586574
rect -5846 550894 -5226 586338
rect -5846 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 -5226 550894
rect -5846 550574 -5226 550658
rect -5846 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 -5226 550574
rect -5846 514894 -5226 550338
rect -5846 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 -5226 514894
rect -5846 514574 -5226 514658
rect -5846 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 -5226 514574
rect -5846 478894 -5226 514338
rect -5846 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 -5226 478894
rect -5846 478574 -5226 478658
rect -5846 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 -5226 478574
rect -5846 442894 -5226 478338
rect -5846 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 -5226 442894
rect -5846 442574 -5226 442658
rect -5846 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 -5226 442574
rect -5846 406894 -5226 442338
rect -5846 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 -5226 406894
rect -5846 406574 -5226 406658
rect -5846 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 -5226 406574
rect -5846 370894 -5226 406338
rect -5846 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 -5226 370894
rect -5846 370574 -5226 370658
rect -5846 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 -5226 370574
rect -5846 334894 -5226 370338
rect -5846 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 -5226 334894
rect -5846 334574 -5226 334658
rect -5846 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 -5226 334574
rect -5846 298894 -5226 334338
rect -5846 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 -5226 298894
rect -5846 298574 -5226 298658
rect -5846 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 -5226 298574
rect -5846 262894 -5226 298338
rect -5846 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 -5226 262894
rect -5846 262574 -5226 262658
rect -5846 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 -5226 262574
rect -5846 226894 -5226 262338
rect -5846 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 -5226 226894
rect -5846 226574 -5226 226658
rect -5846 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 -5226 226574
rect -5846 190894 -5226 226338
rect -5846 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 -5226 190894
rect -5846 190574 -5226 190658
rect -5846 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 -5226 190574
rect -5846 154894 -5226 190338
rect -5846 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 -5226 154894
rect -5846 154574 -5226 154658
rect -5846 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 -5226 154574
rect -5846 118894 -5226 154338
rect -5846 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 -5226 118894
rect -5846 118574 -5226 118658
rect -5846 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 -5226 118574
rect -5846 82894 -5226 118338
rect -5846 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 -5226 82894
rect -5846 82574 -5226 82658
rect -5846 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 -5226 82574
rect -5846 46894 -5226 82338
rect -5846 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 -5226 46894
rect -5846 46574 -5226 46658
rect -5846 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 -5226 46574
rect -5846 10894 -5226 46338
rect -5846 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 -5226 10894
rect -5846 10574 -5226 10658
rect -5846 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 -5226 10574
rect -5846 -4186 -5226 10338
rect -4886 707718 -4266 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 -4266 707718
rect -4886 707398 -4266 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 -4266 707398
rect -4886 673174 -4266 707162
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 -4266 673174
rect -4886 672854 -4266 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 -4266 672854
rect -4886 637174 -4266 672618
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 -4266 637174
rect -4886 636854 -4266 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 -4266 636854
rect -4886 601174 -4266 636618
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 -4266 601174
rect -4886 600854 -4266 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 -4266 600854
rect -4886 565174 -4266 600618
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 -4266 565174
rect -4886 564854 -4266 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 -4266 564854
rect -4886 529174 -4266 564618
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 -4266 529174
rect -4886 528854 -4266 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 -4266 528854
rect -4886 493174 -4266 528618
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 -4266 493174
rect -4886 492854 -4266 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 -4266 492854
rect -4886 457174 -4266 492618
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 -4266 457174
rect -4886 456854 -4266 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 -4266 456854
rect -4886 421174 -4266 456618
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 -4266 421174
rect -4886 420854 -4266 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 -4266 420854
rect -4886 385174 -4266 420618
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 -4266 385174
rect -4886 384854 -4266 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 -4266 384854
rect -4886 349174 -4266 384618
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 -4266 349174
rect -4886 348854 -4266 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 -4266 348854
rect -4886 313174 -4266 348618
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 -4266 313174
rect -4886 312854 -4266 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 -4266 312854
rect -4886 277174 -4266 312618
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 -4266 277174
rect -4886 276854 -4266 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 -4266 276854
rect -4886 241174 -4266 276618
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 -4266 241174
rect -4886 240854 -4266 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 -4266 240854
rect -4886 205174 -4266 240618
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 -4266 205174
rect -4886 204854 -4266 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 -4266 204854
rect -4886 169174 -4266 204618
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 -4266 169174
rect -4886 168854 -4266 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 -4266 168854
rect -4886 133174 -4266 168618
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 -4266 133174
rect -4886 132854 -4266 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 -4266 132854
rect -4886 97174 -4266 132618
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 -4266 97174
rect -4886 96854 -4266 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 -4266 96854
rect -4886 61174 -4266 96618
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 -4266 61174
rect -4886 60854 -4266 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 -4266 60854
rect -4886 25174 -4266 60618
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 -4266 25174
rect -4886 24854 -4266 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 -4266 24854
rect -4886 -3226 -4266 24618
rect -3926 706758 -3306 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 -3306 706758
rect -3926 706438 -3306 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 -3306 706438
rect -3926 691174 -3306 706202
rect 5514 706758 6134 707750
rect 5514 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 6134 706758
rect 5514 706438 6134 706522
rect 5514 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 6134 706438
rect -3926 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 -3306 691174
rect -3926 690854 -3306 690938
rect -3926 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 -3306 690854
rect -3926 655174 -3306 690618
rect -3926 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 -3306 655174
rect -3926 654854 -3306 654938
rect -3926 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 -3306 654854
rect -3926 619174 -3306 654618
rect -3926 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 -3306 619174
rect -3926 618854 -3306 618938
rect -3926 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 -3306 618854
rect -3926 583174 -3306 618618
rect -3926 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 -3306 583174
rect -3926 582854 -3306 582938
rect -3926 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 -3306 582854
rect -3926 547174 -3306 582618
rect -3926 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 -3306 547174
rect -3926 546854 -3306 546938
rect -3926 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 -3306 546854
rect -3926 511174 -3306 546618
rect -3926 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 -3306 511174
rect -3926 510854 -3306 510938
rect -3926 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 -3306 510854
rect -3926 475174 -3306 510618
rect -3926 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 -3306 475174
rect -3926 474854 -3306 474938
rect -3926 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 -3306 474854
rect -3926 439174 -3306 474618
rect -3926 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 -3306 439174
rect -3926 438854 -3306 438938
rect -3926 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 -3306 438854
rect -3926 403174 -3306 438618
rect -3926 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 -3306 403174
rect -3926 402854 -3306 402938
rect -3926 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 -3306 402854
rect -3926 367174 -3306 402618
rect -3926 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 -3306 367174
rect -3926 366854 -3306 366938
rect -3926 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 -3306 366854
rect -3926 331174 -3306 366618
rect -3926 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 -3306 331174
rect -3926 330854 -3306 330938
rect -3926 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 -3306 330854
rect -3926 295174 -3306 330618
rect -3926 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 -3306 295174
rect -3926 294854 -3306 294938
rect -3926 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 -3306 294854
rect -3926 259174 -3306 294618
rect -3926 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 -3306 259174
rect -3926 258854 -3306 258938
rect -3926 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 -3306 258854
rect -3926 223174 -3306 258618
rect -3926 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 -3306 223174
rect -3926 222854 -3306 222938
rect -3926 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 -3306 222854
rect -3926 187174 -3306 222618
rect -3926 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 -3306 187174
rect -3926 186854 -3306 186938
rect -3926 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 -3306 186854
rect -3926 151174 -3306 186618
rect -3926 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 -3306 151174
rect -3926 150854 -3306 150938
rect -3926 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 -3306 150854
rect -3926 115174 -3306 150618
rect -3926 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 -3306 115174
rect -3926 114854 -3306 114938
rect -3926 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 -3306 114854
rect -3926 79174 -3306 114618
rect -3926 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 -3306 79174
rect -3926 78854 -3306 78938
rect -3926 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 -3306 78854
rect -3926 43174 -3306 78618
rect -3926 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 -3306 43174
rect -3926 42854 -3306 42938
rect -3926 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 -3306 42854
rect -3926 7174 -3306 42618
rect -3926 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 -3306 7174
rect -3926 6854 -3306 6938
rect -3926 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 -3306 6854
rect -3926 -2266 -3306 6618
rect -2966 705798 -2346 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 -2346 705798
rect -2966 705478 -2346 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 -2346 705478
rect -2966 669454 -2346 705242
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 -2346 669454
rect -2966 669134 -2346 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 -2346 669134
rect -2966 633454 -2346 668898
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 -2346 633454
rect -2966 633134 -2346 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 -2346 633134
rect -2966 597454 -2346 632898
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 -2346 597454
rect -2966 597134 -2346 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 -2346 597134
rect -2966 561454 -2346 596898
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 -2346 561454
rect -2966 561134 -2346 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 -2346 561134
rect -2966 525454 -2346 560898
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 -2346 525454
rect -2966 525134 -2346 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 -2346 525134
rect -2966 489454 -2346 524898
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 -2346 489454
rect -2966 489134 -2346 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 -2346 489134
rect -2966 453454 -2346 488898
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 -2346 453454
rect -2966 453134 -2346 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 -2346 453134
rect -2966 417454 -2346 452898
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 -2346 417454
rect -2966 417134 -2346 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 -2346 417134
rect -2966 381454 -2346 416898
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 -2346 381454
rect -2966 381134 -2346 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 -2346 381134
rect -2966 345454 -2346 380898
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 -2346 345454
rect -2966 345134 -2346 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 -2346 345134
rect -2966 309454 -2346 344898
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 -2346 309454
rect -2966 309134 -2346 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 -2346 309134
rect -2966 273454 -2346 308898
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 -2346 273454
rect -2966 273134 -2346 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 -2346 273134
rect -2966 237454 -2346 272898
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 -2346 237454
rect -2966 237134 -2346 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 -2346 237134
rect -2966 201454 -2346 236898
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 -2346 201454
rect -2966 201134 -2346 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 -2346 201134
rect -2966 165454 -2346 200898
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 -2346 165454
rect -2966 165134 -2346 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 -2346 165134
rect -2966 129454 -2346 164898
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 -2346 129454
rect -2966 129134 -2346 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 -2346 129134
rect -2966 93454 -2346 128898
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 -2346 93454
rect -2966 93134 -2346 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 -2346 93134
rect -2966 57454 -2346 92898
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 -2346 57454
rect -2966 57134 -2346 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 -2346 57134
rect -2966 21454 -2346 56898
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 -2346 21454
rect -2966 21134 -2346 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 -2346 21134
rect -2966 -1306 -2346 20898
rect -2006 704838 -1386 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 -1386 704838
rect -2006 704518 -1386 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 -1386 704518
rect -2006 687454 -1386 704282
rect 1794 704838 2414 705830
rect 1794 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 2414 704838
rect 1794 704518 2414 704602
rect 1794 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 2414 704518
rect 1794 702000 2414 704282
rect 5514 702000 6134 706202
rect 9234 702000 9854 708122
rect 12954 702000 13574 710042
rect 30954 711558 31574 711590
rect 30954 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 31574 711558
rect 30954 711238 31574 711322
rect 30954 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 31574 711238
rect 27234 709638 27854 709670
rect 27234 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 27854 709638
rect 27234 709318 27854 709402
rect 27234 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 27854 709318
rect 23514 707718 24134 707750
rect 23514 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 24134 707718
rect 23514 707398 24134 707482
rect 23514 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 24134 707398
rect 19794 705798 20414 705830
rect 19794 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 20414 705798
rect 19794 705478 20414 705562
rect 19794 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 20414 705478
rect 19794 702000 20414 705242
rect 23514 702000 24134 707162
rect 27234 702000 27854 709082
rect 30954 702000 31574 711002
rect 48954 710598 49574 711590
rect 48954 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 49574 710598
rect 48954 710278 49574 710362
rect 48954 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 49574 710278
rect 45234 708678 45854 709670
rect 45234 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 45854 708678
rect 45234 708358 45854 708442
rect 45234 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 45854 708358
rect 41514 706758 42134 707750
rect 41514 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 42134 706758
rect 41514 706438 42134 706522
rect 41514 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 42134 706438
rect 37794 704838 38414 705830
rect 37794 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 38414 704838
rect 37794 704518 38414 704602
rect 37794 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 38414 704518
rect 37794 702000 38414 704282
rect 41514 702000 42134 706202
rect 45234 702000 45854 708122
rect 48954 702000 49574 710042
rect 66954 711558 67574 711590
rect 66954 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 67574 711558
rect 66954 711238 67574 711322
rect 66954 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 67574 711238
rect 63234 709638 63854 709670
rect 63234 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 63854 709638
rect 63234 709318 63854 709402
rect 63234 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 63854 709318
rect 59514 707718 60134 707750
rect 59514 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 60134 707718
rect 59514 707398 60134 707482
rect 59514 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 60134 707398
rect 55794 705798 56414 705830
rect 55794 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 56414 705798
rect 55794 705478 56414 705562
rect 55794 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 56414 705478
rect 55794 702000 56414 705242
rect 59514 702000 60134 707162
rect 63234 702000 63854 709082
rect 66954 702000 67574 711002
rect 84954 710598 85574 711590
rect 84954 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 85574 710598
rect 84954 710278 85574 710362
rect 84954 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 85574 710278
rect 81234 708678 81854 709670
rect 81234 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 81854 708678
rect 81234 708358 81854 708442
rect 81234 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 81854 708358
rect 77514 706758 78134 707750
rect 77514 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 78134 706758
rect 77514 706438 78134 706522
rect 77514 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 78134 706438
rect 73794 704838 74414 705830
rect 73794 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 74414 704838
rect 73794 704518 74414 704602
rect 73794 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 74414 704518
rect 73794 702000 74414 704282
rect 77514 702000 78134 706202
rect 81234 702000 81854 708122
rect 84954 702000 85574 710042
rect 102954 711558 103574 711590
rect 102954 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 103574 711558
rect 102954 711238 103574 711322
rect 102954 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 103574 711238
rect 99234 709638 99854 709670
rect 99234 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 99854 709638
rect 99234 709318 99854 709402
rect 99234 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 99854 709318
rect 95514 707718 96134 707750
rect 95514 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 96134 707718
rect 95514 707398 96134 707482
rect 95514 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 96134 707398
rect 91794 705798 92414 705830
rect 91794 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 92414 705798
rect 91794 705478 92414 705562
rect 91794 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 92414 705478
rect 91794 702000 92414 705242
rect 95514 702000 96134 707162
rect 99234 702000 99854 709082
rect 102954 702000 103574 711002
rect 120954 710598 121574 711590
rect 120954 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 121574 710598
rect 120954 710278 121574 710362
rect 120954 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 121574 710278
rect 117234 708678 117854 709670
rect 117234 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 117854 708678
rect 117234 708358 117854 708442
rect 117234 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 117854 708358
rect 113514 706758 114134 707750
rect 113514 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 114134 706758
rect 113514 706438 114134 706522
rect 113514 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 114134 706438
rect 109794 704838 110414 705830
rect 109794 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 110414 704838
rect 109794 704518 110414 704602
rect 109794 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 110414 704518
rect 109794 702000 110414 704282
rect 113514 702000 114134 706202
rect 117234 702000 117854 708122
rect 120954 702000 121574 710042
rect 138954 711558 139574 711590
rect 138954 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 139574 711558
rect 138954 711238 139574 711322
rect 138954 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 139574 711238
rect 135234 709638 135854 709670
rect 135234 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 135854 709638
rect 135234 709318 135854 709402
rect 135234 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 135854 709318
rect 131514 707718 132134 707750
rect 131514 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 132134 707718
rect 131514 707398 132134 707482
rect 131514 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 132134 707398
rect 127794 705798 128414 705830
rect 127794 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 128414 705798
rect 127794 705478 128414 705562
rect 127794 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 128414 705478
rect 127794 702000 128414 705242
rect 131514 702000 132134 707162
rect 135234 702000 135854 709082
rect 138954 702000 139574 711002
rect 156954 710598 157574 711590
rect 156954 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 157574 710598
rect 156954 710278 157574 710362
rect 156954 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 157574 710278
rect 153234 708678 153854 709670
rect 153234 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 153854 708678
rect 153234 708358 153854 708442
rect 153234 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 153854 708358
rect 149514 706758 150134 707750
rect 149514 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 150134 706758
rect 149514 706438 150134 706522
rect 149514 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 150134 706438
rect 145794 704838 146414 705830
rect 145794 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 146414 704838
rect 145794 704518 146414 704602
rect 145794 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 146414 704518
rect 145794 702000 146414 704282
rect 149514 702000 150134 706202
rect 153234 702000 153854 708122
rect 156954 702000 157574 710042
rect 174954 711558 175574 711590
rect 174954 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 175574 711558
rect 174954 711238 175574 711322
rect 174954 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 175574 711238
rect 171234 709638 171854 709670
rect 171234 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 171854 709638
rect 171234 709318 171854 709402
rect 171234 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 171854 709318
rect 167514 707718 168134 707750
rect 167514 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 168134 707718
rect 167514 707398 168134 707482
rect 167514 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 168134 707398
rect 163794 705798 164414 705830
rect 163794 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 164414 705798
rect 163794 705478 164414 705562
rect 163794 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 164414 705478
rect 163794 702000 164414 705242
rect 167514 702000 168134 707162
rect 171234 702000 171854 709082
rect 174954 702000 175574 711002
rect 192954 710598 193574 711590
rect 192954 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 193574 710598
rect 192954 710278 193574 710362
rect 192954 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 193574 710278
rect 189234 708678 189854 709670
rect 189234 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 189854 708678
rect 189234 708358 189854 708442
rect 189234 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 189854 708358
rect 185514 706758 186134 707750
rect 185514 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 186134 706758
rect 185514 706438 186134 706522
rect 185514 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 186134 706438
rect 181794 704838 182414 705830
rect 181794 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 182414 704838
rect 181794 704518 182414 704602
rect 181794 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 182414 704518
rect 181794 702000 182414 704282
rect 185514 702000 186134 706202
rect 189234 702000 189854 708122
rect 192954 702000 193574 710042
rect 210954 711558 211574 711590
rect 210954 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 211574 711558
rect 210954 711238 211574 711322
rect 210954 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 211574 711238
rect 207234 709638 207854 709670
rect 207234 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 207854 709638
rect 207234 709318 207854 709402
rect 207234 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 207854 709318
rect 203514 707718 204134 707750
rect 203514 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 204134 707718
rect 203514 707398 204134 707482
rect 203514 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 204134 707398
rect 199794 705798 200414 705830
rect 199794 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 200414 705798
rect 199794 705478 200414 705562
rect 199794 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 200414 705478
rect 199794 702000 200414 705242
rect 203514 702000 204134 707162
rect 207234 702000 207854 709082
rect 210954 702000 211574 711002
rect 228954 710598 229574 711590
rect 228954 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 229574 710598
rect 228954 710278 229574 710362
rect 228954 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 229574 710278
rect 225234 708678 225854 709670
rect 225234 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 225854 708678
rect 225234 708358 225854 708442
rect 225234 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 225854 708358
rect 221514 706758 222134 707750
rect 221514 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 222134 706758
rect 221514 706438 222134 706522
rect 221514 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 222134 706438
rect 217794 704838 218414 705830
rect 217794 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 218414 704838
rect 217794 704518 218414 704602
rect 217794 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 218414 704518
rect 217794 702000 218414 704282
rect 221514 702000 222134 706202
rect 225234 702000 225854 708122
rect 228954 702000 229574 710042
rect 246954 711558 247574 711590
rect 246954 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 247574 711558
rect 246954 711238 247574 711322
rect 246954 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 247574 711238
rect 243234 709638 243854 709670
rect 243234 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 243854 709638
rect 243234 709318 243854 709402
rect 243234 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 243854 709318
rect 239514 707718 240134 707750
rect 239514 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 240134 707718
rect 239514 707398 240134 707482
rect 239514 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 240134 707398
rect 235794 705798 236414 705830
rect 235794 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 236414 705798
rect 235794 705478 236414 705562
rect 235794 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 236414 705478
rect 235794 702000 236414 705242
rect 239514 702000 240134 707162
rect 243234 702000 243854 709082
rect 246954 702000 247574 711002
rect 264954 710598 265574 711590
rect 264954 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 265574 710598
rect 264954 710278 265574 710362
rect 264954 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 265574 710278
rect 261234 708678 261854 709670
rect 261234 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 261854 708678
rect 261234 708358 261854 708442
rect 261234 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 261854 708358
rect 257514 706758 258134 707750
rect 257514 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 258134 706758
rect 257514 706438 258134 706522
rect 257514 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 258134 706438
rect 253794 704838 254414 705830
rect 253794 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 254414 704838
rect 253794 704518 254414 704602
rect 253794 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 254414 704518
rect 253794 702000 254414 704282
rect 257514 702000 258134 706202
rect 261234 702000 261854 708122
rect 264954 702000 265574 710042
rect 282954 711558 283574 711590
rect 282954 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 283574 711558
rect 282954 711238 283574 711322
rect 282954 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 283574 711238
rect 279234 709638 279854 709670
rect 279234 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 279854 709638
rect 279234 709318 279854 709402
rect 279234 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 279854 709318
rect 275514 707718 276134 707750
rect 275514 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 276134 707718
rect 275514 707398 276134 707482
rect 275514 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 276134 707398
rect 271794 705798 272414 705830
rect 271794 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 272414 705798
rect 271794 705478 272414 705562
rect 271794 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 272414 705478
rect 271794 702000 272414 705242
rect 275514 702000 276134 707162
rect 279234 702000 279854 709082
rect 282954 702000 283574 711002
rect 300954 710598 301574 711590
rect 300954 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 301574 710598
rect 300954 710278 301574 710362
rect 300954 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 301574 710278
rect 297234 708678 297854 709670
rect 297234 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 297854 708678
rect 297234 708358 297854 708442
rect 297234 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 297854 708358
rect 293514 706758 294134 707750
rect 293514 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 294134 706758
rect 293514 706438 294134 706522
rect 293514 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 294134 706438
rect 289794 704838 290414 705830
rect 289794 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 290414 704838
rect 289794 704518 290414 704602
rect 289794 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 290414 704518
rect 289794 702000 290414 704282
rect 293514 702000 294134 706202
rect 297234 702000 297854 708122
rect 300954 702000 301574 710042
rect 318954 711558 319574 711590
rect 318954 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 319574 711558
rect 318954 711238 319574 711322
rect 318954 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 319574 711238
rect 315234 709638 315854 709670
rect 315234 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 315854 709638
rect 315234 709318 315854 709402
rect 315234 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 315854 709318
rect 311514 707718 312134 707750
rect 311514 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 312134 707718
rect 311514 707398 312134 707482
rect 311514 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 312134 707398
rect 307794 705798 308414 705830
rect 307794 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 308414 705798
rect 307794 705478 308414 705562
rect 307794 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 308414 705478
rect 307794 702000 308414 705242
rect 311514 702000 312134 707162
rect 315234 702000 315854 709082
rect 318954 702000 319574 711002
rect 336954 710598 337574 711590
rect 336954 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 337574 710598
rect 336954 710278 337574 710362
rect 336954 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 337574 710278
rect 333234 708678 333854 709670
rect 333234 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 333854 708678
rect 333234 708358 333854 708442
rect 333234 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 333854 708358
rect 329514 706758 330134 707750
rect 329514 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 330134 706758
rect 329514 706438 330134 706522
rect 329514 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 330134 706438
rect 325794 704838 326414 705830
rect 325794 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 326414 704838
rect 325794 704518 326414 704602
rect 325794 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 326414 704518
rect 325794 702000 326414 704282
rect 329514 702000 330134 706202
rect 333234 702000 333854 708122
rect 336954 702000 337574 710042
rect 354954 711558 355574 711590
rect 354954 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 355574 711558
rect 354954 711238 355574 711322
rect 354954 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 355574 711238
rect 351234 709638 351854 709670
rect 351234 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 351854 709638
rect 351234 709318 351854 709402
rect 351234 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 351854 709318
rect 347514 707718 348134 707750
rect 347514 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 348134 707718
rect 347514 707398 348134 707482
rect 347514 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 348134 707398
rect 343794 705798 344414 705830
rect 343794 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 344414 705798
rect 343794 705478 344414 705562
rect 343794 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 344414 705478
rect 343794 702000 344414 705242
rect 347514 702000 348134 707162
rect 351234 702000 351854 709082
rect 354954 702000 355574 711002
rect 372954 710598 373574 711590
rect 372954 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 373574 710598
rect 372954 710278 373574 710362
rect 372954 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 373574 710278
rect 369234 708678 369854 709670
rect 369234 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 369854 708678
rect 369234 708358 369854 708442
rect 369234 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 369854 708358
rect 365514 706758 366134 707750
rect 365514 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 366134 706758
rect 365514 706438 366134 706522
rect 365514 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 366134 706438
rect 361794 704838 362414 705830
rect 361794 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 362414 704838
rect 361794 704518 362414 704602
rect 361794 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 362414 704518
rect 361794 702000 362414 704282
rect 365514 702000 366134 706202
rect 369234 702000 369854 708122
rect 372954 702000 373574 710042
rect 390954 711558 391574 711590
rect 390954 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 391574 711558
rect 390954 711238 391574 711322
rect 390954 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 391574 711238
rect 387234 709638 387854 709670
rect 387234 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 387854 709638
rect 387234 709318 387854 709402
rect 387234 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 387854 709318
rect 383514 707718 384134 707750
rect 383514 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 384134 707718
rect 383514 707398 384134 707482
rect 383514 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 384134 707398
rect 379794 705798 380414 705830
rect 379794 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 380414 705798
rect 379794 705478 380414 705562
rect 379794 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 380414 705478
rect 379794 702000 380414 705242
rect 383514 702000 384134 707162
rect 387234 702000 387854 709082
rect 390954 702000 391574 711002
rect 408954 710598 409574 711590
rect 408954 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 409574 710598
rect 408954 710278 409574 710362
rect 408954 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 409574 710278
rect 405234 708678 405854 709670
rect 405234 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 405854 708678
rect 405234 708358 405854 708442
rect 405234 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 405854 708358
rect 401514 706758 402134 707750
rect 401514 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 402134 706758
rect 401514 706438 402134 706522
rect 401514 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 402134 706438
rect 397794 704838 398414 705830
rect 397794 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 398414 704838
rect 397794 704518 398414 704602
rect 397794 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 398414 704518
rect 397794 702000 398414 704282
rect 401514 702000 402134 706202
rect 405234 702000 405854 708122
rect 408954 702000 409574 710042
rect 426954 711558 427574 711590
rect 426954 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 427574 711558
rect 426954 711238 427574 711322
rect 426954 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 427574 711238
rect 423234 709638 423854 709670
rect 423234 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 423854 709638
rect 423234 709318 423854 709402
rect 423234 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 423854 709318
rect 419514 707718 420134 707750
rect 419514 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 420134 707718
rect 419514 707398 420134 707482
rect 419514 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 420134 707398
rect 415794 705798 416414 705830
rect 415794 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 416414 705798
rect 415794 705478 416414 705562
rect 415794 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 416414 705478
rect 415794 702000 416414 705242
rect 419514 702000 420134 707162
rect 423234 702000 423854 709082
rect 426954 702000 427574 711002
rect 444954 710598 445574 711590
rect 444954 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 445574 710598
rect 444954 710278 445574 710362
rect 444954 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 445574 710278
rect 441234 708678 441854 709670
rect 441234 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 441854 708678
rect 441234 708358 441854 708442
rect 441234 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 441854 708358
rect 437514 706758 438134 707750
rect 437514 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 438134 706758
rect 437514 706438 438134 706522
rect 437514 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 438134 706438
rect 433794 704838 434414 705830
rect 433794 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 434414 704838
rect 433794 704518 434414 704602
rect 433794 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 434414 704518
rect 433794 702000 434414 704282
rect 437514 702000 438134 706202
rect 441234 702000 441854 708122
rect 444954 702000 445574 710042
rect 462954 711558 463574 711590
rect 462954 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 463574 711558
rect 462954 711238 463574 711322
rect 462954 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 463574 711238
rect 459234 709638 459854 709670
rect 459234 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 459854 709638
rect 459234 709318 459854 709402
rect 459234 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 459854 709318
rect 455514 707718 456134 707750
rect 455514 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 456134 707718
rect 455514 707398 456134 707482
rect 455514 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 456134 707398
rect 451794 705798 452414 705830
rect 451794 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 452414 705798
rect 451794 705478 452414 705562
rect 451794 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 452414 705478
rect 451794 702000 452414 705242
rect 455514 702000 456134 707162
rect 459234 702000 459854 709082
rect 462954 702000 463574 711002
rect 480954 710598 481574 711590
rect 480954 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 481574 710598
rect 480954 710278 481574 710362
rect 480954 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 481574 710278
rect 477234 708678 477854 709670
rect 477234 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 477854 708678
rect 477234 708358 477854 708442
rect 477234 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 477854 708358
rect 473514 706758 474134 707750
rect 473514 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 474134 706758
rect 473514 706438 474134 706522
rect 473514 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 474134 706438
rect 469794 704838 470414 705830
rect 469794 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 470414 704838
rect 469794 704518 470414 704602
rect 469794 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 470414 704518
rect 469794 702000 470414 704282
rect 473514 702000 474134 706202
rect 477234 702000 477854 708122
rect 480954 702000 481574 710042
rect 498954 711558 499574 711590
rect 498954 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 499574 711558
rect 498954 711238 499574 711322
rect 498954 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 499574 711238
rect 495234 709638 495854 709670
rect 495234 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 495854 709638
rect 495234 709318 495854 709402
rect 495234 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 495854 709318
rect 491514 707718 492134 707750
rect 491514 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 492134 707718
rect 491514 707398 492134 707482
rect 491514 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 492134 707398
rect 487794 705798 488414 705830
rect 487794 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 488414 705798
rect 487794 705478 488414 705562
rect 487794 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 488414 705478
rect 487794 702000 488414 705242
rect 491514 702000 492134 707162
rect 495234 702000 495854 709082
rect 498954 702000 499574 711002
rect 516954 710598 517574 711590
rect 516954 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 517574 710598
rect 516954 710278 517574 710362
rect 516954 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 517574 710278
rect 513234 708678 513854 709670
rect 513234 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 513854 708678
rect 513234 708358 513854 708442
rect 513234 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 513854 708358
rect 509514 706758 510134 707750
rect 509514 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 510134 706758
rect 509514 706438 510134 706522
rect 509514 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 510134 706438
rect 505794 704838 506414 705830
rect 505794 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 506414 704838
rect 505794 704518 506414 704602
rect 505794 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 506414 704518
rect 505794 702000 506414 704282
rect 509514 702000 510134 706202
rect 513234 702000 513854 708122
rect 516954 702000 517574 710042
rect 534954 711558 535574 711590
rect 534954 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 535574 711558
rect 534954 711238 535574 711322
rect 534954 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 535574 711238
rect 531234 709638 531854 709670
rect 531234 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 531854 709638
rect 531234 709318 531854 709402
rect 531234 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 531854 709318
rect 527514 707718 528134 707750
rect 527514 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 528134 707718
rect 527514 707398 528134 707482
rect 527514 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 528134 707398
rect 523794 705798 524414 705830
rect 523794 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 524414 705798
rect 523794 705478 524414 705562
rect 523794 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 524414 705478
rect 523794 702000 524414 705242
rect 527514 702000 528134 707162
rect 531234 702000 531854 709082
rect 534954 702000 535574 711002
rect 552954 710598 553574 711590
rect 552954 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 553574 710598
rect 552954 710278 553574 710362
rect 552954 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 553574 710278
rect 549234 708678 549854 709670
rect 549234 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 549854 708678
rect 549234 708358 549854 708442
rect 549234 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 549854 708358
rect 545514 706758 546134 707750
rect 545514 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 546134 706758
rect 545514 706438 546134 706522
rect 545514 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 546134 706438
rect 541794 704838 542414 705830
rect 541794 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 542414 704838
rect 541794 704518 542414 704602
rect 541794 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 542414 704518
rect 541794 702000 542414 704282
rect 545514 702000 546134 706202
rect 549234 702000 549854 708122
rect 552954 702000 553574 710042
rect 570954 711558 571574 711590
rect 570954 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 571574 711558
rect 570954 711238 571574 711322
rect 570954 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 571574 711238
rect 567234 709638 567854 709670
rect 567234 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 567854 709638
rect 567234 709318 567854 709402
rect 567234 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 567854 709318
rect 563514 707718 564134 707750
rect 563514 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 564134 707718
rect 563514 707398 564134 707482
rect 563514 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 564134 707398
rect 559794 705798 560414 705830
rect 559794 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 560414 705798
rect 559794 705478 560414 705562
rect 559794 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 560414 705478
rect 559794 702000 560414 705242
rect 563514 702000 564134 707162
rect 453987 701996 454053 701997
rect 453987 701932 453988 701996
rect 454052 701932 454053 701996
rect 453987 701931 454053 701932
rect 259131 701724 259197 701725
rect 259131 701660 259132 701724
rect 259196 701660 259197 701724
rect 259131 701659 259197 701660
rect 13859 699412 13925 699413
rect 13859 699348 13860 699412
rect 13924 699348 13925 699412
rect 13859 699347 13925 699348
rect 43115 699412 43181 699413
rect 43115 699348 43116 699412
rect 43180 699348 43181 699412
rect 43115 699347 43181 699348
rect 52867 699412 52933 699413
rect 52867 699348 52868 699412
rect 52932 699348 52933 699412
rect 52867 699347 52933 699348
rect 60227 699412 60293 699413
rect 60227 699348 60228 699412
rect 60292 699348 60293 699412
rect 60227 699347 60293 699348
rect 124627 699412 124693 699413
rect 124627 699348 124628 699412
rect 124692 699348 124693 699412
rect 124627 699347 124693 699348
rect 13862 698325 13922 699347
rect 43118 698597 43178 699347
rect 52870 698733 52930 699347
rect 60230 698869 60290 699347
rect 124443 699140 124509 699141
rect 124443 699076 124444 699140
rect 124508 699076 124509 699140
rect 124443 699075 124509 699076
rect 60227 698868 60293 698869
rect 60227 698804 60228 698868
rect 60292 698804 60293 698868
rect 60227 698803 60293 698804
rect 52867 698732 52933 698733
rect 52867 698668 52868 698732
rect 52932 698668 52933 698732
rect 52867 698667 52933 698668
rect 43115 698596 43181 698597
rect 43115 698532 43116 698596
rect 43180 698532 43181 698596
rect 43115 698531 43181 698532
rect 13859 698324 13925 698325
rect 13859 698260 13860 698324
rect 13924 698260 13925 698324
rect 13859 698259 13925 698260
rect 124446 697917 124506 699075
rect 124630 697917 124690 699347
rect 259134 699141 259194 701659
rect 453990 699549 454050 701931
rect 453987 699548 454053 699549
rect 453987 699484 453988 699548
rect 454052 699484 454053 699548
rect 453987 699483 454053 699484
rect 418659 699412 418725 699413
rect 418659 699348 418660 699412
rect 418724 699348 418725 699412
rect 418659 699347 418725 699348
rect 433379 699412 433445 699413
rect 433379 699348 433380 699412
rect 433444 699348 433445 699412
rect 433379 699347 433445 699348
rect 462819 699412 462885 699413
rect 462819 699348 462820 699412
rect 462884 699348 462885 699412
rect 462819 699347 462885 699348
rect 492627 699412 492693 699413
rect 492627 699348 492628 699412
rect 492692 699348 492693 699412
rect 492627 699347 492693 699348
rect 510659 699412 510725 699413
rect 510659 699348 510660 699412
rect 510724 699348 510725 699412
rect 510659 699347 510725 699348
rect 539915 699412 539981 699413
rect 539915 699348 539916 699412
rect 539980 699348 539981 699412
rect 539915 699347 539981 699348
rect 259131 699140 259197 699141
rect 259131 699076 259132 699140
rect 259196 699076 259197 699140
rect 259131 699075 259197 699076
rect 418662 698189 418722 699347
rect 418659 698188 418725 698189
rect 418659 698124 418660 698188
rect 418724 698124 418725 698188
rect 418659 698123 418725 698124
rect 433382 698053 433442 699347
rect 433379 698052 433445 698053
rect 433379 697988 433380 698052
rect 433444 697988 433445 698052
rect 433379 697987 433445 697988
rect 124443 697916 124509 697917
rect 124443 697852 124444 697916
rect 124508 697852 124509 697916
rect 124443 697851 124509 697852
rect 124627 697916 124693 697917
rect 124627 697852 124628 697916
rect 124692 697852 124693 697916
rect 124627 697851 124693 697852
rect 462822 697781 462882 699347
rect 462819 697780 462885 697781
rect 462819 697716 462820 697780
rect 462884 697716 462885 697780
rect 462819 697715 462885 697716
rect 492630 697645 492690 699347
rect 510662 699005 510722 699347
rect 510659 699004 510725 699005
rect 510659 698940 510660 699004
rect 510724 698940 510725 699004
rect 510659 698939 510725 698940
rect 539918 698461 539978 699347
rect 539915 698460 539981 698461
rect 539915 698396 539916 698460
rect 539980 698396 539981 698460
rect 539915 698395 539981 698396
rect 492627 697644 492693 697645
rect 492627 697580 492628 697644
rect 492692 697580 492693 697644
rect 492627 697579 492693 697580
rect -2006 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 -1386 687454
rect -2006 687134 -1386 687218
rect -2006 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 -1386 687134
rect -2006 651454 -1386 686898
rect 8208 687454 8528 687486
rect 8208 687218 8250 687454
rect 8486 687218 8528 687454
rect 8208 687134 8528 687218
rect 8208 686898 8250 687134
rect 8486 686898 8528 687134
rect 8208 686866 8528 686898
rect 38928 687454 39248 687486
rect 38928 687218 38970 687454
rect 39206 687218 39248 687454
rect 38928 687134 39248 687218
rect 38928 686898 38970 687134
rect 39206 686898 39248 687134
rect 38928 686866 39248 686898
rect 69648 687454 69968 687486
rect 69648 687218 69690 687454
rect 69926 687218 69968 687454
rect 69648 687134 69968 687218
rect 69648 686898 69690 687134
rect 69926 686898 69968 687134
rect 69648 686866 69968 686898
rect 100368 687454 100688 687486
rect 100368 687218 100410 687454
rect 100646 687218 100688 687454
rect 100368 687134 100688 687218
rect 100368 686898 100410 687134
rect 100646 686898 100688 687134
rect 100368 686866 100688 686898
rect 131088 687454 131408 687486
rect 131088 687218 131130 687454
rect 131366 687218 131408 687454
rect 131088 687134 131408 687218
rect 131088 686898 131130 687134
rect 131366 686898 131408 687134
rect 131088 686866 131408 686898
rect 161808 687454 162128 687486
rect 161808 687218 161850 687454
rect 162086 687218 162128 687454
rect 161808 687134 162128 687218
rect 161808 686898 161850 687134
rect 162086 686898 162128 687134
rect 161808 686866 162128 686898
rect 192528 687454 192848 687486
rect 192528 687218 192570 687454
rect 192806 687218 192848 687454
rect 192528 687134 192848 687218
rect 192528 686898 192570 687134
rect 192806 686898 192848 687134
rect 192528 686866 192848 686898
rect 223248 687454 223568 687486
rect 223248 687218 223290 687454
rect 223526 687218 223568 687454
rect 223248 687134 223568 687218
rect 223248 686898 223290 687134
rect 223526 686898 223568 687134
rect 223248 686866 223568 686898
rect 253968 687454 254288 687486
rect 253968 687218 254010 687454
rect 254246 687218 254288 687454
rect 253968 687134 254288 687218
rect 253968 686898 254010 687134
rect 254246 686898 254288 687134
rect 253968 686866 254288 686898
rect 284688 687454 285008 687486
rect 284688 687218 284730 687454
rect 284966 687218 285008 687454
rect 284688 687134 285008 687218
rect 284688 686898 284730 687134
rect 284966 686898 285008 687134
rect 284688 686866 285008 686898
rect 315408 687454 315728 687486
rect 315408 687218 315450 687454
rect 315686 687218 315728 687454
rect 315408 687134 315728 687218
rect 315408 686898 315450 687134
rect 315686 686898 315728 687134
rect 315408 686866 315728 686898
rect 346128 687454 346448 687486
rect 346128 687218 346170 687454
rect 346406 687218 346448 687454
rect 346128 687134 346448 687218
rect 346128 686898 346170 687134
rect 346406 686898 346448 687134
rect 346128 686866 346448 686898
rect 376848 687454 377168 687486
rect 376848 687218 376890 687454
rect 377126 687218 377168 687454
rect 376848 687134 377168 687218
rect 376848 686898 376890 687134
rect 377126 686898 377168 687134
rect 376848 686866 377168 686898
rect 407568 687454 407888 687486
rect 407568 687218 407610 687454
rect 407846 687218 407888 687454
rect 407568 687134 407888 687218
rect 407568 686898 407610 687134
rect 407846 686898 407888 687134
rect 407568 686866 407888 686898
rect 438288 687454 438608 687486
rect 438288 687218 438330 687454
rect 438566 687218 438608 687454
rect 438288 687134 438608 687218
rect 438288 686898 438330 687134
rect 438566 686898 438608 687134
rect 438288 686866 438608 686898
rect 469008 687454 469328 687486
rect 469008 687218 469050 687454
rect 469286 687218 469328 687454
rect 469008 687134 469328 687218
rect 469008 686898 469050 687134
rect 469286 686898 469328 687134
rect 469008 686866 469328 686898
rect 499728 687454 500048 687486
rect 499728 687218 499770 687454
rect 500006 687218 500048 687454
rect 499728 687134 500048 687218
rect 499728 686898 499770 687134
rect 500006 686898 500048 687134
rect 499728 686866 500048 686898
rect 530448 687454 530768 687486
rect 530448 687218 530490 687454
rect 530726 687218 530768 687454
rect 530448 687134 530768 687218
rect 530448 686898 530490 687134
rect 530726 686898 530768 687134
rect 530448 686866 530768 686898
rect 561168 687454 561488 687486
rect 561168 687218 561210 687454
rect 561446 687218 561488 687454
rect 561168 687134 561488 687218
rect 561168 686898 561210 687134
rect 561446 686898 561488 687134
rect 561168 686866 561488 686898
rect 567234 676894 567854 709082
rect 567234 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 567854 676894
rect 567234 676574 567854 676658
rect 567234 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 567854 676574
rect 23568 669454 23888 669486
rect 23568 669218 23610 669454
rect 23846 669218 23888 669454
rect 23568 669134 23888 669218
rect 23568 668898 23610 669134
rect 23846 668898 23888 669134
rect 23568 668866 23888 668898
rect 54288 669454 54608 669486
rect 54288 669218 54330 669454
rect 54566 669218 54608 669454
rect 54288 669134 54608 669218
rect 54288 668898 54330 669134
rect 54566 668898 54608 669134
rect 54288 668866 54608 668898
rect 85008 669454 85328 669486
rect 85008 669218 85050 669454
rect 85286 669218 85328 669454
rect 85008 669134 85328 669218
rect 85008 668898 85050 669134
rect 85286 668898 85328 669134
rect 85008 668866 85328 668898
rect 115728 669454 116048 669486
rect 115728 669218 115770 669454
rect 116006 669218 116048 669454
rect 115728 669134 116048 669218
rect 115728 668898 115770 669134
rect 116006 668898 116048 669134
rect 115728 668866 116048 668898
rect 146448 669454 146768 669486
rect 146448 669218 146490 669454
rect 146726 669218 146768 669454
rect 146448 669134 146768 669218
rect 146448 668898 146490 669134
rect 146726 668898 146768 669134
rect 146448 668866 146768 668898
rect 177168 669454 177488 669486
rect 177168 669218 177210 669454
rect 177446 669218 177488 669454
rect 177168 669134 177488 669218
rect 177168 668898 177210 669134
rect 177446 668898 177488 669134
rect 177168 668866 177488 668898
rect 207888 669454 208208 669486
rect 207888 669218 207930 669454
rect 208166 669218 208208 669454
rect 207888 669134 208208 669218
rect 207888 668898 207930 669134
rect 208166 668898 208208 669134
rect 207888 668866 208208 668898
rect 238608 669454 238928 669486
rect 238608 669218 238650 669454
rect 238886 669218 238928 669454
rect 238608 669134 238928 669218
rect 238608 668898 238650 669134
rect 238886 668898 238928 669134
rect 238608 668866 238928 668898
rect 269328 669454 269648 669486
rect 269328 669218 269370 669454
rect 269606 669218 269648 669454
rect 269328 669134 269648 669218
rect 269328 668898 269370 669134
rect 269606 668898 269648 669134
rect 269328 668866 269648 668898
rect 300048 669454 300368 669486
rect 300048 669218 300090 669454
rect 300326 669218 300368 669454
rect 300048 669134 300368 669218
rect 300048 668898 300090 669134
rect 300326 668898 300368 669134
rect 300048 668866 300368 668898
rect 330768 669454 331088 669486
rect 330768 669218 330810 669454
rect 331046 669218 331088 669454
rect 330768 669134 331088 669218
rect 330768 668898 330810 669134
rect 331046 668898 331088 669134
rect 330768 668866 331088 668898
rect 361488 669454 361808 669486
rect 361488 669218 361530 669454
rect 361766 669218 361808 669454
rect 361488 669134 361808 669218
rect 361488 668898 361530 669134
rect 361766 668898 361808 669134
rect 361488 668866 361808 668898
rect 392208 669454 392528 669486
rect 392208 669218 392250 669454
rect 392486 669218 392528 669454
rect 392208 669134 392528 669218
rect 392208 668898 392250 669134
rect 392486 668898 392528 669134
rect 392208 668866 392528 668898
rect 422928 669454 423248 669486
rect 422928 669218 422970 669454
rect 423206 669218 423248 669454
rect 422928 669134 423248 669218
rect 422928 668898 422970 669134
rect 423206 668898 423248 669134
rect 422928 668866 423248 668898
rect 453648 669454 453968 669486
rect 453648 669218 453690 669454
rect 453926 669218 453968 669454
rect 453648 669134 453968 669218
rect 453648 668898 453690 669134
rect 453926 668898 453968 669134
rect 453648 668866 453968 668898
rect 484368 669454 484688 669486
rect 484368 669218 484410 669454
rect 484646 669218 484688 669454
rect 484368 669134 484688 669218
rect 484368 668898 484410 669134
rect 484646 668898 484688 669134
rect 484368 668866 484688 668898
rect 515088 669454 515408 669486
rect 515088 669218 515130 669454
rect 515366 669218 515408 669454
rect 515088 669134 515408 669218
rect 515088 668898 515130 669134
rect 515366 668898 515408 669134
rect 515088 668866 515408 668898
rect 545808 669454 546128 669486
rect 545808 669218 545850 669454
rect 546086 669218 546128 669454
rect 545808 669134 546128 669218
rect 545808 668898 545850 669134
rect 546086 668898 546128 669134
rect 545808 668866 546128 668898
rect -2006 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 -1386 651454
rect -2006 651134 -1386 651218
rect -2006 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 -1386 651134
rect -2006 615454 -1386 650898
rect 8208 651454 8528 651486
rect 8208 651218 8250 651454
rect 8486 651218 8528 651454
rect 8208 651134 8528 651218
rect 8208 650898 8250 651134
rect 8486 650898 8528 651134
rect 8208 650866 8528 650898
rect 38928 651454 39248 651486
rect 38928 651218 38970 651454
rect 39206 651218 39248 651454
rect 38928 651134 39248 651218
rect 38928 650898 38970 651134
rect 39206 650898 39248 651134
rect 38928 650866 39248 650898
rect 69648 651454 69968 651486
rect 69648 651218 69690 651454
rect 69926 651218 69968 651454
rect 69648 651134 69968 651218
rect 69648 650898 69690 651134
rect 69926 650898 69968 651134
rect 69648 650866 69968 650898
rect 100368 651454 100688 651486
rect 100368 651218 100410 651454
rect 100646 651218 100688 651454
rect 100368 651134 100688 651218
rect 100368 650898 100410 651134
rect 100646 650898 100688 651134
rect 100368 650866 100688 650898
rect 131088 651454 131408 651486
rect 131088 651218 131130 651454
rect 131366 651218 131408 651454
rect 131088 651134 131408 651218
rect 131088 650898 131130 651134
rect 131366 650898 131408 651134
rect 131088 650866 131408 650898
rect 161808 651454 162128 651486
rect 161808 651218 161850 651454
rect 162086 651218 162128 651454
rect 161808 651134 162128 651218
rect 161808 650898 161850 651134
rect 162086 650898 162128 651134
rect 161808 650866 162128 650898
rect 192528 651454 192848 651486
rect 192528 651218 192570 651454
rect 192806 651218 192848 651454
rect 192528 651134 192848 651218
rect 192528 650898 192570 651134
rect 192806 650898 192848 651134
rect 192528 650866 192848 650898
rect 223248 651454 223568 651486
rect 223248 651218 223290 651454
rect 223526 651218 223568 651454
rect 223248 651134 223568 651218
rect 223248 650898 223290 651134
rect 223526 650898 223568 651134
rect 223248 650866 223568 650898
rect 253968 651454 254288 651486
rect 253968 651218 254010 651454
rect 254246 651218 254288 651454
rect 253968 651134 254288 651218
rect 253968 650898 254010 651134
rect 254246 650898 254288 651134
rect 253968 650866 254288 650898
rect 284688 651454 285008 651486
rect 284688 651218 284730 651454
rect 284966 651218 285008 651454
rect 284688 651134 285008 651218
rect 284688 650898 284730 651134
rect 284966 650898 285008 651134
rect 284688 650866 285008 650898
rect 315408 651454 315728 651486
rect 315408 651218 315450 651454
rect 315686 651218 315728 651454
rect 315408 651134 315728 651218
rect 315408 650898 315450 651134
rect 315686 650898 315728 651134
rect 315408 650866 315728 650898
rect 346128 651454 346448 651486
rect 346128 651218 346170 651454
rect 346406 651218 346448 651454
rect 346128 651134 346448 651218
rect 346128 650898 346170 651134
rect 346406 650898 346448 651134
rect 346128 650866 346448 650898
rect 376848 651454 377168 651486
rect 376848 651218 376890 651454
rect 377126 651218 377168 651454
rect 376848 651134 377168 651218
rect 376848 650898 376890 651134
rect 377126 650898 377168 651134
rect 376848 650866 377168 650898
rect 407568 651454 407888 651486
rect 407568 651218 407610 651454
rect 407846 651218 407888 651454
rect 407568 651134 407888 651218
rect 407568 650898 407610 651134
rect 407846 650898 407888 651134
rect 407568 650866 407888 650898
rect 438288 651454 438608 651486
rect 438288 651218 438330 651454
rect 438566 651218 438608 651454
rect 438288 651134 438608 651218
rect 438288 650898 438330 651134
rect 438566 650898 438608 651134
rect 438288 650866 438608 650898
rect 469008 651454 469328 651486
rect 469008 651218 469050 651454
rect 469286 651218 469328 651454
rect 469008 651134 469328 651218
rect 469008 650898 469050 651134
rect 469286 650898 469328 651134
rect 469008 650866 469328 650898
rect 499728 651454 500048 651486
rect 499728 651218 499770 651454
rect 500006 651218 500048 651454
rect 499728 651134 500048 651218
rect 499728 650898 499770 651134
rect 500006 650898 500048 651134
rect 499728 650866 500048 650898
rect 530448 651454 530768 651486
rect 530448 651218 530490 651454
rect 530726 651218 530768 651454
rect 530448 651134 530768 651218
rect 530448 650898 530490 651134
rect 530726 650898 530768 651134
rect 530448 650866 530768 650898
rect 561168 651454 561488 651486
rect 561168 651218 561210 651454
rect 561446 651218 561488 651454
rect 561168 651134 561488 651218
rect 561168 650898 561210 651134
rect 561446 650898 561488 651134
rect 561168 650866 561488 650898
rect 567234 640894 567854 676338
rect 567234 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 567854 640894
rect 567234 640574 567854 640658
rect 567234 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 567854 640574
rect 23568 633454 23888 633486
rect 23568 633218 23610 633454
rect 23846 633218 23888 633454
rect 23568 633134 23888 633218
rect 23568 632898 23610 633134
rect 23846 632898 23888 633134
rect 23568 632866 23888 632898
rect 54288 633454 54608 633486
rect 54288 633218 54330 633454
rect 54566 633218 54608 633454
rect 54288 633134 54608 633218
rect 54288 632898 54330 633134
rect 54566 632898 54608 633134
rect 54288 632866 54608 632898
rect 85008 633454 85328 633486
rect 85008 633218 85050 633454
rect 85286 633218 85328 633454
rect 85008 633134 85328 633218
rect 85008 632898 85050 633134
rect 85286 632898 85328 633134
rect 85008 632866 85328 632898
rect 115728 633454 116048 633486
rect 115728 633218 115770 633454
rect 116006 633218 116048 633454
rect 115728 633134 116048 633218
rect 115728 632898 115770 633134
rect 116006 632898 116048 633134
rect 115728 632866 116048 632898
rect 146448 633454 146768 633486
rect 146448 633218 146490 633454
rect 146726 633218 146768 633454
rect 146448 633134 146768 633218
rect 146448 632898 146490 633134
rect 146726 632898 146768 633134
rect 146448 632866 146768 632898
rect 177168 633454 177488 633486
rect 177168 633218 177210 633454
rect 177446 633218 177488 633454
rect 177168 633134 177488 633218
rect 177168 632898 177210 633134
rect 177446 632898 177488 633134
rect 177168 632866 177488 632898
rect 207888 633454 208208 633486
rect 207888 633218 207930 633454
rect 208166 633218 208208 633454
rect 207888 633134 208208 633218
rect 207888 632898 207930 633134
rect 208166 632898 208208 633134
rect 207888 632866 208208 632898
rect 238608 633454 238928 633486
rect 238608 633218 238650 633454
rect 238886 633218 238928 633454
rect 238608 633134 238928 633218
rect 238608 632898 238650 633134
rect 238886 632898 238928 633134
rect 238608 632866 238928 632898
rect 269328 633454 269648 633486
rect 269328 633218 269370 633454
rect 269606 633218 269648 633454
rect 269328 633134 269648 633218
rect 269328 632898 269370 633134
rect 269606 632898 269648 633134
rect 269328 632866 269648 632898
rect 300048 633454 300368 633486
rect 300048 633218 300090 633454
rect 300326 633218 300368 633454
rect 300048 633134 300368 633218
rect 300048 632898 300090 633134
rect 300326 632898 300368 633134
rect 300048 632866 300368 632898
rect 330768 633454 331088 633486
rect 330768 633218 330810 633454
rect 331046 633218 331088 633454
rect 330768 633134 331088 633218
rect 330768 632898 330810 633134
rect 331046 632898 331088 633134
rect 330768 632866 331088 632898
rect 361488 633454 361808 633486
rect 361488 633218 361530 633454
rect 361766 633218 361808 633454
rect 361488 633134 361808 633218
rect 361488 632898 361530 633134
rect 361766 632898 361808 633134
rect 361488 632866 361808 632898
rect 392208 633454 392528 633486
rect 392208 633218 392250 633454
rect 392486 633218 392528 633454
rect 392208 633134 392528 633218
rect 392208 632898 392250 633134
rect 392486 632898 392528 633134
rect 392208 632866 392528 632898
rect 422928 633454 423248 633486
rect 422928 633218 422970 633454
rect 423206 633218 423248 633454
rect 422928 633134 423248 633218
rect 422928 632898 422970 633134
rect 423206 632898 423248 633134
rect 422928 632866 423248 632898
rect 453648 633454 453968 633486
rect 453648 633218 453690 633454
rect 453926 633218 453968 633454
rect 453648 633134 453968 633218
rect 453648 632898 453690 633134
rect 453926 632898 453968 633134
rect 453648 632866 453968 632898
rect 484368 633454 484688 633486
rect 484368 633218 484410 633454
rect 484646 633218 484688 633454
rect 484368 633134 484688 633218
rect 484368 632898 484410 633134
rect 484646 632898 484688 633134
rect 484368 632866 484688 632898
rect 515088 633454 515408 633486
rect 515088 633218 515130 633454
rect 515366 633218 515408 633454
rect 515088 633134 515408 633218
rect 515088 632898 515130 633134
rect 515366 632898 515408 633134
rect 515088 632866 515408 632898
rect 545808 633454 546128 633486
rect 545808 633218 545850 633454
rect 546086 633218 546128 633454
rect 545808 633134 546128 633218
rect 545808 632898 545850 633134
rect 546086 632898 546128 633134
rect 545808 632866 546128 632898
rect -2006 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 -1386 615454
rect -2006 615134 -1386 615218
rect -2006 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 -1386 615134
rect -2006 579454 -1386 614898
rect 8208 615454 8528 615486
rect 8208 615218 8250 615454
rect 8486 615218 8528 615454
rect 8208 615134 8528 615218
rect 8208 614898 8250 615134
rect 8486 614898 8528 615134
rect 8208 614866 8528 614898
rect 38928 615454 39248 615486
rect 38928 615218 38970 615454
rect 39206 615218 39248 615454
rect 38928 615134 39248 615218
rect 38928 614898 38970 615134
rect 39206 614898 39248 615134
rect 38928 614866 39248 614898
rect 69648 615454 69968 615486
rect 69648 615218 69690 615454
rect 69926 615218 69968 615454
rect 69648 615134 69968 615218
rect 69648 614898 69690 615134
rect 69926 614898 69968 615134
rect 69648 614866 69968 614898
rect 100368 615454 100688 615486
rect 100368 615218 100410 615454
rect 100646 615218 100688 615454
rect 100368 615134 100688 615218
rect 100368 614898 100410 615134
rect 100646 614898 100688 615134
rect 100368 614866 100688 614898
rect 131088 615454 131408 615486
rect 131088 615218 131130 615454
rect 131366 615218 131408 615454
rect 131088 615134 131408 615218
rect 131088 614898 131130 615134
rect 131366 614898 131408 615134
rect 131088 614866 131408 614898
rect 161808 615454 162128 615486
rect 161808 615218 161850 615454
rect 162086 615218 162128 615454
rect 161808 615134 162128 615218
rect 161808 614898 161850 615134
rect 162086 614898 162128 615134
rect 161808 614866 162128 614898
rect 192528 615454 192848 615486
rect 192528 615218 192570 615454
rect 192806 615218 192848 615454
rect 192528 615134 192848 615218
rect 192528 614898 192570 615134
rect 192806 614898 192848 615134
rect 192528 614866 192848 614898
rect 223248 615454 223568 615486
rect 223248 615218 223290 615454
rect 223526 615218 223568 615454
rect 223248 615134 223568 615218
rect 223248 614898 223290 615134
rect 223526 614898 223568 615134
rect 223248 614866 223568 614898
rect 253968 615454 254288 615486
rect 253968 615218 254010 615454
rect 254246 615218 254288 615454
rect 253968 615134 254288 615218
rect 253968 614898 254010 615134
rect 254246 614898 254288 615134
rect 253968 614866 254288 614898
rect 284688 615454 285008 615486
rect 284688 615218 284730 615454
rect 284966 615218 285008 615454
rect 284688 615134 285008 615218
rect 284688 614898 284730 615134
rect 284966 614898 285008 615134
rect 284688 614866 285008 614898
rect 315408 615454 315728 615486
rect 315408 615218 315450 615454
rect 315686 615218 315728 615454
rect 315408 615134 315728 615218
rect 315408 614898 315450 615134
rect 315686 614898 315728 615134
rect 315408 614866 315728 614898
rect 346128 615454 346448 615486
rect 346128 615218 346170 615454
rect 346406 615218 346448 615454
rect 346128 615134 346448 615218
rect 346128 614898 346170 615134
rect 346406 614898 346448 615134
rect 346128 614866 346448 614898
rect 376848 615454 377168 615486
rect 376848 615218 376890 615454
rect 377126 615218 377168 615454
rect 376848 615134 377168 615218
rect 376848 614898 376890 615134
rect 377126 614898 377168 615134
rect 376848 614866 377168 614898
rect 407568 615454 407888 615486
rect 407568 615218 407610 615454
rect 407846 615218 407888 615454
rect 407568 615134 407888 615218
rect 407568 614898 407610 615134
rect 407846 614898 407888 615134
rect 407568 614866 407888 614898
rect 438288 615454 438608 615486
rect 438288 615218 438330 615454
rect 438566 615218 438608 615454
rect 438288 615134 438608 615218
rect 438288 614898 438330 615134
rect 438566 614898 438608 615134
rect 438288 614866 438608 614898
rect 469008 615454 469328 615486
rect 469008 615218 469050 615454
rect 469286 615218 469328 615454
rect 469008 615134 469328 615218
rect 469008 614898 469050 615134
rect 469286 614898 469328 615134
rect 469008 614866 469328 614898
rect 499728 615454 500048 615486
rect 499728 615218 499770 615454
rect 500006 615218 500048 615454
rect 499728 615134 500048 615218
rect 499728 614898 499770 615134
rect 500006 614898 500048 615134
rect 499728 614866 500048 614898
rect 530448 615454 530768 615486
rect 530448 615218 530490 615454
rect 530726 615218 530768 615454
rect 530448 615134 530768 615218
rect 530448 614898 530490 615134
rect 530726 614898 530768 615134
rect 530448 614866 530768 614898
rect 561168 615454 561488 615486
rect 561168 615218 561210 615454
rect 561446 615218 561488 615454
rect 561168 615134 561488 615218
rect 561168 614898 561210 615134
rect 561446 614898 561488 615134
rect 561168 614866 561488 614898
rect 567234 604894 567854 640338
rect 567234 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 567854 604894
rect 567234 604574 567854 604658
rect 567234 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 567854 604574
rect 23568 597454 23888 597486
rect 23568 597218 23610 597454
rect 23846 597218 23888 597454
rect 23568 597134 23888 597218
rect 23568 596898 23610 597134
rect 23846 596898 23888 597134
rect 23568 596866 23888 596898
rect 54288 597454 54608 597486
rect 54288 597218 54330 597454
rect 54566 597218 54608 597454
rect 54288 597134 54608 597218
rect 54288 596898 54330 597134
rect 54566 596898 54608 597134
rect 54288 596866 54608 596898
rect 85008 597454 85328 597486
rect 85008 597218 85050 597454
rect 85286 597218 85328 597454
rect 85008 597134 85328 597218
rect 85008 596898 85050 597134
rect 85286 596898 85328 597134
rect 85008 596866 85328 596898
rect 115728 597454 116048 597486
rect 115728 597218 115770 597454
rect 116006 597218 116048 597454
rect 115728 597134 116048 597218
rect 115728 596898 115770 597134
rect 116006 596898 116048 597134
rect 115728 596866 116048 596898
rect 146448 597454 146768 597486
rect 146448 597218 146490 597454
rect 146726 597218 146768 597454
rect 146448 597134 146768 597218
rect 146448 596898 146490 597134
rect 146726 596898 146768 597134
rect 146448 596866 146768 596898
rect 177168 597454 177488 597486
rect 177168 597218 177210 597454
rect 177446 597218 177488 597454
rect 177168 597134 177488 597218
rect 177168 596898 177210 597134
rect 177446 596898 177488 597134
rect 177168 596866 177488 596898
rect 207888 597454 208208 597486
rect 207888 597218 207930 597454
rect 208166 597218 208208 597454
rect 207888 597134 208208 597218
rect 207888 596898 207930 597134
rect 208166 596898 208208 597134
rect 207888 596866 208208 596898
rect 238608 597454 238928 597486
rect 238608 597218 238650 597454
rect 238886 597218 238928 597454
rect 238608 597134 238928 597218
rect 238608 596898 238650 597134
rect 238886 596898 238928 597134
rect 238608 596866 238928 596898
rect 269328 597454 269648 597486
rect 269328 597218 269370 597454
rect 269606 597218 269648 597454
rect 269328 597134 269648 597218
rect 269328 596898 269370 597134
rect 269606 596898 269648 597134
rect 269328 596866 269648 596898
rect 300048 597454 300368 597486
rect 300048 597218 300090 597454
rect 300326 597218 300368 597454
rect 300048 597134 300368 597218
rect 300048 596898 300090 597134
rect 300326 596898 300368 597134
rect 300048 596866 300368 596898
rect 330768 597454 331088 597486
rect 330768 597218 330810 597454
rect 331046 597218 331088 597454
rect 330768 597134 331088 597218
rect 330768 596898 330810 597134
rect 331046 596898 331088 597134
rect 330768 596866 331088 596898
rect 361488 597454 361808 597486
rect 361488 597218 361530 597454
rect 361766 597218 361808 597454
rect 361488 597134 361808 597218
rect 361488 596898 361530 597134
rect 361766 596898 361808 597134
rect 361488 596866 361808 596898
rect 392208 597454 392528 597486
rect 392208 597218 392250 597454
rect 392486 597218 392528 597454
rect 392208 597134 392528 597218
rect 392208 596898 392250 597134
rect 392486 596898 392528 597134
rect 392208 596866 392528 596898
rect 422928 597454 423248 597486
rect 422928 597218 422970 597454
rect 423206 597218 423248 597454
rect 422928 597134 423248 597218
rect 422928 596898 422970 597134
rect 423206 596898 423248 597134
rect 422928 596866 423248 596898
rect 453648 597454 453968 597486
rect 453648 597218 453690 597454
rect 453926 597218 453968 597454
rect 453648 597134 453968 597218
rect 453648 596898 453690 597134
rect 453926 596898 453968 597134
rect 453648 596866 453968 596898
rect 484368 597454 484688 597486
rect 484368 597218 484410 597454
rect 484646 597218 484688 597454
rect 484368 597134 484688 597218
rect 484368 596898 484410 597134
rect 484646 596898 484688 597134
rect 484368 596866 484688 596898
rect 515088 597454 515408 597486
rect 515088 597218 515130 597454
rect 515366 597218 515408 597454
rect 515088 597134 515408 597218
rect 515088 596898 515130 597134
rect 515366 596898 515408 597134
rect 515088 596866 515408 596898
rect 545808 597454 546128 597486
rect 545808 597218 545850 597454
rect 546086 597218 546128 597454
rect 545808 597134 546128 597218
rect 545808 596898 545850 597134
rect 546086 596898 546128 597134
rect 545808 596866 546128 596898
rect -2006 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 -1386 579454
rect -2006 579134 -1386 579218
rect -2006 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 -1386 579134
rect -2006 543454 -1386 578898
rect 8208 579454 8528 579486
rect 8208 579218 8250 579454
rect 8486 579218 8528 579454
rect 8208 579134 8528 579218
rect 8208 578898 8250 579134
rect 8486 578898 8528 579134
rect 8208 578866 8528 578898
rect 38928 579454 39248 579486
rect 38928 579218 38970 579454
rect 39206 579218 39248 579454
rect 38928 579134 39248 579218
rect 38928 578898 38970 579134
rect 39206 578898 39248 579134
rect 38928 578866 39248 578898
rect 69648 579454 69968 579486
rect 69648 579218 69690 579454
rect 69926 579218 69968 579454
rect 69648 579134 69968 579218
rect 69648 578898 69690 579134
rect 69926 578898 69968 579134
rect 69648 578866 69968 578898
rect 100368 579454 100688 579486
rect 100368 579218 100410 579454
rect 100646 579218 100688 579454
rect 100368 579134 100688 579218
rect 100368 578898 100410 579134
rect 100646 578898 100688 579134
rect 100368 578866 100688 578898
rect 131088 579454 131408 579486
rect 131088 579218 131130 579454
rect 131366 579218 131408 579454
rect 131088 579134 131408 579218
rect 131088 578898 131130 579134
rect 131366 578898 131408 579134
rect 131088 578866 131408 578898
rect 161808 579454 162128 579486
rect 161808 579218 161850 579454
rect 162086 579218 162128 579454
rect 161808 579134 162128 579218
rect 161808 578898 161850 579134
rect 162086 578898 162128 579134
rect 161808 578866 162128 578898
rect 192528 579454 192848 579486
rect 192528 579218 192570 579454
rect 192806 579218 192848 579454
rect 192528 579134 192848 579218
rect 192528 578898 192570 579134
rect 192806 578898 192848 579134
rect 192528 578866 192848 578898
rect 223248 579454 223568 579486
rect 223248 579218 223290 579454
rect 223526 579218 223568 579454
rect 223248 579134 223568 579218
rect 223248 578898 223290 579134
rect 223526 578898 223568 579134
rect 223248 578866 223568 578898
rect 253968 579454 254288 579486
rect 253968 579218 254010 579454
rect 254246 579218 254288 579454
rect 253968 579134 254288 579218
rect 253968 578898 254010 579134
rect 254246 578898 254288 579134
rect 253968 578866 254288 578898
rect 284688 579454 285008 579486
rect 284688 579218 284730 579454
rect 284966 579218 285008 579454
rect 284688 579134 285008 579218
rect 284688 578898 284730 579134
rect 284966 578898 285008 579134
rect 284688 578866 285008 578898
rect 315408 579454 315728 579486
rect 315408 579218 315450 579454
rect 315686 579218 315728 579454
rect 315408 579134 315728 579218
rect 315408 578898 315450 579134
rect 315686 578898 315728 579134
rect 315408 578866 315728 578898
rect 346128 579454 346448 579486
rect 346128 579218 346170 579454
rect 346406 579218 346448 579454
rect 346128 579134 346448 579218
rect 346128 578898 346170 579134
rect 346406 578898 346448 579134
rect 346128 578866 346448 578898
rect 376848 579454 377168 579486
rect 376848 579218 376890 579454
rect 377126 579218 377168 579454
rect 376848 579134 377168 579218
rect 376848 578898 376890 579134
rect 377126 578898 377168 579134
rect 376848 578866 377168 578898
rect 407568 579454 407888 579486
rect 407568 579218 407610 579454
rect 407846 579218 407888 579454
rect 407568 579134 407888 579218
rect 407568 578898 407610 579134
rect 407846 578898 407888 579134
rect 407568 578866 407888 578898
rect 438288 579454 438608 579486
rect 438288 579218 438330 579454
rect 438566 579218 438608 579454
rect 438288 579134 438608 579218
rect 438288 578898 438330 579134
rect 438566 578898 438608 579134
rect 438288 578866 438608 578898
rect 469008 579454 469328 579486
rect 469008 579218 469050 579454
rect 469286 579218 469328 579454
rect 469008 579134 469328 579218
rect 469008 578898 469050 579134
rect 469286 578898 469328 579134
rect 469008 578866 469328 578898
rect 499728 579454 500048 579486
rect 499728 579218 499770 579454
rect 500006 579218 500048 579454
rect 499728 579134 500048 579218
rect 499728 578898 499770 579134
rect 500006 578898 500048 579134
rect 499728 578866 500048 578898
rect 530448 579454 530768 579486
rect 530448 579218 530490 579454
rect 530726 579218 530768 579454
rect 530448 579134 530768 579218
rect 530448 578898 530490 579134
rect 530726 578898 530768 579134
rect 530448 578866 530768 578898
rect 561168 579454 561488 579486
rect 561168 579218 561210 579454
rect 561446 579218 561488 579454
rect 561168 579134 561488 579218
rect 561168 578898 561210 579134
rect 561446 578898 561488 579134
rect 561168 578866 561488 578898
rect 567234 568894 567854 604338
rect 567234 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 567854 568894
rect 567234 568574 567854 568658
rect 567234 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 567854 568574
rect 23568 561454 23888 561486
rect 23568 561218 23610 561454
rect 23846 561218 23888 561454
rect 23568 561134 23888 561218
rect 23568 560898 23610 561134
rect 23846 560898 23888 561134
rect 23568 560866 23888 560898
rect 54288 561454 54608 561486
rect 54288 561218 54330 561454
rect 54566 561218 54608 561454
rect 54288 561134 54608 561218
rect 54288 560898 54330 561134
rect 54566 560898 54608 561134
rect 54288 560866 54608 560898
rect 85008 561454 85328 561486
rect 85008 561218 85050 561454
rect 85286 561218 85328 561454
rect 85008 561134 85328 561218
rect 85008 560898 85050 561134
rect 85286 560898 85328 561134
rect 85008 560866 85328 560898
rect 115728 561454 116048 561486
rect 115728 561218 115770 561454
rect 116006 561218 116048 561454
rect 115728 561134 116048 561218
rect 115728 560898 115770 561134
rect 116006 560898 116048 561134
rect 115728 560866 116048 560898
rect 146448 561454 146768 561486
rect 146448 561218 146490 561454
rect 146726 561218 146768 561454
rect 146448 561134 146768 561218
rect 146448 560898 146490 561134
rect 146726 560898 146768 561134
rect 146448 560866 146768 560898
rect 177168 561454 177488 561486
rect 177168 561218 177210 561454
rect 177446 561218 177488 561454
rect 177168 561134 177488 561218
rect 177168 560898 177210 561134
rect 177446 560898 177488 561134
rect 177168 560866 177488 560898
rect 207888 561454 208208 561486
rect 207888 561218 207930 561454
rect 208166 561218 208208 561454
rect 207888 561134 208208 561218
rect 207888 560898 207930 561134
rect 208166 560898 208208 561134
rect 207888 560866 208208 560898
rect 238608 561454 238928 561486
rect 238608 561218 238650 561454
rect 238886 561218 238928 561454
rect 238608 561134 238928 561218
rect 238608 560898 238650 561134
rect 238886 560898 238928 561134
rect 238608 560866 238928 560898
rect 269328 561454 269648 561486
rect 269328 561218 269370 561454
rect 269606 561218 269648 561454
rect 269328 561134 269648 561218
rect 269328 560898 269370 561134
rect 269606 560898 269648 561134
rect 269328 560866 269648 560898
rect 300048 561454 300368 561486
rect 300048 561218 300090 561454
rect 300326 561218 300368 561454
rect 300048 561134 300368 561218
rect 300048 560898 300090 561134
rect 300326 560898 300368 561134
rect 300048 560866 300368 560898
rect 330768 561454 331088 561486
rect 330768 561218 330810 561454
rect 331046 561218 331088 561454
rect 330768 561134 331088 561218
rect 330768 560898 330810 561134
rect 331046 560898 331088 561134
rect 330768 560866 331088 560898
rect 361488 561454 361808 561486
rect 361488 561218 361530 561454
rect 361766 561218 361808 561454
rect 361488 561134 361808 561218
rect 361488 560898 361530 561134
rect 361766 560898 361808 561134
rect 361488 560866 361808 560898
rect 392208 561454 392528 561486
rect 392208 561218 392250 561454
rect 392486 561218 392528 561454
rect 392208 561134 392528 561218
rect 392208 560898 392250 561134
rect 392486 560898 392528 561134
rect 392208 560866 392528 560898
rect 422928 561454 423248 561486
rect 422928 561218 422970 561454
rect 423206 561218 423248 561454
rect 422928 561134 423248 561218
rect 422928 560898 422970 561134
rect 423206 560898 423248 561134
rect 422928 560866 423248 560898
rect 453648 561454 453968 561486
rect 453648 561218 453690 561454
rect 453926 561218 453968 561454
rect 453648 561134 453968 561218
rect 453648 560898 453690 561134
rect 453926 560898 453968 561134
rect 453648 560866 453968 560898
rect 484368 561454 484688 561486
rect 484368 561218 484410 561454
rect 484646 561218 484688 561454
rect 484368 561134 484688 561218
rect 484368 560898 484410 561134
rect 484646 560898 484688 561134
rect 484368 560866 484688 560898
rect 515088 561454 515408 561486
rect 515088 561218 515130 561454
rect 515366 561218 515408 561454
rect 515088 561134 515408 561218
rect 515088 560898 515130 561134
rect 515366 560898 515408 561134
rect 515088 560866 515408 560898
rect 545808 561454 546128 561486
rect 545808 561218 545850 561454
rect 546086 561218 546128 561454
rect 545808 561134 546128 561218
rect 545808 560898 545850 561134
rect 546086 560898 546128 561134
rect 545808 560866 546128 560898
rect -2006 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 -1386 543454
rect -2006 543134 -1386 543218
rect -2006 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 -1386 543134
rect -2006 507454 -1386 542898
rect 8208 543454 8528 543486
rect 8208 543218 8250 543454
rect 8486 543218 8528 543454
rect 8208 543134 8528 543218
rect 8208 542898 8250 543134
rect 8486 542898 8528 543134
rect 8208 542866 8528 542898
rect 38928 543454 39248 543486
rect 38928 543218 38970 543454
rect 39206 543218 39248 543454
rect 38928 543134 39248 543218
rect 38928 542898 38970 543134
rect 39206 542898 39248 543134
rect 38928 542866 39248 542898
rect 69648 543454 69968 543486
rect 69648 543218 69690 543454
rect 69926 543218 69968 543454
rect 69648 543134 69968 543218
rect 69648 542898 69690 543134
rect 69926 542898 69968 543134
rect 69648 542866 69968 542898
rect 100368 543454 100688 543486
rect 100368 543218 100410 543454
rect 100646 543218 100688 543454
rect 100368 543134 100688 543218
rect 100368 542898 100410 543134
rect 100646 542898 100688 543134
rect 100368 542866 100688 542898
rect 131088 543454 131408 543486
rect 131088 543218 131130 543454
rect 131366 543218 131408 543454
rect 131088 543134 131408 543218
rect 131088 542898 131130 543134
rect 131366 542898 131408 543134
rect 131088 542866 131408 542898
rect 161808 543454 162128 543486
rect 161808 543218 161850 543454
rect 162086 543218 162128 543454
rect 161808 543134 162128 543218
rect 161808 542898 161850 543134
rect 162086 542898 162128 543134
rect 161808 542866 162128 542898
rect 192528 543454 192848 543486
rect 192528 543218 192570 543454
rect 192806 543218 192848 543454
rect 192528 543134 192848 543218
rect 192528 542898 192570 543134
rect 192806 542898 192848 543134
rect 192528 542866 192848 542898
rect 223248 543454 223568 543486
rect 223248 543218 223290 543454
rect 223526 543218 223568 543454
rect 223248 543134 223568 543218
rect 223248 542898 223290 543134
rect 223526 542898 223568 543134
rect 223248 542866 223568 542898
rect 253968 543454 254288 543486
rect 253968 543218 254010 543454
rect 254246 543218 254288 543454
rect 253968 543134 254288 543218
rect 253968 542898 254010 543134
rect 254246 542898 254288 543134
rect 253968 542866 254288 542898
rect 284688 543454 285008 543486
rect 284688 543218 284730 543454
rect 284966 543218 285008 543454
rect 284688 543134 285008 543218
rect 284688 542898 284730 543134
rect 284966 542898 285008 543134
rect 284688 542866 285008 542898
rect 315408 543454 315728 543486
rect 315408 543218 315450 543454
rect 315686 543218 315728 543454
rect 315408 543134 315728 543218
rect 315408 542898 315450 543134
rect 315686 542898 315728 543134
rect 315408 542866 315728 542898
rect 346128 543454 346448 543486
rect 346128 543218 346170 543454
rect 346406 543218 346448 543454
rect 346128 543134 346448 543218
rect 346128 542898 346170 543134
rect 346406 542898 346448 543134
rect 346128 542866 346448 542898
rect 376848 543454 377168 543486
rect 376848 543218 376890 543454
rect 377126 543218 377168 543454
rect 376848 543134 377168 543218
rect 376848 542898 376890 543134
rect 377126 542898 377168 543134
rect 376848 542866 377168 542898
rect 407568 543454 407888 543486
rect 407568 543218 407610 543454
rect 407846 543218 407888 543454
rect 407568 543134 407888 543218
rect 407568 542898 407610 543134
rect 407846 542898 407888 543134
rect 407568 542866 407888 542898
rect 438288 543454 438608 543486
rect 438288 543218 438330 543454
rect 438566 543218 438608 543454
rect 438288 543134 438608 543218
rect 438288 542898 438330 543134
rect 438566 542898 438608 543134
rect 438288 542866 438608 542898
rect 469008 543454 469328 543486
rect 469008 543218 469050 543454
rect 469286 543218 469328 543454
rect 469008 543134 469328 543218
rect 469008 542898 469050 543134
rect 469286 542898 469328 543134
rect 469008 542866 469328 542898
rect 499728 543454 500048 543486
rect 499728 543218 499770 543454
rect 500006 543218 500048 543454
rect 499728 543134 500048 543218
rect 499728 542898 499770 543134
rect 500006 542898 500048 543134
rect 499728 542866 500048 542898
rect 530448 543454 530768 543486
rect 530448 543218 530490 543454
rect 530726 543218 530768 543454
rect 530448 543134 530768 543218
rect 530448 542898 530490 543134
rect 530726 542898 530768 543134
rect 530448 542866 530768 542898
rect 561168 543454 561488 543486
rect 561168 543218 561210 543454
rect 561446 543218 561488 543454
rect 561168 543134 561488 543218
rect 561168 542898 561210 543134
rect 561446 542898 561488 543134
rect 561168 542866 561488 542898
rect 567234 532894 567854 568338
rect 567234 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 567854 532894
rect 567234 532574 567854 532658
rect 567234 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 567854 532574
rect 23568 525454 23888 525486
rect 23568 525218 23610 525454
rect 23846 525218 23888 525454
rect 23568 525134 23888 525218
rect 23568 524898 23610 525134
rect 23846 524898 23888 525134
rect 23568 524866 23888 524898
rect 54288 525454 54608 525486
rect 54288 525218 54330 525454
rect 54566 525218 54608 525454
rect 54288 525134 54608 525218
rect 54288 524898 54330 525134
rect 54566 524898 54608 525134
rect 54288 524866 54608 524898
rect 85008 525454 85328 525486
rect 85008 525218 85050 525454
rect 85286 525218 85328 525454
rect 85008 525134 85328 525218
rect 85008 524898 85050 525134
rect 85286 524898 85328 525134
rect 85008 524866 85328 524898
rect 115728 525454 116048 525486
rect 115728 525218 115770 525454
rect 116006 525218 116048 525454
rect 115728 525134 116048 525218
rect 115728 524898 115770 525134
rect 116006 524898 116048 525134
rect 115728 524866 116048 524898
rect 146448 525454 146768 525486
rect 146448 525218 146490 525454
rect 146726 525218 146768 525454
rect 146448 525134 146768 525218
rect 146448 524898 146490 525134
rect 146726 524898 146768 525134
rect 146448 524866 146768 524898
rect 177168 525454 177488 525486
rect 177168 525218 177210 525454
rect 177446 525218 177488 525454
rect 177168 525134 177488 525218
rect 177168 524898 177210 525134
rect 177446 524898 177488 525134
rect 177168 524866 177488 524898
rect 207888 525454 208208 525486
rect 207888 525218 207930 525454
rect 208166 525218 208208 525454
rect 207888 525134 208208 525218
rect 207888 524898 207930 525134
rect 208166 524898 208208 525134
rect 207888 524866 208208 524898
rect 238608 525454 238928 525486
rect 238608 525218 238650 525454
rect 238886 525218 238928 525454
rect 238608 525134 238928 525218
rect 238608 524898 238650 525134
rect 238886 524898 238928 525134
rect 238608 524866 238928 524898
rect 269328 525454 269648 525486
rect 269328 525218 269370 525454
rect 269606 525218 269648 525454
rect 269328 525134 269648 525218
rect 269328 524898 269370 525134
rect 269606 524898 269648 525134
rect 269328 524866 269648 524898
rect 300048 525454 300368 525486
rect 300048 525218 300090 525454
rect 300326 525218 300368 525454
rect 300048 525134 300368 525218
rect 300048 524898 300090 525134
rect 300326 524898 300368 525134
rect 300048 524866 300368 524898
rect 330768 525454 331088 525486
rect 330768 525218 330810 525454
rect 331046 525218 331088 525454
rect 330768 525134 331088 525218
rect 330768 524898 330810 525134
rect 331046 524898 331088 525134
rect 330768 524866 331088 524898
rect 361488 525454 361808 525486
rect 361488 525218 361530 525454
rect 361766 525218 361808 525454
rect 361488 525134 361808 525218
rect 361488 524898 361530 525134
rect 361766 524898 361808 525134
rect 361488 524866 361808 524898
rect 392208 525454 392528 525486
rect 392208 525218 392250 525454
rect 392486 525218 392528 525454
rect 392208 525134 392528 525218
rect 392208 524898 392250 525134
rect 392486 524898 392528 525134
rect 392208 524866 392528 524898
rect 422928 525454 423248 525486
rect 422928 525218 422970 525454
rect 423206 525218 423248 525454
rect 422928 525134 423248 525218
rect 422928 524898 422970 525134
rect 423206 524898 423248 525134
rect 422928 524866 423248 524898
rect 453648 525454 453968 525486
rect 453648 525218 453690 525454
rect 453926 525218 453968 525454
rect 453648 525134 453968 525218
rect 453648 524898 453690 525134
rect 453926 524898 453968 525134
rect 453648 524866 453968 524898
rect 484368 525454 484688 525486
rect 484368 525218 484410 525454
rect 484646 525218 484688 525454
rect 484368 525134 484688 525218
rect 484368 524898 484410 525134
rect 484646 524898 484688 525134
rect 484368 524866 484688 524898
rect 515088 525454 515408 525486
rect 515088 525218 515130 525454
rect 515366 525218 515408 525454
rect 515088 525134 515408 525218
rect 515088 524898 515130 525134
rect 515366 524898 515408 525134
rect 515088 524866 515408 524898
rect 545808 525454 546128 525486
rect 545808 525218 545850 525454
rect 546086 525218 546128 525454
rect 545808 525134 546128 525218
rect 545808 524898 545850 525134
rect 546086 524898 546128 525134
rect 545808 524866 546128 524898
rect -2006 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 -1386 507454
rect -2006 507134 -1386 507218
rect -2006 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 -1386 507134
rect -2006 471454 -1386 506898
rect 8208 507454 8528 507486
rect 8208 507218 8250 507454
rect 8486 507218 8528 507454
rect 8208 507134 8528 507218
rect 8208 506898 8250 507134
rect 8486 506898 8528 507134
rect 8208 506866 8528 506898
rect 38928 507454 39248 507486
rect 38928 507218 38970 507454
rect 39206 507218 39248 507454
rect 38928 507134 39248 507218
rect 38928 506898 38970 507134
rect 39206 506898 39248 507134
rect 38928 506866 39248 506898
rect 69648 507454 69968 507486
rect 69648 507218 69690 507454
rect 69926 507218 69968 507454
rect 69648 507134 69968 507218
rect 69648 506898 69690 507134
rect 69926 506898 69968 507134
rect 69648 506866 69968 506898
rect 100368 507454 100688 507486
rect 100368 507218 100410 507454
rect 100646 507218 100688 507454
rect 100368 507134 100688 507218
rect 100368 506898 100410 507134
rect 100646 506898 100688 507134
rect 100368 506866 100688 506898
rect 131088 507454 131408 507486
rect 131088 507218 131130 507454
rect 131366 507218 131408 507454
rect 131088 507134 131408 507218
rect 131088 506898 131130 507134
rect 131366 506898 131408 507134
rect 131088 506866 131408 506898
rect 161808 507454 162128 507486
rect 161808 507218 161850 507454
rect 162086 507218 162128 507454
rect 161808 507134 162128 507218
rect 161808 506898 161850 507134
rect 162086 506898 162128 507134
rect 161808 506866 162128 506898
rect 192528 507454 192848 507486
rect 192528 507218 192570 507454
rect 192806 507218 192848 507454
rect 192528 507134 192848 507218
rect 192528 506898 192570 507134
rect 192806 506898 192848 507134
rect 192528 506866 192848 506898
rect 223248 507454 223568 507486
rect 223248 507218 223290 507454
rect 223526 507218 223568 507454
rect 223248 507134 223568 507218
rect 223248 506898 223290 507134
rect 223526 506898 223568 507134
rect 223248 506866 223568 506898
rect 253968 507454 254288 507486
rect 253968 507218 254010 507454
rect 254246 507218 254288 507454
rect 253968 507134 254288 507218
rect 253968 506898 254010 507134
rect 254246 506898 254288 507134
rect 253968 506866 254288 506898
rect 284688 507454 285008 507486
rect 284688 507218 284730 507454
rect 284966 507218 285008 507454
rect 284688 507134 285008 507218
rect 284688 506898 284730 507134
rect 284966 506898 285008 507134
rect 284688 506866 285008 506898
rect 315408 507454 315728 507486
rect 315408 507218 315450 507454
rect 315686 507218 315728 507454
rect 315408 507134 315728 507218
rect 315408 506898 315450 507134
rect 315686 506898 315728 507134
rect 315408 506866 315728 506898
rect 346128 507454 346448 507486
rect 346128 507218 346170 507454
rect 346406 507218 346448 507454
rect 346128 507134 346448 507218
rect 346128 506898 346170 507134
rect 346406 506898 346448 507134
rect 346128 506866 346448 506898
rect 376848 507454 377168 507486
rect 376848 507218 376890 507454
rect 377126 507218 377168 507454
rect 376848 507134 377168 507218
rect 376848 506898 376890 507134
rect 377126 506898 377168 507134
rect 376848 506866 377168 506898
rect 407568 507454 407888 507486
rect 407568 507218 407610 507454
rect 407846 507218 407888 507454
rect 407568 507134 407888 507218
rect 407568 506898 407610 507134
rect 407846 506898 407888 507134
rect 407568 506866 407888 506898
rect 438288 507454 438608 507486
rect 438288 507218 438330 507454
rect 438566 507218 438608 507454
rect 438288 507134 438608 507218
rect 438288 506898 438330 507134
rect 438566 506898 438608 507134
rect 438288 506866 438608 506898
rect 469008 507454 469328 507486
rect 469008 507218 469050 507454
rect 469286 507218 469328 507454
rect 469008 507134 469328 507218
rect 469008 506898 469050 507134
rect 469286 506898 469328 507134
rect 469008 506866 469328 506898
rect 499728 507454 500048 507486
rect 499728 507218 499770 507454
rect 500006 507218 500048 507454
rect 499728 507134 500048 507218
rect 499728 506898 499770 507134
rect 500006 506898 500048 507134
rect 499728 506866 500048 506898
rect 530448 507454 530768 507486
rect 530448 507218 530490 507454
rect 530726 507218 530768 507454
rect 530448 507134 530768 507218
rect 530448 506898 530490 507134
rect 530726 506898 530768 507134
rect 530448 506866 530768 506898
rect 561168 507454 561488 507486
rect 561168 507218 561210 507454
rect 561446 507218 561488 507454
rect 561168 507134 561488 507218
rect 561168 506898 561210 507134
rect 561446 506898 561488 507134
rect 561168 506866 561488 506898
rect 567234 496894 567854 532338
rect 567234 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 567854 496894
rect 567234 496574 567854 496658
rect 567234 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 567854 496574
rect 23568 489454 23888 489486
rect 23568 489218 23610 489454
rect 23846 489218 23888 489454
rect 23568 489134 23888 489218
rect 23568 488898 23610 489134
rect 23846 488898 23888 489134
rect 23568 488866 23888 488898
rect 54288 489454 54608 489486
rect 54288 489218 54330 489454
rect 54566 489218 54608 489454
rect 54288 489134 54608 489218
rect 54288 488898 54330 489134
rect 54566 488898 54608 489134
rect 54288 488866 54608 488898
rect 85008 489454 85328 489486
rect 85008 489218 85050 489454
rect 85286 489218 85328 489454
rect 85008 489134 85328 489218
rect 85008 488898 85050 489134
rect 85286 488898 85328 489134
rect 85008 488866 85328 488898
rect 115728 489454 116048 489486
rect 115728 489218 115770 489454
rect 116006 489218 116048 489454
rect 115728 489134 116048 489218
rect 115728 488898 115770 489134
rect 116006 488898 116048 489134
rect 115728 488866 116048 488898
rect 146448 489454 146768 489486
rect 146448 489218 146490 489454
rect 146726 489218 146768 489454
rect 146448 489134 146768 489218
rect 146448 488898 146490 489134
rect 146726 488898 146768 489134
rect 146448 488866 146768 488898
rect 177168 489454 177488 489486
rect 177168 489218 177210 489454
rect 177446 489218 177488 489454
rect 177168 489134 177488 489218
rect 177168 488898 177210 489134
rect 177446 488898 177488 489134
rect 177168 488866 177488 488898
rect 207888 489454 208208 489486
rect 207888 489218 207930 489454
rect 208166 489218 208208 489454
rect 207888 489134 208208 489218
rect 207888 488898 207930 489134
rect 208166 488898 208208 489134
rect 207888 488866 208208 488898
rect 238608 489454 238928 489486
rect 238608 489218 238650 489454
rect 238886 489218 238928 489454
rect 238608 489134 238928 489218
rect 238608 488898 238650 489134
rect 238886 488898 238928 489134
rect 238608 488866 238928 488898
rect 269328 489454 269648 489486
rect 269328 489218 269370 489454
rect 269606 489218 269648 489454
rect 269328 489134 269648 489218
rect 269328 488898 269370 489134
rect 269606 488898 269648 489134
rect 269328 488866 269648 488898
rect 300048 489454 300368 489486
rect 300048 489218 300090 489454
rect 300326 489218 300368 489454
rect 300048 489134 300368 489218
rect 300048 488898 300090 489134
rect 300326 488898 300368 489134
rect 300048 488866 300368 488898
rect 330768 489454 331088 489486
rect 330768 489218 330810 489454
rect 331046 489218 331088 489454
rect 330768 489134 331088 489218
rect 330768 488898 330810 489134
rect 331046 488898 331088 489134
rect 330768 488866 331088 488898
rect 361488 489454 361808 489486
rect 361488 489218 361530 489454
rect 361766 489218 361808 489454
rect 361488 489134 361808 489218
rect 361488 488898 361530 489134
rect 361766 488898 361808 489134
rect 361488 488866 361808 488898
rect 392208 489454 392528 489486
rect 392208 489218 392250 489454
rect 392486 489218 392528 489454
rect 392208 489134 392528 489218
rect 392208 488898 392250 489134
rect 392486 488898 392528 489134
rect 392208 488866 392528 488898
rect 422928 489454 423248 489486
rect 422928 489218 422970 489454
rect 423206 489218 423248 489454
rect 422928 489134 423248 489218
rect 422928 488898 422970 489134
rect 423206 488898 423248 489134
rect 422928 488866 423248 488898
rect 453648 489454 453968 489486
rect 453648 489218 453690 489454
rect 453926 489218 453968 489454
rect 453648 489134 453968 489218
rect 453648 488898 453690 489134
rect 453926 488898 453968 489134
rect 453648 488866 453968 488898
rect 484368 489454 484688 489486
rect 484368 489218 484410 489454
rect 484646 489218 484688 489454
rect 484368 489134 484688 489218
rect 484368 488898 484410 489134
rect 484646 488898 484688 489134
rect 484368 488866 484688 488898
rect 515088 489454 515408 489486
rect 515088 489218 515130 489454
rect 515366 489218 515408 489454
rect 515088 489134 515408 489218
rect 515088 488898 515130 489134
rect 515366 488898 515408 489134
rect 515088 488866 515408 488898
rect 545808 489454 546128 489486
rect 545808 489218 545850 489454
rect 546086 489218 546128 489454
rect 545808 489134 546128 489218
rect 545808 488898 545850 489134
rect 546086 488898 546128 489134
rect 545808 488866 546128 488898
rect -2006 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 -1386 471454
rect -2006 471134 -1386 471218
rect -2006 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 -1386 471134
rect -2006 435454 -1386 470898
rect 8208 471454 8528 471486
rect 8208 471218 8250 471454
rect 8486 471218 8528 471454
rect 8208 471134 8528 471218
rect 8208 470898 8250 471134
rect 8486 470898 8528 471134
rect 8208 470866 8528 470898
rect 38928 471454 39248 471486
rect 38928 471218 38970 471454
rect 39206 471218 39248 471454
rect 38928 471134 39248 471218
rect 38928 470898 38970 471134
rect 39206 470898 39248 471134
rect 38928 470866 39248 470898
rect 69648 471454 69968 471486
rect 69648 471218 69690 471454
rect 69926 471218 69968 471454
rect 69648 471134 69968 471218
rect 69648 470898 69690 471134
rect 69926 470898 69968 471134
rect 69648 470866 69968 470898
rect 100368 471454 100688 471486
rect 100368 471218 100410 471454
rect 100646 471218 100688 471454
rect 100368 471134 100688 471218
rect 100368 470898 100410 471134
rect 100646 470898 100688 471134
rect 100368 470866 100688 470898
rect 131088 471454 131408 471486
rect 131088 471218 131130 471454
rect 131366 471218 131408 471454
rect 131088 471134 131408 471218
rect 131088 470898 131130 471134
rect 131366 470898 131408 471134
rect 131088 470866 131408 470898
rect 161808 471454 162128 471486
rect 161808 471218 161850 471454
rect 162086 471218 162128 471454
rect 161808 471134 162128 471218
rect 161808 470898 161850 471134
rect 162086 470898 162128 471134
rect 161808 470866 162128 470898
rect 192528 471454 192848 471486
rect 192528 471218 192570 471454
rect 192806 471218 192848 471454
rect 192528 471134 192848 471218
rect 192528 470898 192570 471134
rect 192806 470898 192848 471134
rect 192528 470866 192848 470898
rect 223248 471454 223568 471486
rect 223248 471218 223290 471454
rect 223526 471218 223568 471454
rect 223248 471134 223568 471218
rect 223248 470898 223290 471134
rect 223526 470898 223568 471134
rect 223248 470866 223568 470898
rect 253968 471454 254288 471486
rect 253968 471218 254010 471454
rect 254246 471218 254288 471454
rect 253968 471134 254288 471218
rect 253968 470898 254010 471134
rect 254246 470898 254288 471134
rect 253968 470866 254288 470898
rect 284688 471454 285008 471486
rect 284688 471218 284730 471454
rect 284966 471218 285008 471454
rect 284688 471134 285008 471218
rect 284688 470898 284730 471134
rect 284966 470898 285008 471134
rect 284688 470866 285008 470898
rect 315408 471454 315728 471486
rect 315408 471218 315450 471454
rect 315686 471218 315728 471454
rect 315408 471134 315728 471218
rect 315408 470898 315450 471134
rect 315686 470898 315728 471134
rect 315408 470866 315728 470898
rect 346128 471454 346448 471486
rect 346128 471218 346170 471454
rect 346406 471218 346448 471454
rect 346128 471134 346448 471218
rect 346128 470898 346170 471134
rect 346406 470898 346448 471134
rect 346128 470866 346448 470898
rect 376848 471454 377168 471486
rect 376848 471218 376890 471454
rect 377126 471218 377168 471454
rect 376848 471134 377168 471218
rect 376848 470898 376890 471134
rect 377126 470898 377168 471134
rect 376848 470866 377168 470898
rect 407568 471454 407888 471486
rect 407568 471218 407610 471454
rect 407846 471218 407888 471454
rect 407568 471134 407888 471218
rect 407568 470898 407610 471134
rect 407846 470898 407888 471134
rect 407568 470866 407888 470898
rect 438288 471454 438608 471486
rect 438288 471218 438330 471454
rect 438566 471218 438608 471454
rect 438288 471134 438608 471218
rect 438288 470898 438330 471134
rect 438566 470898 438608 471134
rect 438288 470866 438608 470898
rect 469008 471454 469328 471486
rect 469008 471218 469050 471454
rect 469286 471218 469328 471454
rect 469008 471134 469328 471218
rect 469008 470898 469050 471134
rect 469286 470898 469328 471134
rect 469008 470866 469328 470898
rect 499728 471454 500048 471486
rect 499728 471218 499770 471454
rect 500006 471218 500048 471454
rect 499728 471134 500048 471218
rect 499728 470898 499770 471134
rect 500006 470898 500048 471134
rect 499728 470866 500048 470898
rect 530448 471454 530768 471486
rect 530448 471218 530490 471454
rect 530726 471218 530768 471454
rect 530448 471134 530768 471218
rect 530448 470898 530490 471134
rect 530726 470898 530768 471134
rect 530448 470866 530768 470898
rect 561168 471454 561488 471486
rect 561168 471218 561210 471454
rect 561446 471218 561488 471454
rect 561168 471134 561488 471218
rect 561168 470898 561210 471134
rect 561446 470898 561488 471134
rect 561168 470866 561488 470898
rect 567234 460894 567854 496338
rect 567234 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 567854 460894
rect 567234 460574 567854 460658
rect 567234 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 567854 460574
rect 23568 453454 23888 453486
rect 23568 453218 23610 453454
rect 23846 453218 23888 453454
rect 23568 453134 23888 453218
rect 23568 452898 23610 453134
rect 23846 452898 23888 453134
rect 23568 452866 23888 452898
rect 54288 453454 54608 453486
rect 54288 453218 54330 453454
rect 54566 453218 54608 453454
rect 54288 453134 54608 453218
rect 54288 452898 54330 453134
rect 54566 452898 54608 453134
rect 54288 452866 54608 452898
rect 85008 453454 85328 453486
rect 85008 453218 85050 453454
rect 85286 453218 85328 453454
rect 85008 453134 85328 453218
rect 85008 452898 85050 453134
rect 85286 452898 85328 453134
rect 85008 452866 85328 452898
rect 115728 453454 116048 453486
rect 115728 453218 115770 453454
rect 116006 453218 116048 453454
rect 115728 453134 116048 453218
rect 115728 452898 115770 453134
rect 116006 452898 116048 453134
rect 115728 452866 116048 452898
rect 146448 453454 146768 453486
rect 146448 453218 146490 453454
rect 146726 453218 146768 453454
rect 146448 453134 146768 453218
rect 146448 452898 146490 453134
rect 146726 452898 146768 453134
rect 146448 452866 146768 452898
rect 177168 453454 177488 453486
rect 177168 453218 177210 453454
rect 177446 453218 177488 453454
rect 177168 453134 177488 453218
rect 177168 452898 177210 453134
rect 177446 452898 177488 453134
rect 177168 452866 177488 452898
rect 207888 453454 208208 453486
rect 207888 453218 207930 453454
rect 208166 453218 208208 453454
rect 207888 453134 208208 453218
rect 207888 452898 207930 453134
rect 208166 452898 208208 453134
rect 207888 452866 208208 452898
rect 238608 453454 238928 453486
rect 238608 453218 238650 453454
rect 238886 453218 238928 453454
rect 238608 453134 238928 453218
rect 238608 452898 238650 453134
rect 238886 452898 238928 453134
rect 238608 452866 238928 452898
rect 269328 453454 269648 453486
rect 269328 453218 269370 453454
rect 269606 453218 269648 453454
rect 269328 453134 269648 453218
rect 269328 452898 269370 453134
rect 269606 452898 269648 453134
rect 269328 452866 269648 452898
rect 300048 453454 300368 453486
rect 300048 453218 300090 453454
rect 300326 453218 300368 453454
rect 300048 453134 300368 453218
rect 300048 452898 300090 453134
rect 300326 452898 300368 453134
rect 300048 452866 300368 452898
rect 330768 453454 331088 453486
rect 330768 453218 330810 453454
rect 331046 453218 331088 453454
rect 330768 453134 331088 453218
rect 330768 452898 330810 453134
rect 331046 452898 331088 453134
rect 330768 452866 331088 452898
rect 361488 453454 361808 453486
rect 361488 453218 361530 453454
rect 361766 453218 361808 453454
rect 361488 453134 361808 453218
rect 361488 452898 361530 453134
rect 361766 452898 361808 453134
rect 361488 452866 361808 452898
rect 392208 453454 392528 453486
rect 392208 453218 392250 453454
rect 392486 453218 392528 453454
rect 392208 453134 392528 453218
rect 392208 452898 392250 453134
rect 392486 452898 392528 453134
rect 392208 452866 392528 452898
rect 422928 453454 423248 453486
rect 422928 453218 422970 453454
rect 423206 453218 423248 453454
rect 422928 453134 423248 453218
rect 422928 452898 422970 453134
rect 423206 452898 423248 453134
rect 422928 452866 423248 452898
rect 453648 453454 453968 453486
rect 453648 453218 453690 453454
rect 453926 453218 453968 453454
rect 453648 453134 453968 453218
rect 453648 452898 453690 453134
rect 453926 452898 453968 453134
rect 453648 452866 453968 452898
rect 484368 453454 484688 453486
rect 484368 453218 484410 453454
rect 484646 453218 484688 453454
rect 484368 453134 484688 453218
rect 484368 452898 484410 453134
rect 484646 452898 484688 453134
rect 484368 452866 484688 452898
rect 515088 453454 515408 453486
rect 515088 453218 515130 453454
rect 515366 453218 515408 453454
rect 515088 453134 515408 453218
rect 515088 452898 515130 453134
rect 515366 452898 515408 453134
rect 515088 452866 515408 452898
rect 545808 453454 546128 453486
rect 545808 453218 545850 453454
rect 546086 453218 546128 453454
rect 545808 453134 546128 453218
rect 545808 452898 545850 453134
rect 546086 452898 546128 453134
rect 545808 452866 546128 452898
rect -2006 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 -1386 435454
rect -2006 435134 -1386 435218
rect -2006 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 -1386 435134
rect -2006 399454 -1386 434898
rect 8208 435454 8528 435486
rect 8208 435218 8250 435454
rect 8486 435218 8528 435454
rect 8208 435134 8528 435218
rect 8208 434898 8250 435134
rect 8486 434898 8528 435134
rect 8208 434866 8528 434898
rect 38928 435454 39248 435486
rect 38928 435218 38970 435454
rect 39206 435218 39248 435454
rect 38928 435134 39248 435218
rect 38928 434898 38970 435134
rect 39206 434898 39248 435134
rect 38928 434866 39248 434898
rect 69648 435454 69968 435486
rect 69648 435218 69690 435454
rect 69926 435218 69968 435454
rect 69648 435134 69968 435218
rect 69648 434898 69690 435134
rect 69926 434898 69968 435134
rect 69648 434866 69968 434898
rect 100368 435454 100688 435486
rect 100368 435218 100410 435454
rect 100646 435218 100688 435454
rect 100368 435134 100688 435218
rect 100368 434898 100410 435134
rect 100646 434898 100688 435134
rect 100368 434866 100688 434898
rect 131088 435454 131408 435486
rect 131088 435218 131130 435454
rect 131366 435218 131408 435454
rect 131088 435134 131408 435218
rect 131088 434898 131130 435134
rect 131366 434898 131408 435134
rect 131088 434866 131408 434898
rect 161808 435454 162128 435486
rect 161808 435218 161850 435454
rect 162086 435218 162128 435454
rect 161808 435134 162128 435218
rect 161808 434898 161850 435134
rect 162086 434898 162128 435134
rect 161808 434866 162128 434898
rect 192528 435454 192848 435486
rect 192528 435218 192570 435454
rect 192806 435218 192848 435454
rect 192528 435134 192848 435218
rect 192528 434898 192570 435134
rect 192806 434898 192848 435134
rect 192528 434866 192848 434898
rect 223248 435454 223568 435486
rect 223248 435218 223290 435454
rect 223526 435218 223568 435454
rect 223248 435134 223568 435218
rect 223248 434898 223290 435134
rect 223526 434898 223568 435134
rect 223248 434866 223568 434898
rect 253968 435454 254288 435486
rect 253968 435218 254010 435454
rect 254246 435218 254288 435454
rect 253968 435134 254288 435218
rect 253968 434898 254010 435134
rect 254246 434898 254288 435134
rect 253968 434866 254288 434898
rect 284688 435454 285008 435486
rect 284688 435218 284730 435454
rect 284966 435218 285008 435454
rect 284688 435134 285008 435218
rect 284688 434898 284730 435134
rect 284966 434898 285008 435134
rect 284688 434866 285008 434898
rect 315408 435454 315728 435486
rect 315408 435218 315450 435454
rect 315686 435218 315728 435454
rect 315408 435134 315728 435218
rect 315408 434898 315450 435134
rect 315686 434898 315728 435134
rect 315408 434866 315728 434898
rect 346128 435454 346448 435486
rect 346128 435218 346170 435454
rect 346406 435218 346448 435454
rect 346128 435134 346448 435218
rect 346128 434898 346170 435134
rect 346406 434898 346448 435134
rect 346128 434866 346448 434898
rect 376848 435454 377168 435486
rect 376848 435218 376890 435454
rect 377126 435218 377168 435454
rect 376848 435134 377168 435218
rect 376848 434898 376890 435134
rect 377126 434898 377168 435134
rect 376848 434866 377168 434898
rect 407568 435454 407888 435486
rect 407568 435218 407610 435454
rect 407846 435218 407888 435454
rect 407568 435134 407888 435218
rect 407568 434898 407610 435134
rect 407846 434898 407888 435134
rect 407568 434866 407888 434898
rect 438288 435454 438608 435486
rect 438288 435218 438330 435454
rect 438566 435218 438608 435454
rect 438288 435134 438608 435218
rect 438288 434898 438330 435134
rect 438566 434898 438608 435134
rect 438288 434866 438608 434898
rect 469008 435454 469328 435486
rect 469008 435218 469050 435454
rect 469286 435218 469328 435454
rect 469008 435134 469328 435218
rect 469008 434898 469050 435134
rect 469286 434898 469328 435134
rect 469008 434866 469328 434898
rect 499728 435454 500048 435486
rect 499728 435218 499770 435454
rect 500006 435218 500048 435454
rect 499728 435134 500048 435218
rect 499728 434898 499770 435134
rect 500006 434898 500048 435134
rect 499728 434866 500048 434898
rect 530448 435454 530768 435486
rect 530448 435218 530490 435454
rect 530726 435218 530768 435454
rect 530448 435134 530768 435218
rect 530448 434898 530490 435134
rect 530726 434898 530768 435134
rect 530448 434866 530768 434898
rect 561168 435454 561488 435486
rect 561168 435218 561210 435454
rect 561446 435218 561488 435454
rect 561168 435134 561488 435218
rect 561168 434898 561210 435134
rect 561446 434898 561488 435134
rect 561168 434866 561488 434898
rect 567234 424894 567854 460338
rect 567234 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 567854 424894
rect 567234 424574 567854 424658
rect 567234 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 567854 424574
rect 23568 417454 23888 417486
rect 23568 417218 23610 417454
rect 23846 417218 23888 417454
rect 23568 417134 23888 417218
rect 23568 416898 23610 417134
rect 23846 416898 23888 417134
rect 23568 416866 23888 416898
rect 54288 417454 54608 417486
rect 54288 417218 54330 417454
rect 54566 417218 54608 417454
rect 54288 417134 54608 417218
rect 54288 416898 54330 417134
rect 54566 416898 54608 417134
rect 54288 416866 54608 416898
rect 85008 417454 85328 417486
rect 85008 417218 85050 417454
rect 85286 417218 85328 417454
rect 85008 417134 85328 417218
rect 85008 416898 85050 417134
rect 85286 416898 85328 417134
rect 85008 416866 85328 416898
rect 115728 417454 116048 417486
rect 115728 417218 115770 417454
rect 116006 417218 116048 417454
rect 115728 417134 116048 417218
rect 115728 416898 115770 417134
rect 116006 416898 116048 417134
rect 115728 416866 116048 416898
rect 146448 417454 146768 417486
rect 146448 417218 146490 417454
rect 146726 417218 146768 417454
rect 146448 417134 146768 417218
rect 146448 416898 146490 417134
rect 146726 416898 146768 417134
rect 146448 416866 146768 416898
rect 177168 417454 177488 417486
rect 177168 417218 177210 417454
rect 177446 417218 177488 417454
rect 177168 417134 177488 417218
rect 177168 416898 177210 417134
rect 177446 416898 177488 417134
rect 177168 416866 177488 416898
rect 207888 417454 208208 417486
rect 207888 417218 207930 417454
rect 208166 417218 208208 417454
rect 207888 417134 208208 417218
rect 207888 416898 207930 417134
rect 208166 416898 208208 417134
rect 207888 416866 208208 416898
rect 238608 417454 238928 417486
rect 238608 417218 238650 417454
rect 238886 417218 238928 417454
rect 238608 417134 238928 417218
rect 238608 416898 238650 417134
rect 238886 416898 238928 417134
rect 238608 416866 238928 416898
rect 269328 417454 269648 417486
rect 269328 417218 269370 417454
rect 269606 417218 269648 417454
rect 269328 417134 269648 417218
rect 269328 416898 269370 417134
rect 269606 416898 269648 417134
rect 269328 416866 269648 416898
rect 300048 417454 300368 417486
rect 300048 417218 300090 417454
rect 300326 417218 300368 417454
rect 300048 417134 300368 417218
rect 300048 416898 300090 417134
rect 300326 416898 300368 417134
rect 300048 416866 300368 416898
rect 330768 417454 331088 417486
rect 330768 417218 330810 417454
rect 331046 417218 331088 417454
rect 330768 417134 331088 417218
rect 330768 416898 330810 417134
rect 331046 416898 331088 417134
rect 330768 416866 331088 416898
rect 361488 417454 361808 417486
rect 361488 417218 361530 417454
rect 361766 417218 361808 417454
rect 361488 417134 361808 417218
rect 361488 416898 361530 417134
rect 361766 416898 361808 417134
rect 361488 416866 361808 416898
rect 392208 417454 392528 417486
rect 392208 417218 392250 417454
rect 392486 417218 392528 417454
rect 392208 417134 392528 417218
rect 392208 416898 392250 417134
rect 392486 416898 392528 417134
rect 392208 416866 392528 416898
rect 422928 417454 423248 417486
rect 422928 417218 422970 417454
rect 423206 417218 423248 417454
rect 422928 417134 423248 417218
rect 422928 416898 422970 417134
rect 423206 416898 423248 417134
rect 422928 416866 423248 416898
rect 453648 417454 453968 417486
rect 453648 417218 453690 417454
rect 453926 417218 453968 417454
rect 453648 417134 453968 417218
rect 453648 416898 453690 417134
rect 453926 416898 453968 417134
rect 453648 416866 453968 416898
rect 484368 417454 484688 417486
rect 484368 417218 484410 417454
rect 484646 417218 484688 417454
rect 484368 417134 484688 417218
rect 484368 416898 484410 417134
rect 484646 416898 484688 417134
rect 484368 416866 484688 416898
rect 515088 417454 515408 417486
rect 515088 417218 515130 417454
rect 515366 417218 515408 417454
rect 515088 417134 515408 417218
rect 515088 416898 515130 417134
rect 515366 416898 515408 417134
rect 515088 416866 515408 416898
rect 545808 417454 546128 417486
rect 545808 417218 545850 417454
rect 546086 417218 546128 417454
rect 545808 417134 546128 417218
rect 545808 416898 545850 417134
rect 546086 416898 546128 417134
rect 545808 416866 546128 416898
rect -2006 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 -1386 399454
rect -2006 399134 -1386 399218
rect -2006 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 -1386 399134
rect -2006 363454 -1386 398898
rect 8208 399454 8528 399486
rect 8208 399218 8250 399454
rect 8486 399218 8528 399454
rect 8208 399134 8528 399218
rect 8208 398898 8250 399134
rect 8486 398898 8528 399134
rect 8208 398866 8528 398898
rect 38928 399454 39248 399486
rect 38928 399218 38970 399454
rect 39206 399218 39248 399454
rect 38928 399134 39248 399218
rect 38928 398898 38970 399134
rect 39206 398898 39248 399134
rect 38928 398866 39248 398898
rect 69648 399454 69968 399486
rect 69648 399218 69690 399454
rect 69926 399218 69968 399454
rect 69648 399134 69968 399218
rect 69648 398898 69690 399134
rect 69926 398898 69968 399134
rect 69648 398866 69968 398898
rect 100368 399454 100688 399486
rect 100368 399218 100410 399454
rect 100646 399218 100688 399454
rect 100368 399134 100688 399218
rect 100368 398898 100410 399134
rect 100646 398898 100688 399134
rect 100368 398866 100688 398898
rect 131088 399454 131408 399486
rect 131088 399218 131130 399454
rect 131366 399218 131408 399454
rect 131088 399134 131408 399218
rect 131088 398898 131130 399134
rect 131366 398898 131408 399134
rect 131088 398866 131408 398898
rect 161808 399454 162128 399486
rect 161808 399218 161850 399454
rect 162086 399218 162128 399454
rect 161808 399134 162128 399218
rect 161808 398898 161850 399134
rect 162086 398898 162128 399134
rect 161808 398866 162128 398898
rect 192528 399454 192848 399486
rect 192528 399218 192570 399454
rect 192806 399218 192848 399454
rect 192528 399134 192848 399218
rect 192528 398898 192570 399134
rect 192806 398898 192848 399134
rect 192528 398866 192848 398898
rect 223248 399454 223568 399486
rect 223248 399218 223290 399454
rect 223526 399218 223568 399454
rect 223248 399134 223568 399218
rect 223248 398898 223290 399134
rect 223526 398898 223568 399134
rect 223248 398866 223568 398898
rect 253968 399454 254288 399486
rect 253968 399218 254010 399454
rect 254246 399218 254288 399454
rect 253968 399134 254288 399218
rect 253968 398898 254010 399134
rect 254246 398898 254288 399134
rect 253968 398866 254288 398898
rect 284688 399454 285008 399486
rect 284688 399218 284730 399454
rect 284966 399218 285008 399454
rect 284688 399134 285008 399218
rect 284688 398898 284730 399134
rect 284966 398898 285008 399134
rect 284688 398866 285008 398898
rect 315408 399454 315728 399486
rect 315408 399218 315450 399454
rect 315686 399218 315728 399454
rect 315408 399134 315728 399218
rect 315408 398898 315450 399134
rect 315686 398898 315728 399134
rect 315408 398866 315728 398898
rect 346128 399454 346448 399486
rect 346128 399218 346170 399454
rect 346406 399218 346448 399454
rect 346128 399134 346448 399218
rect 346128 398898 346170 399134
rect 346406 398898 346448 399134
rect 346128 398866 346448 398898
rect 376848 399454 377168 399486
rect 376848 399218 376890 399454
rect 377126 399218 377168 399454
rect 376848 399134 377168 399218
rect 376848 398898 376890 399134
rect 377126 398898 377168 399134
rect 376848 398866 377168 398898
rect 407568 399454 407888 399486
rect 407568 399218 407610 399454
rect 407846 399218 407888 399454
rect 407568 399134 407888 399218
rect 407568 398898 407610 399134
rect 407846 398898 407888 399134
rect 407568 398866 407888 398898
rect 438288 399454 438608 399486
rect 438288 399218 438330 399454
rect 438566 399218 438608 399454
rect 438288 399134 438608 399218
rect 438288 398898 438330 399134
rect 438566 398898 438608 399134
rect 438288 398866 438608 398898
rect 469008 399454 469328 399486
rect 469008 399218 469050 399454
rect 469286 399218 469328 399454
rect 469008 399134 469328 399218
rect 469008 398898 469050 399134
rect 469286 398898 469328 399134
rect 469008 398866 469328 398898
rect 499728 399454 500048 399486
rect 499728 399218 499770 399454
rect 500006 399218 500048 399454
rect 499728 399134 500048 399218
rect 499728 398898 499770 399134
rect 500006 398898 500048 399134
rect 499728 398866 500048 398898
rect 530448 399454 530768 399486
rect 530448 399218 530490 399454
rect 530726 399218 530768 399454
rect 530448 399134 530768 399218
rect 530448 398898 530490 399134
rect 530726 398898 530768 399134
rect 530448 398866 530768 398898
rect 561168 399454 561488 399486
rect 561168 399218 561210 399454
rect 561446 399218 561488 399454
rect 561168 399134 561488 399218
rect 561168 398898 561210 399134
rect 561446 398898 561488 399134
rect 561168 398866 561488 398898
rect 567234 388894 567854 424338
rect 567234 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 567854 388894
rect 567234 388574 567854 388658
rect 567234 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 567854 388574
rect 23568 381454 23888 381486
rect 23568 381218 23610 381454
rect 23846 381218 23888 381454
rect 23568 381134 23888 381218
rect 23568 380898 23610 381134
rect 23846 380898 23888 381134
rect 23568 380866 23888 380898
rect 54288 381454 54608 381486
rect 54288 381218 54330 381454
rect 54566 381218 54608 381454
rect 54288 381134 54608 381218
rect 54288 380898 54330 381134
rect 54566 380898 54608 381134
rect 54288 380866 54608 380898
rect 85008 381454 85328 381486
rect 85008 381218 85050 381454
rect 85286 381218 85328 381454
rect 85008 381134 85328 381218
rect 85008 380898 85050 381134
rect 85286 380898 85328 381134
rect 85008 380866 85328 380898
rect 115728 381454 116048 381486
rect 115728 381218 115770 381454
rect 116006 381218 116048 381454
rect 115728 381134 116048 381218
rect 115728 380898 115770 381134
rect 116006 380898 116048 381134
rect 115728 380866 116048 380898
rect 146448 381454 146768 381486
rect 146448 381218 146490 381454
rect 146726 381218 146768 381454
rect 146448 381134 146768 381218
rect 146448 380898 146490 381134
rect 146726 380898 146768 381134
rect 146448 380866 146768 380898
rect 177168 381454 177488 381486
rect 177168 381218 177210 381454
rect 177446 381218 177488 381454
rect 177168 381134 177488 381218
rect 177168 380898 177210 381134
rect 177446 380898 177488 381134
rect 177168 380866 177488 380898
rect 207888 381454 208208 381486
rect 207888 381218 207930 381454
rect 208166 381218 208208 381454
rect 207888 381134 208208 381218
rect 207888 380898 207930 381134
rect 208166 380898 208208 381134
rect 207888 380866 208208 380898
rect 238608 381454 238928 381486
rect 238608 381218 238650 381454
rect 238886 381218 238928 381454
rect 238608 381134 238928 381218
rect 238608 380898 238650 381134
rect 238886 380898 238928 381134
rect 238608 380866 238928 380898
rect 269328 381454 269648 381486
rect 269328 381218 269370 381454
rect 269606 381218 269648 381454
rect 269328 381134 269648 381218
rect 269328 380898 269370 381134
rect 269606 380898 269648 381134
rect 269328 380866 269648 380898
rect 300048 381454 300368 381486
rect 300048 381218 300090 381454
rect 300326 381218 300368 381454
rect 300048 381134 300368 381218
rect 300048 380898 300090 381134
rect 300326 380898 300368 381134
rect 300048 380866 300368 380898
rect 330768 381454 331088 381486
rect 330768 381218 330810 381454
rect 331046 381218 331088 381454
rect 330768 381134 331088 381218
rect 330768 380898 330810 381134
rect 331046 380898 331088 381134
rect 330768 380866 331088 380898
rect 361488 381454 361808 381486
rect 361488 381218 361530 381454
rect 361766 381218 361808 381454
rect 361488 381134 361808 381218
rect 361488 380898 361530 381134
rect 361766 380898 361808 381134
rect 361488 380866 361808 380898
rect 392208 381454 392528 381486
rect 392208 381218 392250 381454
rect 392486 381218 392528 381454
rect 392208 381134 392528 381218
rect 392208 380898 392250 381134
rect 392486 380898 392528 381134
rect 392208 380866 392528 380898
rect 422928 381454 423248 381486
rect 422928 381218 422970 381454
rect 423206 381218 423248 381454
rect 422928 381134 423248 381218
rect 422928 380898 422970 381134
rect 423206 380898 423248 381134
rect 422928 380866 423248 380898
rect 453648 381454 453968 381486
rect 453648 381218 453690 381454
rect 453926 381218 453968 381454
rect 453648 381134 453968 381218
rect 453648 380898 453690 381134
rect 453926 380898 453968 381134
rect 453648 380866 453968 380898
rect 484368 381454 484688 381486
rect 484368 381218 484410 381454
rect 484646 381218 484688 381454
rect 484368 381134 484688 381218
rect 484368 380898 484410 381134
rect 484646 380898 484688 381134
rect 484368 380866 484688 380898
rect 515088 381454 515408 381486
rect 515088 381218 515130 381454
rect 515366 381218 515408 381454
rect 515088 381134 515408 381218
rect 515088 380898 515130 381134
rect 515366 380898 515408 381134
rect 515088 380866 515408 380898
rect 545808 381454 546128 381486
rect 545808 381218 545850 381454
rect 546086 381218 546128 381454
rect 545808 381134 546128 381218
rect 545808 380898 545850 381134
rect 546086 380898 546128 381134
rect 545808 380866 546128 380898
rect -2006 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 -1386 363454
rect -2006 363134 -1386 363218
rect -2006 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 -1386 363134
rect -2006 327454 -1386 362898
rect 8208 363454 8528 363486
rect 8208 363218 8250 363454
rect 8486 363218 8528 363454
rect 8208 363134 8528 363218
rect 8208 362898 8250 363134
rect 8486 362898 8528 363134
rect 8208 362866 8528 362898
rect 38928 363454 39248 363486
rect 38928 363218 38970 363454
rect 39206 363218 39248 363454
rect 38928 363134 39248 363218
rect 38928 362898 38970 363134
rect 39206 362898 39248 363134
rect 38928 362866 39248 362898
rect 69648 363454 69968 363486
rect 69648 363218 69690 363454
rect 69926 363218 69968 363454
rect 69648 363134 69968 363218
rect 69648 362898 69690 363134
rect 69926 362898 69968 363134
rect 69648 362866 69968 362898
rect 100368 363454 100688 363486
rect 100368 363218 100410 363454
rect 100646 363218 100688 363454
rect 100368 363134 100688 363218
rect 100368 362898 100410 363134
rect 100646 362898 100688 363134
rect 100368 362866 100688 362898
rect 131088 363454 131408 363486
rect 131088 363218 131130 363454
rect 131366 363218 131408 363454
rect 131088 363134 131408 363218
rect 131088 362898 131130 363134
rect 131366 362898 131408 363134
rect 131088 362866 131408 362898
rect 161808 363454 162128 363486
rect 161808 363218 161850 363454
rect 162086 363218 162128 363454
rect 161808 363134 162128 363218
rect 161808 362898 161850 363134
rect 162086 362898 162128 363134
rect 161808 362866 162128 362898
rect 192528 363454 192848 363486
rect 192528 363218 192570 363454
rect 192806 363218 192848 363454
rect 192528 363134 192848 363218
rect 192528 362898 192570 363134
rect 192806 362898 192848 363134
rect 192528 362866 192848 362898
rect 223248 363454 223568 363486
rect 223248 363218 223290 363454
rect 223526 363218 223568 363454
rect 223248 363134 223568 363218
rect 223248 362898 223290 363134
rect 223526 362898 223568 363134
rect 223248 362866 223568 362898
rect 253968 363454 254288 363486
rect 253968 363218 254010 363454
rect 254246 363218 254288 363454
rect 253968 363134 254288 363218
rect 253968 362898 254010 363134
rect 254246 362898 254288 363134
rect 253968 362866 254288 362898
rect 284688 363454 285008 363486
rect 284688 363218 284730 363454
rect 284966 363218 285008 363454
rect 284688 363134 285008 363218
rect 284688 362898 284730 363134
rect 284966 362898 285008 363134
rect 284688 362866 285008 362898
rect 315408 363454 315728 363486
rect 315408 363218 315450 363454
rect 315686 363218 315728 363454
rect 315408 363134 315728 363218
rect 315408 362898 315450 363134
rect 315686 362898 315728 363134
rect 315408 362866 315728 362898
rect 346128 363454 346448 363486
rect 346128 363218 346170 363454
rect 346406 363218 346448 363454
rect 346128 363134 346448 363218
rect 346128 362898 346170 363134
rect 346406 362898 346448 363134
rect 346128 362866 346448 362898
rect 376848 363454 377168 363486
rect 376848 363218 376890 363454
rect 377126 363218 377168 363454
rect 376848 363134 377168 363218
rect 376848 362898 376890 363134
rect 377126 362898 377168 363134
rect 376848 362866 377168 362898
rect 407568 363454 407888 363486
rect 407568 363218 407610 363454
rect 407846 363218 407888 363454
rect 407568 363134 407888 363218
rect 407568 362898 407610 363134
rect 407846 362898 407888 363134
rect 407568 362866 407888 362898
rect 438288 363454 438608 363486
rect 438288 363218 438330 363454
rect 438566 363218 438608 363454
rect 438288 363134 438608 363218
rect 438288 362898 438330 363134
rect 438566 362898 438608 363134
rect 438288 362866 438608 362898
rect 469008 363454 469328 363486
rect 469008 363218 469050 363454
rect 469286 363218 469328 363454
rect 469008 363134 469328 363218
rect 469008 362898 469050 363134
rect 469286 362898 469328 363134
rect 469008 362866 469328 362898
rect 499728 363454 500048 363486
rect 499728 363218 499770 363454
rect 500006 363218 500048 363454
rect 499728 363134 500048 363218
rect 499728 362898 499770 363134
rect 500006 362898 500048 363134
rect 499728 362866 500048 362898
rect 530448 363454 530768 363486
rect 530448 363218 530490 363454
rect 530726 363218 530768 363454
rect 530448 363134 530768 363218
rect 530448 362898 530490 363134
rect 530726 362898 530768 363134
rect 530448 362866 530768 362898
rect 561168 363454 561488 363486
rect 561168 363218 561210 363454
rect 561446 363218 561488 363454
rect 561168 363134 561488 363218
rect 561168 362898 561210 363134
rect 561446 362898 561488 363134
rect 561168 362866 561488 362898
rect 567234 352894 567854 388338
rect 567234 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 567854 352894
rect 567234 352574 567854 352658
rect 567234 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 567854 352574
rect 23568 345454 23888 345486
rect 23568 345218 23610 345454
rect 23846 345218 23888 345454
rect 23568 345134 23888 345218
rect 23568 344898 23610 345134
rect 23846 344898 23888 345134
rect 23568 344866 23888 344898
rect 54288 345454 54608 345486
rect 54288 345218 54330 345454
rect 54566 345218 54608 345454
rect 54288 345134 54608 345218
rect 54288 344898 54330 345134
rect 54566 344898 54608 345134
rect 54288 344866 54608 344898
rect 85008 345454 85328 345486
rect 85008 345218 85050 345454
rect 85286 345218 85328 345454
rect 85008 345134 85328 345218
rect 85008 344898 85050 345134
rect 85286 344898 85328 345134
rect 85008 344866 85328 344898
rect 115728 345454 116048 345486
rect 115728 345218 115770 345454
rect 116006 345218 116048 345454
rect 115728 345134 116048 345218
rect 115728 344898 115770 345134
rect 116006 344898 116048 345134
rect 115728 344866 116048 344898
rect 146448 345454 146768 345486
rect 146448 345218 146490 345454
rect 146726 345218 146768 345454
rect 146448 345134 146768 345218
rect 146448 344898 146490 345134
rect 146726 344898 146768 345134
rect 146448 344866 146768 344898
rect 177168 345454 177488 345486
rect 177168 345218 177210 345454
rect 177446 345218 177488 345454
rect 177168 345134 177488 345218
rect 177168 344898 177210 345134
rect 177446 344898 177488 345134
rect 177168 344866 177488 344898
rect 207888 345454 208208 345486
rect 207888 345218 207930 345454
rect 208166 345218 208208 345454
rect 207888 345134 208208 345218
rect 207888 344898 207930 345134
rect 208166 344898 208208 345134
rect 207888 344866 208208 344898
rect 238608 345454 238928 345486
rect 238608 345218 238650 345454
rect 238886 345218 238928 345454
rect 238608 345134 238928 345218
rect 238608 344898 238650 345134
rect 238886 344898 238928 345134
rect 238608 344866 238928 344898
rect 269328 345454 269648 345486
rect 269328 345218 269370 345454
rect 269606 345218 269648 345454
rect 269328 345134 269648 345218
rect 269328 344898 269370 345134
rect 269606 344898 269648 345134
rect 269328 344866 269648 344898
rect 300048 345454 300368 345486
rect 300048 345218 300090 345454
rect 300326 345218 300368 345454
rect 300048 345134 300368 345218
rect 300048 344898 300090 345134
rect 300326 344898 300368 345134
rect 300048 344866 300368 344898
rect 330768 345454 331088 345486
rect 330768 345218 330810 345454
rect 331046 345218 331088 345454
rect 330768 345134 331088 345218
rect 330768 344898 330810 345134
rect 331046 344898 331088 345134
rect 330768 344866 331088 344898
rect 361488 345454 361808 345486
rect 361488 345218 361530 345454
rect 361766 345218 361808 345454
rect 361488 345134 361808 345218
rect 361488 344898 361530 345134
rect 361766 344898 361808 345134
rect 361488 344866 361808 344898
rect 392208 345454 392528 345486
rect 392208 345218 392250 345454
rect 392486 345218 392528 345454
rect 392208 345134 392528 345218
rect 392208 344898 392250 345134
rect 392486 344898 392528 345134
rect 392208 344866 392528 344898
rect 422928 345454 423248 345486
rect 422928 345218 422970 345454
rect 423206 345218 423248 345454
rect 422928 345134 423248 345218
rect 422928 344898 422970 345134
rect 423206 344898 423248 345134
rect 422928 344866 423248 344898
rect 453648 345454 453968 345486
rect 453648 345218 453690 345454
rect 453926 345218 453968 345454
rect 453648 345134 453968 345218
rect 453648 344898 453690 345134
rect 453926 344898 453968 345134
rect 453648 344866 453968 344898
rect 484368 345454 484688 345486
rect 484368 345218 484410 345454
rect 484646 345218 484688 345454
rect 484368 345134 484688 345218
rect 484368 344898 484410 345134
rect 484646 344898 484688 345134
rect 484368 344866 484688 344898
rect 515088 345454 515408 345486
rect 515088 345218 515130 345454
rect 515366 345218 515408 345454
rect 515088 345134 515408 345218
rect 515088 344898 515130 345134
rect 515366 344898 515408 345134
rect 515088 344866 515408 344898
rect 545808 345454 546128 345486
rect 545808 345218 545850 345454
rect 546086 345218 546128 345454
rect 545808 345134 546128 345218
rect 545808 344898 545850 345134
rect 546086 344898 546128 345134
rect 545808 344866 546128 344898
rect -2006 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 -1386 327454
rect -2006 327134 -1386 327218
rect -2006 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 -1386 327134
rect -2006 291454 -1386 326898
rect 8208 327454 8528 327486
rect 8208 327218 8250 327454
rect 8486 327218 8528 327454
rect 8208 327134 8528 327218
rect 8208 326898 8250 327134
rect 8486 326898 8528 327134
rect 8208 326866 8528 326898
rect 38928 327454 39248 327486
rect 38928 327218 38970 327454
rect 39206 327218 39248 327454
rect 38928 327134 39248 327218
rect 38928 326898 38970 327134
rect 39206 326898 39248 327134
rect 38928 326866 39248 326898
rect 69648 327454 69968 327486
rect 69648 327218 69690 327454
rect 69926 327218 69968 327454
rect 69648 327134 69968 327218
rect 69648 326898 69690 327134
rect 69926 326898 69968 327134
rect 69648 326866 69968 326898
rect 100368 327454 100688 327486
rect 100368 327218 100410 327454
rect 100646 327218 100688 327454
rect 100368 327134 100688 327218
rect 100368 326898 100410 327134
rect 100646 326898 100688 327134
rect 100368 326866 100688 326898
rect 131088 327454 131408 327486
rect 131088 327218 131130 327454
rect 131366 327218 131408 327454
rect 131088 327134 131408 327218
rect 131088 326898 131130 327134
rect 131366 326898 131408 327134
rect 131088 326866 131408 326898
rect 161808 327454 162128 327486
rect 161808 327218 161850 327454
rect 162086 327218 162128 327454
rect 161808 327134 162128 327218
rect 161808 326898 161850 327134
rect 162086 326898 162128 327134
rect 161808 326866 162128 326898
rect 192528 327454 192848 327486
rect 192528 327218 192570 327454
rect 192806 327218 192848 327454
rect 192528 327134 192848 327218
rect 192528 326898 192570 327134
rect 192806 326898 192848 327134
rect 192528 326866 192848 326898
rect 223248 327454 223568 327486
rect 223248 327218 223290 327454
rect 223526 327218 223568 327454
rect 223248 327134 223568 327218
rect 223248 326898 223290 327134
rect 223526 326898 223568 327134
rect 223248 326866 223568 326898
rect 253968 327454 254288 327486
rect 253968 327218 254010 327454
rect 254246 327218 254288 327454
rect 253968 327134 254288 327218
rect 253968 326898 254010 327134
rect 254246 326898 254288 327134
rect 253968 326866 254288 326898
rect 284688 327454 285008 327486
rect 284688 327218 284730 327454
rect 284966 327218 285008 327454
rect 284688 327134 285008 327218
rect 284688 326898 284730 327134
rect 284966 326898 285008 327134
rect 284688 326866 285008 326898
rect 315408 327454 315728 327486
rect 315408 327218 315450 327454
rect 315686 327218 315728 327454
rect 315408 327134 315728 327218
rect 315408 326898 315450 327134
rect 315686 326898 315728 327134
rect 315408 326866 315728 326898
rect 346128 327454 346448 327486
rect 346128 327218 346170 327454
rect 346406 327218 346448 327454
rect 346128 327134 346448 327218
rect 346128 326898 346170 327134
rect 346406 326898 346448 327134
rect 346128 326866 346448 326898
rect 376848 327454 377168 327486
rect 376848 327218 376890 327454
rect 377126 327218 377168 327454
rect 376848 327134 377168 327218
rect 376848 326898 376890 327134
rect 377126 326898 377168 327134
rect 376848 326866 377168 326898
rect 407568 327454 407888 327486
rect 407568 327218 407610 327454
rect 407846 327218 407888 327454
rect 407568 327134 407888 327218
rect 407568 326898 407610 327134
rect 407846 326898 407888 327134
rect 407568 326866 407888 326898
rect 438288 327454 438608 327486
rect 438288 327218 438330 327454
rect 438566 327218 438608 327454
rect 438288 327134 438608 327218
rect 438288 326898 438330 327134
rect 438566 326898 438608 327134
rect 438288 326866 438608 326898
rect 469008 327454 469328 327486
rect 469008 327218 469050 327454
rect 469286 327218 469328 327454
rect 469008 327134 469328 327218
rect 469008 326898 469050 327134
rect 469286 326898 469328 327134
rect 469008 326866 469328 326898
rect 499728 327454 500048 327486
rect 499728 327218 499770 327454
rect 500006 327218 500048 327454
rect 499728 327134 500048 327218
rect 499728 326898 499770 327134
rect 500006 326898 500048 327134
rect 499728 326866 500048 326898
rect 530448 327454 530768 327486
rect 530448 327218 530490 327454
rect 530726 327218 530768 327454
rect 530448 327134 530768 327218
rect 530448 326898 530490 327134
rect 530726 326898 530768 327134
rect 530448 326866 530768 326898
rect 561168 327454 561488 327486
rect 561168 327218 561210 327454
rect 561446 327218 561488 327454
rect 561168 327134 561488 327218
rect 561168 326898 561210 327134
rect 561446 326898 561488 327134
rect 561168 326866 561488 326898
rect 567234 316894 567854 352338
rect 567234 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 567854 316894
rect 567234 316574 567854 316658
rect 567234 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 567854 316574
rect 23568 309454 23888 309486
rect 23568 309218 23610 309454
rect 23846 309218 23888 309454
rect 23568 309134 23888 309218
rect 23568 308898 23610 309134
rect 23846 308898 23888 309134
rect 23568 308866 23888 308898
rect 54288 309454 54608 309486
rect 54288 309218 54330 309454
rect 54566 309218 54608 309454
rect 54288 309134 54608 309218
rect 54288 308898 54330 309134
rect 54566 308898 54608 309134
rect 54288 308866 54608 308898
rect 85008 309454 85328 309486
rect 85008 309218 85050 309454
rect 85286 309218 85328 309454
rect 85008 309134 85328 309218
rect 85008 308898 85050 309134
rect 85286 308898 85328 309134
rect 85008 308866 85328 308898
rect 115728 309454 116048 309486
rect 115728 309218 115770 309454
rect 116006 309218 116048 309454
rect 115728 309134 116048 309218
rect 115728 308898 115770 309134
rect 116006 308898 116048 309134
rect 115728 308866 116048 308898
rect 146448 309454 146768 309486
rect 146448 309218 146490 309454
rect 146726 309218 146768 309454
rect 146448 309134 146768 309218
rect 146448 308898 146490 309134
rect 146726 308898 146768 309134
rect 146448 308866 146768 308898
rect 177168 309454 177488 309486
rect 177168 309218 177210 309454
rect 177446 309218 177488 309454
rect 177168 309134 177488 309218
rect 177168 308898 177210 309134
rect 177446 308898 177488 309134
rect 177168 308866 177488 308898
rect 207888 309454 208208 309486
rect 207888 309218 207930 309454
rect 208166 309218 208208 309454
rect 207888 309134 208208 309218
rect 207888 308898 207930 309134
rect 208166 308898 208208 309134
rect 207888 308866 208208 308898
rect 238608 309454 238928 309486
rect 238608 309218 238650 309454
rect 238886 309218 238928 309454
rect 238608 309134 238928 309218
rect 238608 308898 238650 309134
rect 238886 308898 238928 309134
rect 238608 308866 238928 308898
rect 269328 309454 269648 309486
rect 269328 309218 269370 309454
rect 269606 309218 269648 309454
rect 269328 309134 269648 309218
rect 269328 308898 269370 309134
rect 269606 308898 269648 309134
rect 269328 308866 269648 308898
rect 300048 309454 300368 309486
rect 300048 309218 300090 309454
rect 300326 309218 300368 309454
rect 300048 309134 300368 309218
rect 300048 308898 300090 309134
rect 300326 308898 300368 309134
rect 300048 308866 300368 308898
rect 330768 309454 331088 309486
rect 330768 309218 330810 309454
rect 331046 309218 331088 309454
rect 330768 309134 331088 309218
rect 330768 308898 330810 309134
rect 331046 308898 331088 309134
rect 330768 308866 331088 308898
rect 361488 309454 361808 309486
rect 361488 309218 361530 309454
rect 361766 309218 361808 309454
rect 361488 309134 361808 309218
rect 361488 308898 361530 309134
rect 361766 308898 361808 309134
rect 361488 308866 361808 308898
rect 392208 309454 392528 309486
rect 392208 309218 392250 309454
rect 392486 309218 392528 309454
rect 392208 309134 392528 309218
rect 392208 308898 392250 309134
rect 392486 308898 392528 309134
rect 392208 308866 392528 308898
rect 422928 309454 423248 309486
rect 422928 309218 422970 309454
rect 423206 309218 423248 309454
rect 422928 309134 423248 309218
rect 422928 308898 422970 309134
rect 423206 308898 423248 309134
rect 422928 308866 423248 308898
rect 453648 309454 453968 309486
rect 453648 309218 453690 309454
rect 453926 309218 453968 309454
rect 453648 309134 453968 309218
rect 453648 308898 453690 309134
rect 453926 308898 453968 309134
rect 453648 308866 453968 308898
rect 484368 309454 484688 309486
rect 484368 309218 484410 309454
rect 484646 309218 484688 309454
rect 484368 309134 484688 309218
rect 484368 308898 484410 309134
rect 484646 308898 484688 309134
rect 484368 308866 484688 308898
rect 515088 309454 515408 309486
rect 515088 309218 515130 309454
rect 515366 309218 515408 309454
rect 515088 309134 515408 309218
rect 515088 308898 515130 309134
rect 515366 308898 515408 309134
rect 515088 308866 515408 308898
rect 545808 309454 546128 309486
rect 545808 309218 545850 309454
rect 546086 309218 546128 309454
rect 545808 309134 546128 309218
rect 545808 308898 545850 309134
rect 546086 308898 546128 309134
rect 545808 308866 546128 308898
rect -2006 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 -1386 291454
rect -2006 291134 -1386 291218
rect -2006 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 -1386 291134
rect -2006 255454 -1386 290898
rect 8208 291454 8528 291486
rect 8208 291218 8250 291454
rect 8486 291218 8528 291454
rect 8208 291134 8528 291218
rect 8208 290898 8250 291134
rect 8486 290898 8528 291134
rect 8208 290866 8528 290898
rect 38928 291454 39248 291486
rect 38928 291218 38970 291454
rect 39206 291218 39248 291454
rect 38928 291134 39248 291218
rect 38928 290898 38970 291134
rect 39206 290898 39248 291134
rect 38928 290866 39248 290898
rect 69648 291454 69968 291486
rect 69648 291218 69690 291454
rect 69926 291218 69968 291454
rect 69648 291134 69968 291218
rect 69648 290898 69690 291134
rect 69926 290898 69968 291134
rect 69648 290866 69968 290898
rect 100368 291454 100688 291486
rect 100368 291218 100410 291454
rect 100646 291218 100688 291454
rect 100368 291134 100688 291218
rect 100368 290898 100410 291134
rect 100646 290898 100688 291134
rect 100368 290866 100688 290898
rect 131088 291454 131408 291486
rect 131088 291218 131130 291454
rect 131366 291218 131408 291454
rect 131088 291134 131408 291218
rect 131088 290898 131130 291134
rect 131366 290898 131408 291134
rect 131088 290866 131408 290898
rect 161808 291454 162128 291486
rect 161808 291218 161850 291454
rect 162086 291218 162128 291454
rect 161808 291134 162128 291218
rect 161808 290898 161850 291134
rect 162086 290898 162128 291134
rect 161808 290866 162128 290898
rect 192528 291454 192848 291486
rect 192528 291218 192570 291454
rect 192806 291218 192848 291454
rect 192528 291134 192848 291218
rect 192528 290898 192570 291134
rect 192806 290898 192848 291134
rect 192528 290866 192848 290898
rect 223248 291454 223568 291486
rect 223248 291218 223290 291454
rect 223526 291218 223568 291454
rect 223248 291134 223568 291218
rect 223248 290898 223290 291134
rect 223526 290898 223568 291134
rect 223248 290866 223568 290898
rect 253968 291454 254288 291486
rect 253968 291218 254010 291454
rect 254246 291218 254288 291454
rect 253968 291134 254288 291218
rect 253968 290898 254010 291134
rect 254246 290898 254288 291134
rect 253968 290866 254288 290898
rect 284688 291454 285008 291486
rect 284688 291218 284730 291454
rect 284966 291218 285008 291454
rect 284688 291134 285008 291218
rect 284688 290898 284730 291134
rect 284966 290898 285008 291134
rect 284688 290866 285008 290898
rect 315408 291454 315728 291486
rect 315408 291218 315450 291454
rect 315686 291218 315728 291454
rect 315408 291134 315728 291218
rect 315408 290898 315450 291134
rect 315686 290898 315728 291134
rect 315408 290866 315728 290898
rect 346128 291454 346448 291486
rect 346128 291218 346170 291454
rect 346406 291218 346448 291454
rect 346128 291134 346448 291218
rect 346128 290898 346170 291134
rect 346406 290898 346448 291134
rect 346128 290866 346448 290898
rect 376848 291454 377168 291486
rect 376848 291218 376890 291454
rect 377126 291218 377168 291454
rect 376848 291134 377168 291218
rect 376848 290898 376890 291134
rect 377126 290898 377168 291134
rect 376848 290866 377168 290898
rect 407568 291454 407888 291486
rect 407568 291218 407610 291454
rect 407846 291218 407888 291454
rect 407568 291134 407888 291218
rect 407568 290898 407610 291134
rect 407846 290898 407888 291134
rect 407568 290866 407888 290898
rect 438288 291454 438608 291486
rect 438288 291218 438330 291454
rect 438566 291218 438608 291454
rect 438288 291134 438608 291218
rect 438288 290898 438330 291134
rect 438566 290898 438608 291134
rect 438288 290866 438608 290898
rect 469008 291454 469328 291486
rect 469008 291218 469050 291454
rect 469286 291218 469328 291454
rect 469008 291134 469328 291218
rect 469008 290898 469050 291134
rect 469286 290898 469328 291134
rect 469008 290866 469328 290898
rect 499728 291454 500048 291486
rect 499728 291218 499770 291454
rect 500006 291218 500048 291454
rect 499728 291134 500048 291218
rect 499728 290898 499770 291134
rect 500006 290898 500048 291134
rect 499728 290866 500048 290898
rect 530448 291454 530768 291486
rect 530448 291218 530490 291454
rect 530726 291218 530768 291454
rect 530448 291134 530768 291218
rect 530448 290898 530490 291134
rect 530726 290898 530768 291134
rect 530448 290866 530768 290898
rect 561168 291454 561488 291486
rect 561168 291218 561210 291454
rect 561446 291218 561488 291454
rect 561168 291134 561488 291218
rect 561168 290898 561210 291134
rect 561446 290898 561488 291134
rect 561168 290866 561488 290898
rect 567234 280894 567854 316338
rect 567234 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 567854 280894
rect 567234 280574 567854 280658
rect 567234 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 567854 280574
rect 23568 273454 23888 273486
rect 23568 273218 23610 273454
rect 23846 273218 23888 273454
rect 23568 273134 23888 273218
rect 23568 272898 23610 273134
rect 23846 272898 23888 273134
rect 23568 272866 23888 272898
rect 54288 273454 54608 273486
rect 54288 273218 54330 273454
rect 54566 273218 54608 273454
rect 54288 273134 54608 273218
rect 54288 272898 54330 273134
rect 54566 272898 54608 273134
rect 54288 272866 54608 272898
rect 85008 273454 85328 273486
rect 85008 273218 85050 273454
rect 85286 273218 85328 273454
rect 85008 273134 85328 273218
rect 85008 272898 85050 273134
rect 85286 272898 85328 273134
rect 85008 272866 85328 272898
rect 115728 273454 116048 273486
rect 115728 273218 115770 273454
rect 116006 273218 116048 273454
rect 115728 273134 116048 273218
rect 115728 272898 115770 273134
rect 116006 272898 116048 273134
rect 115728 272866 116048 272898
rect 146448 273454 146768 273486
rect 146448 273218 146490 273454
rect 146726 273218 146768 273454
rect 146448 273134 146768 273218
rect 146448 272898 146490 273134
rect 146726 272898 146768 273134
rect 146448 272866 146768 272898
rect 177168 273454 177488 273486
rect 177168 273218 177210 273454
rect 177446 273218 177488 273454
rect 177168 273134 177488 273218
rect 177168 272898 177210 273134
rect 177446 272898 177488 273134
rect 177168 272866 177488 272898
rect 207888 273454 208208 273486
rect 207888 273218 207930 273454
rect 208166 273218 208208 273454
rect 207888 273134 208208 273218
rect 207888 272898 207930 273134
rect 208166 272898 208208 273134
rect 207888 272866 208208 272898
rect 238608 273454 238928 273486
rect 238608 273218 238650 273454
rect 238886 273218 238928 273454
rect 238608 273134 238928 273218
rect 238608 272898 238650 273134
rect 238886 272898 238928 273134
rect 238608 272866 238928 272898
rect 269328 273454 269648 273486
rect 269328 273218 269370 273454
rect 269606 273218 269648 273454
rect 269328 273134 269648 273218
rect 269328 272898 269370 273134
rect 269606 272898 269648 273134
rect 269328 272866 269648 272898
rect 300048 273454 300368 273486
rect 300048 273218 300090 273454
rect 300326 273218 300368 273454
rect 300048 273134 300368 273218
rect 300048 272898 300090 273134
rect 300326 272898 300368 273134
rect 300048 272866 300368 272898
rect 330768 273454 331088 273486
rect 330768 273218 330810 273454
rect 331046 273218 331088 273454
rect 330768 273134 331088 273218
rect 330768 272898 330810 273134
rect 331046 272898 331088 273134
rect 330768 272866 331088 272898
rect 361488 273454 361808 273486
rect 361488 273218 361530 273454
rect 361766 273218 361808 273454
rect 361488 273134 361808 273218
rect 361488 272898 361530 273134
rect 361766 272898 361808 273134
rect 361488 272866 361808 272898
rect 392208 273454 392528 273486
rect 392208 273218 392250 273454
rect 392486 273218 392528 273454
rect 392208 273134 392528 273218
rect 392208 272898 392250 273134
rect 392486 272898 392528 273134
rect 392208 272866 392528 272898
rect 422928 273454 423248 273486
rect 422928 273218 422970 273454
rect 423206 273218 423248 273454
rect 422928 273134 423248 273218
rect 422928 272898 422970 273134
rect 423206 272898 423248 273134
rect 422928 272866 423248 272898
rect 453648 273454 453968 273486
rect 453648 273218 453690 273454
rect 453926 273218 453968 273454
rect 453648 273134 453968 273218
rect 453648 272898 453690 273134
rect 453926 272898 453968 273134
rect 453648 272866 453968 272898
rect 484368 273454 484688 273486
rect 484368 273218 484410 273454
rect 484646 273218 484688 273454
rect 484368 273134 484688 273218
rect 484368 272898 484410 273134
rect 484646 272898 484688 273134
rect 484368 272866 484688 272898
rect 515088 273454 515408 273486
rect 515088 273218 515130 273454
rect 515366 273218 515408 273454
rect 515088 273134 515408 273218
rect 515088 272898 515130 273134
rect 515366 272898 515408 273134
rect 515088 272866 515408 272898
rect 545808 273454 546128 273486
rect 545808 273218 545850 273454
rect 546086 273218 546128 273454
rect 545808 273134 546128 273218
rect 545808 272898 545850 273134
rect 546086 272898 546128 273134
rect 545808 272866 546128 272898
rect -2006 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 -1386 255454
rect -2006 255134 -1386 255218
rect -2006 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 -1386 255134
rect -2006 219454 -1386 254898
rect 8208 255454 8528 255486
rect 8208 255218 8250 255454
rect 8486 255218 8528 255454
rect 8208 255134 8528 255218
rect 8208 254898 8250 255134
rect 8486 254898 8528 255134
rect 8208 254866 8528 254898
rect 38928 255454 39248 255486
rect 38928 255218 38970 255454
rect 39206 255218 39248 255454
rect 38928 255134 39248 255218
rect 38928 254898 38970 255134
rect 39206 254898 39248 255134
rect 38928 254866 39248 254898
rect 69648 255454 69968 255486
rect 69648 255218 69690 255454
rect 69926 255218 69968 255454
rect 69648 255134 69968 255218
rect 69648 254898 69690 255134
rect 69926 254898 69968 255134
rect 69648 254866 69968 254898
rect 100368 255454 100688 255486
rect 100368 255218 100410 255454
rect 100646 255218 100688 255454
rect 100368 255134 100688 255218
rect 100368 254898 100410 255134
rect 100646 254898 100688 255134
rect 100368 254866 100688 254898
rect 131088 255454 131408 255486
rect 131088 255218 131130 255454
rect 131366 255218 131408 255454
rect 131088 255134 131408 255218
rect 131088 254898 131130 255134
rect 131366 254898 131408 255134
rect 131088 254866 131408 254898
rect 161808 255454 162128 255486
rect 161808 255218 161850 255454
rect 162086 255218 162128 255454
rect 161808 255134 162128 255218
rect 161808 254898 161850 255134
rect 162086 254898 162128 255134
rect 161808 254866 162128 254898
rect 192528 255454 192848 255486
rect 192528 255218 192570 255454
rect 192806 255218 192848 255454
rect 192528 255134 192848 255218
rect 192528 254898 192570 255134
rect 192806 254898 192848 255134
rect 192528 254866 192848 254898
rect 223248 255454 223568 255486
rect 223248 255218 223290 255454
rect 223526 255218 223568 255454
rect 223248 255134 223568 255218
rect 223248 254898 223290 255134
rect 223526 254898 223568 255134
rect 223248 254866 223568 254898
rect 253968 255454 254288 255486
rect 253968 255218 254010 255454
rect 254246 255218 254288 255454
rect 253968 255134 254288 255218
rect 253968 254898 254010 255134
rect 254246 254898 254288 255134
rect 253968 254866 254288 254898
rect 284688 255454 285008 255486
rect 284688 255218 284730 255454
rect 284966 255218 285008 255454
rect 284688 255134 285008 255218
rect 284688 254898 284730 255134
rect 284966 254898 285008 255134
rect 284688 254866 285008 254898
rect 315408 255454 315728 255486
rect 315408 255218 315450 255454
rect 315686 255218 315728 255454
rect 315408 255134 315728 255218
rect 315408 254898 315450 255134
rect 315686 254898 315728 255134
rect 315408 254866 315728 254898
rect 346128 255454 346448 255486
rect 346128 255218 346170 255454
rect 346406 255218 346448 255454
rect 346128 255134 346448 255218
rect 346128 254898 346170 255134
rect 346406 254898 346448 255134
rect 346128 254866 346448 254898
rect 376848 255454 377168 255486
rect 376848 255218 376890 255454
rect 377126 255218 377168 255454
rect 376848 255134 377168 255218
rect 376848 254898 376890 255134
rect 377126 254898 377168 255134
rect 376848 254866 377168 254898
rect 407568 255454 407888 255486
rect 407568 255218 407610 255454
rect 407846 255218 407888 255454
rect 407568 255134 407888 255218
rect 407568 254898 407610 255134
rect 407846 254898 407888 255134
rect 407568 254866 407888 254898
rect 438288 255454 438608 255486
rect 438288 255218 438330 255454
rect 438566 255218 438608 255454
rect 438288 255134 438608 255218
rect 438288 254898 438330 255134
rect 438566 254898 438608 255134
rect 438288 254866 438608 254898
rect 469008 255454 469328 255486
rect 469008 255218 469050 255454
rect 469286 255218 469328 255454
rect 469008 255134 469328 255218
rect 469008 254898 469050 255134
rect 469286 254898 469328 255134
rect 469008 254866 469328 254898
rect 499728 255454 500048 255486
rect 499728 255218 499770 255454
rect 500006 255218 500048 255454
rect 499728 255134 500048 255218
rect 499728 254898 499770 255134
rect 500006 254898 500048 255134
rect 499728 254866 500048 254898
rect 530448 255454 530768 255486
rect 530448 255218 530490 255454
rect 530726 255218 530768 255454
rect 530448 255134 530768 255218
rect 530448 254898 530490 255134
rect 530726 254898 530768 255134
rect 530448 254866 530768 254898
rect 561168 255454 561488 255486
rect 561168 255218 561210 255454
rect 561446 255218 561488 255454
rect 561168 255134 561488 255218
rect 561168 254898 561210 255134
rect 561446 254898 561488 255134
rect 561168 254866 561488 254898
rect 567234 244894 567854 280338
rect 567234 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 567854 244894
rect 567234 244574 567854 244658
rect 567234 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 567854 244574
rect 23568 237454 23888 237486
rect 23568 237218 23610 237454
rect 23846 237218 23888 237454
rect 23568 237134 23888 237218
rect 23568 236898 23610 237134
rect 23846 236898 23888 237134
rect 23568 236866 23888 236898
rect 54288 237454 54608 237486
rect 54288 237218 54330 237454
rect 54566 237218 54608 237454
rect 54288 237134 54608 237218
rect 54288 236898 54330 237134
rect 54566 236898 54608 237134
rect 54288 236866 54608 236898
rect 85008 237454 85328 237486
rect 85008 237218 85050 237454
rect 85286 237218 85328 237454
rect 85008 237134 85328 237218
rect 85008 236898 85050 237134
rect 85286 236898 85328 237134
rect 85008 236866 85328 236898
rect 115728 237454 116048 237486
rect 115728 237218 115770 237454
rect 116006 237218 116048 237454
rect 115728 237134 116048 237218
rect 115728 236898 115770 237134
rect 116006 236898 116048 237134
rect 115728 236866 116048 236898
rect 146448 237454 146768 237486
rect 146448 237218 146490 237454
rect 146726 237218 146768 237454
rect 146448 237134 146768 237218
rect 146448 236898 146490 237134
rect 146726 236898 146768 237134
rect 146448 236866 146768 236898
rect 177168 237454 177488 237486
rect 177168 237218 177210 237454
rect 177446 237218 177488 237454
rect 177168 237134 177488 237218
rect 177168 236898 177210 237134
rect 177446 236898 177488 237134
rect 177168 236866 177488 236898
rect 207888 237454 208208 237486
rect 207888 237218 207930 237454
rect 208166 237218 208208 237454
rect 207888 237134 208208 237218
rect 207888 236898 207930 237134
rect 208166 236898 208208 237134
rect 207888 236866 208208 236898
rect 238608 237454 238928 237486
rect 238608 237218 238650 237454
rect 238886 237218 238928 237454
rect 238608 237134 238928 237218
rect 238608 236898 238650 237134
rect 238886 236898 238928 237134
rect 238608 236866 238928 236898
rect 269328 237454 269648 237486
rect 269328 237218 269370 237454
rect 269606 237218 269648 237454
rect 269328 237134 269648 237218
rect 269328 236898 269370 237134
rect 269606 236898 269648 237134
rect 269328 236866 269648 236898
rect 300048 237454 300368 237486
rect 300048 237218 300090 237454
rect 300326 237218 300368 237454
rect 300048 237134 300368 237218
rect 300048 236898 300090 237134
rect 300326 236898 300368 237134
rect 300048 236866 300368 236898
rect 330768 237454 331088 237486
rect 330768 237218 330810 237454
rect 331046 237218 331088 237454
rect 330768 237134 331088 237218
rect 330768 236898 330810 237134
rect 331046 236898 331088 237134
rect 330768 236866 331088 236898
rect 361488 237454 361808 237486
rect 361488 237218 361530 237454
rect 361766 237218 361808 237454
rect 361488 237134 361808 237218
rect 361488 236898 361530 237134
rect 361766 236898 361808 237134
rect 361488 236866 361808 236898
rect 392208 237454 392528 237486
rect 392208 237218 392250 237454
rect 392486 237218 392528 237454
rect 392208 237134 392528 237218
rect 392208 236898 392250 237134
rect 392486 236898 392528 237134
rect 392208 236866 392528 236898
rect 422928 237454 423248 237486
rect 422928 237218 422970 237454
rect 423206 237218 423248 237454
rect 422928 237134 423248 237218
rect 422928 236898 422970 237134
rect 423206 236898 423248 237134
rect 422928 236866 423248 236898
rect 453648 237454 453968 237486
rect 453648 237218 453690 237454
rect 453926 237218 453968 237454
rect 453648 237134 453968 237218
rect 453648 236898 453690 237134
rect 453926 236898 453968 237134
rect 453648 236866 453968 236898
rect 484368 237454 484688 237486
rect 484368 237218 484410 237454
rect 484646 237218 484688 237454
rect 484368 237134 484688 237218
rect 484368 236898 484410 237134
rect 484646 236898 484688 237134
rect 484368 236866 484688 236898
rect 515088 237454 515408 237486
rect 515088 237218 515130 237454
rect 515366 237218 515408 237454
rect 515088 237134 515408 237218
rect 515088 236898 515130 237134
rect 515366 236898 515408 237134
rect 515088 236866 515408 236898
rect 545808 237454 546128 237486
rect 545808 237218 545850 237454
rect 546086 237218 546128 237454
rect 545808 237134 546128 237218
rect 545808 236898 545850 237134
rect 546086 236898 546128 237134
rect 545808 236866 546128 236898
rect -2006 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 -1386 219454
rect -2006 219134 -1386 219218
rect -2006 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 -1386 219134
rect -2006 183454 -1386 218898
rect 8208 219454 8528 219486
rect 8208 219218 8250 219454
rect 8486 219218 8528 219454
rect 8208 219134 8528 219218
rect 8208 218898 8250 219134
rect 8486 218898 8528 219134
rect 8208 218866 8528 218898
rect 38928 219454 39248 219486
rect 38928 219218 38970 219454
rect 39206 219218 39248 219454
rect 38928 219134 39248 219218
rect 38928 218898 38970 219134
rect 39206 218898 39248 219134
rect 38928 218866 39248 218898
rect 69648 219454 69968 219486
rect 69648 219218 69690 219454
rect 69926 219218 69968 219454
rect 69648 219134 69968 219218
rect 69648 218898 69690 219134
rect 69926 218898 69968 219134
rect 69648 218866 69968 218898
rect 100368 219454 100688 219486
rect 100368 219218 100410 219454
rect 100646 219218 100688 219454
rect 100368 219134 100688 219218
rect 100368 218898 100410 219134
rect 100646 218898 100688 219134
rect 100368 218866 100688 218898
rect 131088 219454 131408 219486
rect 131088 219218 131130 219454
rect 131366 219218 131408 219454
rect 131088 219134 131408 219218
rect 131088 218898 131130 219134
rect 131366 218898 131408 219134
rect 131088 218866 131408 218898
rect 161808 219454 162128 219486
rect 161808 219218 161850 219454
rect 162086 219218 162128 219454
rect 161808 219134 162128 219218
rect 161808 218898 161850 219134
rect 162086 218898 162128 219134
rect 161808 218866 162128 218898
rect 192528 219454 192848 219486
rect 192528 219218 192570 219454
rect 192806 219218 192848 219454
rect 192528 219134 192848 219218
rect 192528 218898 192570 219134
rect 192806 218898 192848 219134
rect 192528 218866 192848 218898
rect 223248 219454 223568 219486
rect 223248 219218 223290 219454
rect 223526 219218 223568 219454
rect 223248 219134 223568 219218
rect 223248 218898 223290 219134
rect 223526 218898 223568 219134
rect 223248 218866 223568 218898
rect 253968 219454 254288 219486
rect 253968 219218 254010 219454
rect 254246 219218 254288 219454
rect 253968 219134 254288 219218
rect 253968 218898 254010 219134
rect 254246 218898 254288 219134
rect 253968 218866 254288 218898
rect 284688 219454 285008 219486
rect 284688 219218 284730 219454
rect 284966 219218 285008 219454
rect 284688 219134 285008 219218
rect 284688 218898 284730 219134
rect 284966 218898 285008 219134
rect 284688 218866 285008 218898
rect 315408 219454 315728 219486
rect 315408 219218 315450 219454
rect 315686 219218 315728 219454
rect 315408 219134 315728 219218
rect 315408 218898 315450 219134
rect 315686 218898 315728 219134
rect 315408 218866 315728 218898
rect 346128 219454 346448 219486
rect 346128 219218 346170 219454
rect 346406 219218 346448 219454
rect 346128 219134 346448 219218
rect 346128 218898 346170 219134
rect 346406 218898 346448 219134
rect 346128 218866 346448 218898
rect 376848 219454 377168 219486
rect 376848 219218 376890 219454
rect 377126 219218 377168 219454
rect 376848 219134 377168 219218
rect 376848 218898 376890 219134
rect 377126 218898 377168 219134
rect 376848 218866 377168 218898
rect 407568 219454 407888 219486
rect 407568 219218 407610 219454
rect 407846 219218 407888 219454
rect 407568 219134 407888 219218
rect 407568 218898 407610 219134
rect 407846 218898 407888 219134
rect 407568 218866 407888 218898
rect 438288 219454 438608 219486
rect 438288 219218 438330 219454
rect 438566 219218 438608 219454
rect 438288 219134 438608 219218
rect 438288 218898 438330 219134
rect 438566 218898 438608 219134
rect 438288 218866 438608 218898
rect 469008 219454 469328 219486
rect 469008 219218 469050 219454
rect 469286 219218 469328 219454
rect 469008 219134 469328 219218
rect 469008 218898 469050 219134
rect 469286 218898 469328 219134
rect 469008 218866 469328 218898
rect 499728 219454 500048 219486
rect 499728 219218 499770 219454
rect 500006 219218 500048 219454
rect 499728 219134 500048 219218
rect 499728 218898 499770 219134
rect 500006 218898 500048 219134
rect 499728 218866 500048 218898
rect 530448 219454 530768 219486
rect 530448 219218 530490 219454
rect 530726 219218 530768 219454
rect 530448 219134 530768 219218
rect 530448 218898 530490 219134
rect 530726 218898 530768 219134
rect 530448 218866 530768 218898
rect 561168 219454 561488 219486
rect 561168 219218 561210 219454
rect 561446 219218 561488 219454
rect 561168 219134 561488 219218
rect 561168 218898 561210 219134
rect 561446 218898 561488 219134
rect 561168 218866 561488 218898
rect 567234 208894 567854 244338
rect 567234 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 567854 208894
rect 567234 208574 567854 208658
rect 567234 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 567854 208574
rect 23568 201454 23888 201486
rect 23568 201218 23610 201454
rect 23846 201218 23888 201454
rect 23568 201134 23888 201218
rect 23568 200898 23610 201134
rect 23846 200898 23888 201134
rect 23568 200866 23888 200898
rect 54288 201454 54608 201486
rect 54288 201218 54330 201454
rect 54566 201218 54608 201454
rect 54288 201134 54608 201218
rect 54288 200898 54330 201134
rect 54566 200898 54608 201134
rect 54288 200866 54608 200898
rect 85008 201454 85328 201486
rect 85008 201218 85050 201454
rect 85286 201218 85328 201454
rect 85008 201134 85328 201218
rect 85008 200898 85050 201134
rect 85286 200898 85328 201134
rect 85008 200866 85328 200898
rect 115728 201454 116048 201486
rect 115728 201218 115770 201454
rect 116006 201218 116048 201454
rect 115728 201134 116048 201218
rect 115728 200898 115770 201134
rect 116006 200898 116048 201134
rect 115728 200866 116048 200898
rect 146448 201454 146768 201486
rect 146448 201218 146490 201454
rect 146726 201218 146768 201454
rect 146448 201134 146768 201218
rect 146448 200898 146490 201134
rect 146726 200898 146768 201134
rect 146448 200866 146768 200898
rect 177168 201454 177488 201486
rect 177168 201218 177210 201454
rect 177446 201218 177488 201454
rect 177168 201134 177488 201218
rect 177168 200898 177210 201134
rect 177446 200898 177488 201134
rect 177168 200866 177488 200898
rect 207888 201454 208208 201486
rect 207888 201218 207930 201454
rect 208166 201218 208208 201454
rect 207888 201134 208208 201218
rect 207888 200898 207930 201134
rect 208166 200898 208208 201134
rect 207888 200866 208208 200898
rect 238608 201454 238928 201486
rect 238608 201218 238650 201454
rect 238886 201218 238928 201454
rect 238608 201134 238928 201218
rect 238608 200898 238650 201134
rect 238886 200898 238928 201134
rect 238608 200866 238928 200898
rect 269328 201454 269648 201486
rect 269328 201218 269370 201454
rect 269606 201218 269648 201454
rect 269328 201134 269648 201218
rect 269328 200898 269370 201134
rect 269606 200898 269648 201134
rect 269328 200866 269648 200898
rect 300048 201454 300368 201486
rect 300048 201218 300090 201454
rect 300326 201218 300368 201454
rect 300048 201134 300368 201218
rect 300048 200898 300090 201134
rect 300326 200898 300368 201134
rect 300048 200866 300368 200898
rect 330768 201454 331088 201486
rect 330768 201218 330810 201454
rect 331046 201218 331088 201454
rect 330768 201134 331088 201218
rect 330768 200898 330810 201134
rect 331046 200898 331088 201134
rect 330768 200866 331088 200898
rect 361488 201454 361808 201486
rect 361488 201218 361530 201454
rect 361766 201218 361808 201454
rect 361488 201134 361808 201218
rect 361488 200898 361530 201134
rect 361766 200898 361808 201134
rect 361488 200866 361808 200898
rect 392208 201454 392528 201486
rect 392208 201218 392250 201454
rect 392486 201218 392528 201454
rect 392208 201134 392528 201218
rect 392208 200898 392250 201134
rect 392486 200898 392528 201134
rect 392208 200866 392528 200898
rect 422928 201454 423248 201486
rect 422928 201218 422970 201454
rect 423206 201218 423248 201454
rect 422928 201134 423248 201218
rect 422928 200898 422970 201134
rect 423206 200898 423248 201134
rect 422928 200866 423248 200898
rect 453648 201454 453968 201486
rect 453648 201218 453690 201454
rect 453926 201218 453968 201454
rect 453648 201134 453968 201218
rect 453648 200898 453690 201134
rect 453926 200898 453968 201134
rect 453648 200866 453968 200898
rect 484368 201454 484688 201486
rect 484368 201218 484410 201454
rect 484646 201218 484688 201454
rect 484368 201134 484688 201218
rect 484368 200898 484410 201134
rect 484646 200898 484688 201134
rect 484368 200866 484688 200898
rect 515088 201454 515408 201486
rect 515088 201218 515130 201454
rect 515366 201218 515408 201454
rect 515088 201134 515408 201218
rect 515088 200898 515130 201134
rect 515366 200898 515408 201134
rect 515088 200866 515408 200898
rect 545808 201454 546128 201486
rect 545808 201218 545850 201454
rect 546086 201218 546128 201454
rect 545808 201134 546128 201218
rect 545808 200898 545850 201134
rect 546086 200898 546128 201134
rect 545808 200866 546128 200898
rect -2006 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 -1386 183454
rect -2006 183134 -1386 183218
rect -2006 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 -1386 183134
rect -2006 147454 -1386 182898
rect 8208 183454 8528 183486
rect 8208 183218 8250 183454
rect 8486 183218 8528 183454
rect 8208 183134 8528 183218
rect 8208 182898 8250 183134
rect 8486 182898 8528 183134
rect 8208 182866 8528 182898
rect 38928 183454 39248 183486
rect 38928 183218 38970 183454
rect 39206 183218 39248 183454
rect 38928 183134 39248 183218
rect 38928 182898 38970 183134
rect 39206 182898 39248 183134
rect 38928 182866 39248 182898
rect 69648 183454 69968 183486
rect 69648 183218 69690 183454
rect 69926 183218 69968 183454
rect 69648 183134 69968 183218
rect 69648 182898 69690 183134
rect 69926 182898 69968 183134
rect 69648 182866 69968 182898
rect 100368 183454 100688 183486
rect 100368 183218 100410 183454
rect 100646 183218 100688 183454
rect 100368 183134 100688 183218
rect 100368 182898 100410 183134
rect 100646 182898 100688 183134
rect 100368 182866 100688 182898
rect 131088 183454 131408 183486
rect 131088 183218 131130 183454
rect 131366 183218 131408 183454
rect 131088 183134 131408 183218
rect 131088 182898 131130 183134
rect 131366 182898 131408 183134
rect 131088 182866 131408 182898
rect 161808 183454 162128 183486
rect 161808 183218 161850 183454
rect 162086 183218 162128 183454
rect 161808 183134 162128 183218
rect 161808 182898 161850 183134
rect 162086 182898 162128 183134
rect 161808 182866 162128 182898
rect 192528 183454 192848 183486
rect 192528 183218 192570 183454
rect 192806 183218 192848 183454
rect 192528 183134 192848 183218
rect 192528 182898 192570 183134
rect 192806 182898 192848 183134
rect 192528 182866 192848 182898
rect 223248 183454 223568 183486
rect 223248 183218 223290 183454
rect 223526 183218 223568 183454
rect 223248 183134 223568 183218
rect 223248 182898 223290 183134
rect 223526 182898 223568 183134
rect 223248 182866 223568 182898
rect 253968 183454 254288 183486
rect 253968 183218 254010 183454
rect 254246 183218 254288 183454
rect 253968 183134 254288 183218
rect 253968 182898 254010 183134
rect 254246 182898 254288 183134
rect 253968 182866 254288 182898
rect 284688 183454 285008 183486
rect 284688 183218 284730 183454
rect 284966 183218 285008 183454
rect 284688 183134 285008 183218
rect 284688 182898 284730 183134
rect 284966 182898 285008 183134
rect 284688 182866 285008 182898
rect 315408 183454 315728 183486
rect 315408 183218 315450 183454
rect 315686 183218 315728 183454
rect 315408 183134 315728 183218
rect 315408 182898 315450 183134
rect 315686 182898 315728 183134
rect 315408 182866 315728 182898
rect 346128 183454 346448 183486
rect 346128 183218 346170 183454
rect 346406 183218 346448 183454
rect 346128 183134 346448 183218
rect 346128 182898 346170 183134
rect 346406 182898 346448 183134
rect 346128 182866 346448 182898
rect 376848 183454 377168 183486
rect 376848 183218 376890 183454
rect 377126 183218 377168 183454
rect 376848 183134 377168 183218
rect 376848 182898 376890 183134
rect 377126 182898 377168 183134
rect 376848 182866 377168 182898
rect 407568 183454 407888 183486
rect 407568 183218 407610 183454
rect 407846 183218 407888 183454
rect 407568 183134 407888 183218
rect 407568 182898 407610 183134
rect 407846 182898 407888 183134
rect 407568 182866 407888 182898
rect 438288 183454 438608 183486
rect 438288 183218 438330 183454
rect 438566 183218 438608 183454
rect 438288 183134 438608 183218
rect 438288 182898 438330 183134
rect 438566 182898 438608 183134
rect 438288 182866 438608 182898
rect 469008 183454 469328 183486
rect 469008 183218 469050 183454
rect 469286 183218 469328 183454
rect 469008 183134 469328 183218
rect 469008 182898 469050 183134
rect 469286 182898 469328 183134
rect 469008 182866 469328 182898
rect 499728 183454 500048 183486
rect 499728 183218 499770 183454
rect 500006 183218 500048 183454
rect 499728 183134 500048 183218
rect 499728 182898 499770 183134
rect 500006 182898 500048 183134
rect 499728 182866 500048 182898
rect 530448 183454 530768 183486
rect 530448 183218 530490 183454
rect 530726 183218 530768 183454
rect 530448 183134 530768 183218
rect 530448 182898 530490 183134
rect 530726 182898 530768 183134
rect 530448 182866 530768 182898
rect 561168 183454 561488 183486
rect 561168 183218 561210 183454
rect 561446 183218 561488 183454
rect 561168 183134 561488 183218
rect 561168 182898 561210 183134
rect 561446 182898 561488 183134
rect 561168 182866 561488 182898
rect 567234 172894 567854 208338
rect 567234 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 567854 172894
rect 567234 172574 567854 172658
rect 567234 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 567854 172574
rect 23568 165454 23888 165486
rect 23568 165218 23610 165454
rect 23846 165218 23888 165454
rect 23568 165134 23888 165218
rect 23568 164898 23610 165134
rect 23846 164898 23888 165134
rect 23568 164866 23888 164898
rect 54288 165454 54608 165486
rect 54288 165218 54330 165454
rect 54566 165218 54608 165454
rect 54288 165134 54608 165218
rect 54288 164898 54330 165134
rect 54566 164898 54608 165134
rect 54288 164866 54608 164898
rect 85008 165454 85328 165486
rect 85008 165218 85050 165454
rect 85286 165218 85328 165454
rect 85008 165134 85328 165218
rect 85008 164898 85050 165134
rect 85286 164898 85328 165134
rect 85008 164866 85328 164898
rect 115728 165454 116048 165486
rect 115728 165218 115770 165454
rect 116006 165218 116048 165454
rect 115728 165134 116048 165218
rect 115728 164898 115770 165134
rect 116006 164898 116048 165134
rect 115728 164866 116048 164898
rect 146448 165454 146768 165486
rect 146448 165218 146490 165454
rect 146726 165218 146768 165454
rect 146448 165134 146768 165218
rect 146448 164898 146490 165134
rect 146726 164898 146768 165134
rect 146448 164866 146768 164898
rect 177168 165454 177488 165486
rect 177168 165218 177210 165454
rect 177446 165218 177488 165454
rect 177168 165134 177488 165218
rect 177168 164898 177210 165134
rect 177446 164898 177488 165134
rect 177168 164866 177488 164898
rect 207888 165454 208208 165486
rect 207888 165218 207930 165454
rect 208166 165218 208208 165454
rect 207888 165134 208208 165218
rect 207888 164898 207930 165134
rect 208166 164898 208208 165134
rect 207888 164866 208208 164898
rect 238608 165454 238928 165486
rect 238608 165218 238650 165454
rect 238886 165218 238928 165454
rect 238608 165134 238928 165218
rect 238608 164898 238650 165134
rect 238886 164898 238928 165134
rect 238608 164866 238928 164898
rect 269328 165454 269648 165486
rect 269328 165218 269370 165454
rect 269606 165218 269648 165454
rect 269328 165134 269648 165218
rect 269328 164898 269370 165134
rect 269606 164898 269648 165134
rect 269328 164866 269648 164898
rect 300048 165454 300368 165486
rect 300048 165218 300090 165454
rect 300326 165218 300368 165454
rect 300048 165134 300368 165218
rect 300048 164898 300090 165134
rect 300326 164898 300368 165134
rect 300048 164866 300368 164898
rect 330768 165454 331088 165486
rect 330768 165218 330810 165454
rect 331046 165218 331088 165454
rect 330768 165134 331088 165218
rect 330768 164898 330810 165134
rect 331046 164898 331088 165134
rect 330768 164866 331088 164898
rect 361488 165454 361808 165486
rect 361488 165218 361530 165454
rect 361766 165218 361808 165454
rect 361488 165134 361808 165218
rect 361488 164898 361530 165134
rect 361766 164898 361808 165134
rect 361488 164866 361808 164898
rect 392208 165454 392528 165486
rect 392208 165218 392250 165454
rect 392486 165218 392528 165454
rect 392208 165134 392528 165218
rect 392208 164898 392250 165134
rect 392486 164898 392528 165134
rect 392208 164866 392528 164898
rect 422928 165454 423248 165486
rect 422928 165218 422970 165454
rect 423206 165218 423248 165454
rect 422928 165134 423248 165218
rect 422928 164898 422970 165134
rect 423206 164898 423248 165134
rect 422928 164866 423248 164898
rect 453648 165454 453968 165486
rect 453648 165218 453690 165454
rect 453926 165218 453968 165454
rect 453648 165134 453968 165218
rect 453648 164898 453690 165134
rect 453926 164898 453968 165134
rect 453648 164866 453968 164898
rect 484368 165454 484688 165486
rect 484368 165218 484410 165454
rect 484646 165218 484688 165454
rect 484368 165134 484688 165218
rect 484368 164898 484410 165134
rect 484646 164898 484688 165134
rect 484368 164866 484688 164898
rect 515088 165454 515408 165486
rect 515088 165218 515130 165454
rect 515366 165218 515408 165454
rect 515088 165134 515408 165218
rect 515088 164898 515130 165134
rect 515366 164898 515408 165134
rect 515088 164866 515408 164898
rect 545808 165454 546128 165486
rect 545808 165218 545850 165454
rect 546086 165218 546128 165454
rect 545808 165134 546128 165218
rect 545808 164898 545850 165134
rect 546086 164898 546128 165134
rect 545808 164866 546128 164898
rect -2006 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 -1386 147454
rect -2006 147134 -1386 147218
rect -2006 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 -1386 147134
rect -2006 111454 -1386 146898
rect 8208 147454 8528 147486
rect 8208 147218 8250 147454
rect 8486 147218 8528 147454
rect 8208 147134 8528 147218
rect 8208 146898 8250 147134
rect 8486 146898 8528 147134
rect 8208 146866 8528 146898
rect 38928 147454 39248 147486
rect 38928 147218 38970 147454
rect 39206 147218 39248 147454
rect 38928 147134 39248 147218
rect 38928 146898 38970 147134
rect 39206 146898 39248 147134
rect 38928 146866 39248 146898
rect 69648 147454 69968 147486
rect 69648 147218 69690 147454
rect 69926 147218 69968 147454
rect 69648 147134 69968 147218
rect 69648 146898 69690 147134
rect 69926 146898 69968 147134
rect 69648 146866 69968 146898
rect 100368 147454 100688 147486
rect 100368 147218 100410 147454
rect 100646 147218 100688 147454
rect 100368 147134 100688 147218
rect 100368 146898 100410 147134
rect 100646 146898 100688 147134
rect 100368 146866 100688 146898
rect 131088 147454 131408 147486
rect 131088 147218 131130 147454
rect 131366 147218 131408 147454
rect 131088 147134 131408 147218
rect 131088 146898 131130 147134
rect 131366 146898 131408 147134
rect 131088 146866 131408 146898
rect 161808 147454 162128 147486
rect 161808 147218 161850 147454
rect 162086 147218 162128 147454
rect 161808 147134 162128 147218
rect 161808 146898 161850 147134
rect 162086 146898 162128 147134
rect 161808 146866 162128 146898
rect 192528 147454 192848 147486
rect 192528 147218 192570 147454
rect 192806 147218 192848 147454
rect 192528 147134 192848 147218
rect 192528 146898 192570 147134
rect 192806 146898 192848 147134
rect 192528 146866 192848 146898
rect 223248 147454 223568 147486
rect 223248 147218 223290 147454
rect 223526 147218 223568 147454
rect 223248 147134 223568 147218
rect 223248 146898 223290 147134
rect 223526 146898 223568 147134
rect 223248 146866 223568 146898
rect 253968 147454 254288 147486
rect 253968 147218 254010 147454
rect 254246 147218 254288 147454
rect 253968 147134 254288 147218
rect 253968 146898 254010 147134
rect 254246 146898 254288 147134
rect 253968 146866 254288 146898
rect 284688 147454 285008 147486
rect 284688 147218 284730 147454
rect 284966 147218 285008 147454
rect 284688 147134 285008 147218
rect 284688 146898 284730 147134
rect 284966 146898 285008 147134
rect 284688 146866 285008 146898
rect 315408 147454 315728 147486
rect 315408 147218 315450 147454
rect 315686 147218 315728 147454
rect 315408 147134 315728 147218
rect 315408 146898 315450 147134
rect 315686 146898 315728 147134
rect 315408 146866 315728 146898
rect 346128 147454 346448 147486
rect 346128 147218 346170 147454
rect 346406 147218 346448 147454
rect 346128 147134 346448 147218
rect 346128 146898 346170 147134
rect 346406 146898 346448 147134
rect 346128 146866 346448 146898
rect 376848 147454 377168 147486
rect 376848 147218 376890 147454
rect 377126 147218 377168 147454
rect 376848 147134 377168 147218
rect 376848 146898 376890 147134
rect 377126 146898 377168 147134
rect 376848 146866 377168 146898
rect 407568 147454 407888 147486
rect 407568 147218 407610 147454
rect 407846 147218 407888 147454
rect 407568 147134 407888 147218
rect 407568 146898 407610 147134
rect 407846 146898 407888 147134
rect 407568 146866 407888 146898
rect 438288 147454 438608 147486
rect 438288 147218 438330 147454
rect 438566 147218 438608 147454
rect 438288 147134 438608 147218
rect 438288 146898 438330 147134
rect 438566 146898 438608 147134
rect 438288 146866 438608 146898
rect 469008 147454 469328 147486
rect 469008 147218 469050 147454
rect 469286 147218 469328 147454
rect 469008 147134 469328 147218
rect 469008 146898 469050 147134
rect 469286 146898 469328 147134
rect 469008 146866 469328 146898
rect 499728 147454 500048 147486
rect 499728 147218 499770 147454
rect 500006 147218 500048 147454
rect 499728 147134 500048 147218
rect 499728 146898 499770 147134
rect 500006 146898 500048 147134
rect 499728 146866 500048 146898
rect 530448 147454 530768 147486
rect 530448 147218 530490 147454
rect 530726 147218 530768 147454
rect 530448 147134 530768 147218
rect 530448 146898 530490 147134
rect 530726 146898 530768 147134
rect 530448 146866 530768 146898
rect 561168 147454 561488 147486
rect 561168 147218 561210 147454
rect 561446 147218 561488 147454
rect 561168 147134 561488 147218
rect 561168 146898 561210 147134
rect 561446 146898 561488 147134
rect 561168 146866 561488 146898
rect 567234 136894 567854 172338
rect 567234 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 567854 136894
rect 567234 136574 567854 136658
rect 567234 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 567854 136574
rect 23568 129454 23888 129486
rect 23568 129218 23610 129454
rect 23846 129218 23888 129454
rect 23568 129134 23888 129218
rect 23568 128898 23610 129134
rect 23846 128898 23888 129134
rect 23568 128866 23888 128898
rect 54288 129454 54608 129486
rect 54288 129218 54330 129454
rect 54566 129218 54608 129454
rect 54288 129134 54608 129218
rect 54288 128898 54330 129134
rect 54566 128898 54608 129134
rect 54288 128866 54608 128898
rect 85008 129454 85328 129486
rect 85008 129218 85050 129454
rect 85286 129218 85328 129454
rect 85008 129134 85328 129218
rect 85008 128898 85050 129134
rect 85286 128898 85328 129134
rect 85008 128866 85328 128898
rect 115728 129454 116048 129486
rect 115728 129218 115770 129454
rect 116006 129218 116048 129454
rect 115728 129134 116048 129218
rect 115728 128898 115770 129134
rect 116006 128898 116048 129134
rect 115728 128866 116048 128898
rect 146448 129454 146768 129486
rect 146448 129218 146490 129454
rect 146726 129218 146768 129454
rect 146448 129134 146768 129218
rect 146448 128898 146490 129134
rect 146726 128898 146768 129134
rect 146448 128866 146768 128898
rect 177168 129454 177488 129486
rect 177168 129218 177210 129454
rect 177446 129218 177488 129454
rect 177168 129134 177488 129218
rect 177168 128898 177210 129134
rect 177446 128898 177488 129134
rect 177168 128866 177488 128898
rect 207888 129454 208208 129486
rect 207888 129218 207930 129454
rect 208166 129218 208208 129454
rect 207888 129134 208208 129218
rect 207888 128898 207930 129134
rect 208166 128898 208208 129134
rect 207888 128866 208208 128898
rect 238608 129454 238928 129486
rect 238608 129218 238650 129454
rect 238886 129218 238928 129454
rect 238608 129134 238928 129218
rect 238608 128898 238650 129134
rect 238886 128898 238928 129134
rect 238608 128866 238928 128898
rect 269328 129454 269648 129486
rect 269328 129218 269370 129454
rect 269606 129218 269648 129454
rect 269328 129134 269648 129218
rect 269328 128898 269370 129134
rect 269606 128898 269648 129134
rect 269328 128866 269648 128898
rect 300048 129454 300368 129486
rect 300048 129218 300090 129454
rect 300326 129218 300368 129454
rect 300048 129134 300368 129218
rect 300048 128898 300090 129134
rect 300326 128898 300368 129134
rect 300048 128866 300368 128898
rect 330768 129454 331088 129486
rect 330768 129218 330810 129454
rect 331046 129218 331088 129454
rect 330768 129134 331088 129218
rect 330768 128898 330810 129134
rect 331046 128898 331088 129134
rect 330768 128866 331088 128898
rect 361488 129454 361808 129486
rect 361488 129218 361530 129454
rect 361766 129218 361808 129454
rect 361488 129134 361808 129218
rect 361488 128898 361530 129134
rect 361766 128898 361808 129134
rect 361488 128866 361808 128898
rect 392208 129454 392528 129486
rect 392208 129218 392250 129454
rect 392486 129218 392528 129454
rect 392208 129134 392528 129218
rect 392208 128898 392250 129134
rect 392486 128898 392528 129134
rect 392208 128866 392528 128898
rect 422928 129454 423248 129486
rect 422928 129218 422970 129454
rect 423206 129218 423248 129454
rect 422928 129134 423248 129218
rect 422928 128898 422970 129134
rect 423206 128898 423248 129134
rect 422928 128866 423248 128898
rect 453648 129454 453968 129486
rect 453648 129218 453690 129454
rect 453926 129218 453968 129454
rect 453648 129134 453968 129218
rect 453648 128898 453690 129134
rect 453926 128898 453968 129134
rect 453648 128866 453968 128898
rect 484368 129454 484688 129486
rect 484368 129218 484410 129454
rect 484646 129218 484688 129454
rect 484368 129134 484688 129218
rect 484368 128898 484410 129134
rect 484646 128898 484688 129134
rect 484368 128866 484688 128898
rect 515088 129454 515408 129486
rect 515088 129218 515130 129454
rect 515366 129218 515408 129454
rect 515088 129134 515408 129218
rect 515088 128898 515130 129134
rect 515366 128898 515408 129134
rect 515088 128866 515408 128898
rect 545808 129454 546128 129486
rect 545808 129218 545850 129454
rect 546086 129218 546128 129454
rect 545808 129134 546128 129218
rect 545808 128898 545850 129134
rect 546086 128898 546128 129134
rect 545808 128866 546128 128898
rect -2006 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 -1386 111454
rect -2006 111134 -1386 111218
rect -2006 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 -1386 111134
rect -2006 75454 -1386 110898
rect 8208 111454 8528 111486
rect 8208 111218 8250 111454
rect 8486 111218 8528 111454
rect 8208 111134 8528 111218
rect 8208 110898 8250 111134
rect 8486 110898 8528 111134
rect 8208 110866 8528 110898
rect 38928 111454 39248 111486
rect 38928 111218 38970 111454
rect 39206 111218 39248 111454
rect 38928 111134 39248 111218
rect 38928 110898 38970 111134
rect 39206 110898 39248 111134
rect 38928 110866 39248 110898
rect 69648 111454 69968 111486
rect 69648 111218 69690 111454
rect 69926 111218 69968 111454
rect 69648 111134 69968 111218
rect 69648 110898 69690 111134
rect 69926 110898 69968 111134
rect 69648 110866 69968 110898
rect 100368 111454 100688 111486
rect 100368 111218 100410 111454
rect 100646 111218 100688 111454
rect 100368 111134 100688 111218
rect 100368 110898 100410 111134
rect 100646 110898 100688 111134
rect 100368 110866 100688 110898
rect 131088 111454 131408 111486
rect 131088 111218 131130 111454
rect 131366 111218 131408 111454
rect 131088 111134 131408 111218
rect 131088 110898 131130 111134
rect 131366 110898 131408 111134
rect 131088 110866 131408 110898
rect 161808 111454 162128 111486
rect 161808 111218 161850 111454
rect 162086 111218 162128 111454
rect 161808 111134 162128 111218
rect 161808 110898 161850 111134
rect 162086 110898 162128 111134
rect 161808 110866 162128 110898
rect 192528 111454 192848 111486
rect 192528 111218 192570 111454
rect 192806 111218 192848 111454
rect 192528 111134 192848 111218
rect 192528 110898 192570 111134
rect 192806 110898 192848 111134
rect 192528 110866 192848 110898
rect 223248 111454 223568 111486
rect 223248 111218 223290 111454
rect 223526 111218 223568 111454
rect 223248 111134 223568 111218
rect 223248 110898 223290 111134
rect 223526 110898 223568 111134
rect 223248 110866 223568 110898
rect 253968 111454 254288 111486
rect 253968 111218 254010 111454
rect 254246 111218 254288 111454
rect 253968 111134 254288 111218
rect 253968 110898 254010 111134
rect 254246 110898 254288 111134
rect 253968 110866 254288 110898
rect 284688 111454 285008 111486
rect 284688 111218 284730 111454
rect 284966 111218 285008 111454
rect 284688 111134 285008 111218
rect 284688 110898 284730 111134
rect 284966 110898 285008 111134
rect 284688 110866 285008 110898
rect 315408 111454 315728 111486
rect 315408 111218 315450 111454
rect 315686 111218 315728 111454
rect 315408 111134 315728 111218
rect 315408 110898 315450 111134
rect 315686 110898 315728 111134
rect 315408 110866 315728 110898
rect 346128 111454 346448 111486
rect 346128 111218 346170 111454
rect 346406 111218 346448 111454
rect 346128 111134 346448 111218
rect 346128 110898 346170 111134
rect 346406 110898 346448 111134
rect 346128 110866 346448 110898
rect 376848 111454 377168 111486
rect 376848 111218 376890 111454
rect 377126 111218 377168 111454
rect 376848 111134 377168 111218
rect 376848 110898 376890 111134
rect 377126 110898 377168 111134
rect 376848 110866 377168 110898
rect 407568 111454 407888 111486
rect 407568 111218 407610 111454
rect 407846 111218 407888 111454
rect 407568 111134 407888 111218
rect 407568 110898 407610 111134
rect 407846 110898 407888 111134
rect 407568 110866 407888 110898
rect 438288 111454 438608 111486
rect 438288 111218 438330 111454
rect 438566 111218 438608 111454
rect 438288 111134 438608 111218
rect 438288 110898 438330 111134
rect 438566 110898 438608 111134
rect 438288 110866 438608 110898
rect 469008 111454 469328 111486
rect 469008 111218 469050 111454
rect 469286 111218 469328 111454
rect 469008 111134 469328 111218
rect 469008 110898 469050 111134
rect 469286 110898 469328 111134
rect 469008 110866 469328 110898
rect 499728 111454 500048 111486
rect 499728 111218 499770 111454
rect 500006 111218 500048 111454
rect 499728 111134 500048 111218
rect 499728 110898 499770 111134
rect 500006 110898 500048 111134
rect 499728 110866 500048 110898
rect 530448 111454 530768 111486
rect 530448 111218 530490 111454
rect 530726 111218 530768 111454
rect 530448 111134 530768 111218
rect 530448 110898 530490 111134
rect 530726 110898 530768 111134
rect 530448 110866 530768 110898
rect 561168 111454 561488 111486
rect 561168 111218 561210 111454
rect 561446 111218 561488 111454
rect 561168 111134 561488 111218
rect 561168 110898 561210 111134
rect 561446 110898 561488 111134
rect 561168 110866 561488 110898
rect 567234 100894 567854 136338
rect 567234 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 567854 100894
rect 567234 100574 567854 100658
rect 567234 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 567854 100574
rect 23568 93454 23888 93486
rect 23568 93218 23610 93454
rect 23846 93218 23888 93454
rect 23568 93134 23888 93218
rect 23568 92898 23610 93134
rect 23846 92898 23888 93134
rect 23568 92866 23888 92898
rect 54288 93454 54608 93486
rect 54288 93218 54330 93454
rect 54566 93218 54608 93454
rect 54288 93134 54608 93218
rect 54288 92898 54330 93134
rect 54566 92898 54608 93134
rect 54288 92866 54608 92898
rect 85008 93454 85328 93486
rect 85008 93218 85050 93454
rect 85286 93218 85328 93454
rect 85008 93134 85328 93218
rect 85008 92898 85050 93134
rect 85286 92898 85328 93134
rect 85008 92866 85328 92898
rect 115728 93454 116048 93486
rect 115728 93218 115770 93454
rect 116006 93218 116048 93454
rect 115728 93134 116048 93218
rect 115728 92898 115770 93134
rect 116006 92898 116048 93134
rect 115728 92866 116048 92898
rect 146448 93454 146768 93486
rect 146448 93218 146490 93454
rect 146726 93218 146768 93454
rect 146448 93134 146768 93218
rect 146448 92898 146490 93134
rect 146726 92898 146768 93134
rect 146448 92866 146768 92898
rect 177168 93454 177488 93486
rect 177168 93218 177210 93454
rect 177446 93218 177488 93454
rect 177168 93134 177488 93218
rect 177168 92898 177210 93134
rect 177446 92898 177488 93134
rect 177168 92866 177488 92898
rect 207888 93454 208208 93486
rect 207888 93218 207930 93454
rect 208166 93218 208208 93454
rect 207888 93134 208208 93218
rect 207888 92898 207930 93134
rect 208166 92898 208208 93134
rect 207888 92866 208208 92898
rect 238608 93454 238928 93486
rect 238608 93218 238650 93454
rect 238886 93218 238928 93454
rect 238608 93134 238928 93218
rect 238608 92898 238650 93134
rect 238886 92898 238928 93134
rect 238608 92866 238928 92898
rect 269328 93454 269648 93486
rect 269328 93218 269370 93454
rect 269606 93218 269648 93454
rect 269328 93134 269648 93218
rect 269328 92898 269370 93134
rect 269606 92898 269648 93134
rect 269328 92866 269648 92898
rect 300048 93454 300368 93486
rect 300048 93218 300090 93454
rect 300326 93218 300368 93454
rect 300048 93134 300368 93218
rect 300048 92898 300090 93134
rect 300326 92898 300368 93134
rect 300048 92866 300368 92898
rect 330768 93454 331088 93486
rect 330768 93218 330810 93454
rect 331046 93218 331088 93454
rect 330768 93134 331088 93218
rect 330768 92898 330810 93134
rect 331046 92898 331088 93134
rect 330768 92866 331088 92898
rect 361488 93454 361808 93486
rect 361488 93218 361530 93454
rect 361766 93218 361808 93454
rect 361488 93134 361808 93218
rect 361488 92898 361530 93134
rect 361766 92898 361808 93134
rect 361488 92866 361808 92898
rect 392208 93454 392528 93486
rect 392208 93218 392250 93454
rect 392486 93218 392528 93454
rect 392208 93134 392528 93218
rect 392208 92898 392250 93134
rect 392486 92898 392528 93134
rect 392208 92866 392528 92898
rect 422928 93454 423248 93486
rect 422928 93218 422970 93454
rect 423206 93218 423248 93454
rect 422928 93134 423248 93218
rect 422928 92898 422970 93134
rect 423206 92898 423248 93134
rect 422928 92866 423248 92898
rect 453648 93454 453968 93486
rect 453648 93218 453690 93454
rect 453926 93218 453968 93454
rect 453648 93134 453968 93218
rect 453648 92898 453690 93134
rect 453926 92898 453968 93134
rect 453648 92866 453968 92898
rect 484368 93454 484688 93486
rect 484368 93218 484410 93454
rect 484646 93218 484688 93454
rect 484368 93134 484688 93218
rect 484368 92898 484410 93134
rect 484646 92898 484688 93134
rect 484368 92866 484688 92898
rect 515088 93454 515408 93486
rect 515088 93218 515130 93454
rect 515366 93218 515408 93454
rect 515088 93134 515408 93218
rect 515088 92898 515130 93134
rect 515366 92898 515408 93134
rect 515088 92866 515408 92898
rect 545808 93454 546128 93486
rect 545808 93218 545850 93454
rect 546086 93218 546128 93454
rect 545808 93134 546128 93218
rect 545808 92898 545850 93134
rect 546086 92898 546128 93134
rect 545808 92866 546128 92898
rect -2006 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 -1386 75454
rect -2006 75134 -1386 75218
rect -2006 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 -1386 75134
rect -2006 39454 -1386 74898
rect 8208 75454 8528 75486
rect 8208 75218 8250 75454
rect 8486 75218 8528 75454
rect 8208 75134 8528 75218
rect 8208 74898 8250 75134
rect 8486 74898 8528 75134
rect 8208 74866 8528 74898
rect 38928 75454 39248 75486
rect 38928 75218 38970 75454
rect 39206 75218 39248 75454
rect 38928 75134 39248 75218
rect 38928 74898 38970 75134
rect 39206 74898 39248 75134
rect 38928 74866 39248 74898
rect 69648 75454 69968 75486
rect 69648 75218 69690 75454
rect 69926 75218 69968 75454
rect 69648 75134 69968 75218
rect 69648 74898 69690 75134
rect 69926 74898 69968 75134
rect 69648 74866 69968 74898
rect 100368 75454 100688 75486
rect 100368 75218 100410 75454
rect 100646 75218 100688 75454
rect 100368 75134 100688 75218
rect 100368 74898 100410 75134
rect 100646 74898 100688 75134
rect 100368 74866 100688 74898
rect 131088 75454 131408 75486
rect 131088 75218 131130 75454
rect 131366 75218 131408 75454
rect 131088 75134 131408 75218
rect 131088 74898 131130 75134
rect 131366 74898 131408 75134
rect 131088 74866 131408 74898
rect 161808 75454 162128 75486
rect 161808 75218 161850 75454
rect 162086 75218 162128 75454
rect 161808 75134 162128 75218
rect 161808 74898 161850 75134
rect 162086 74898 162128 75134
rect 161808 74866 162128 74898
rect 192528 75454 192848 75486
rect 192528 75218 192570 75454
rect 192806 75218 192848 75454
rect 192528 75134 192848 75218
rect 192528 74898 192570 75134
rect 192806 74898 192848 75134
rect 192528 74866 192848 74898
rect 223248 75454 223568 75486
rect 223248 75218 223290 75454
rect 223526 75218 223568 75454
rect 223248 75134 223568 75218
rect 223248 74898 223290 75134
rect 223526 74898 223568 75134
rect 223248 74866 223568 74898
rect 253968 75454 254288 75486
rect 253968 75218 254010 75454
rect 254246 75218 254288 75454
rect 253968 75134 254288 75218
rect 253968 74898 254010 75134
rect 254246 74898 254288 75134
rect 253968 74866 254288 74898
rect 284688 75454 285008 75486
rect 284688 75218 284730 75454
rect 284966 75218 285008 75454
rect 284688 75134 285008 75218
rect 284688 74898 284730 75134
rect 284966 74898 285008 75134
rect 284688 74866 285008 74898
rect 315408 75454 315728 75486
rect 315408 75218 315450 75454
rect 315686 75218 315728 75454
rect 315408 75134 315728 75218
rect 315408 74898 315450 75134
rect 315686 74898 315728 75134
rect 315408 74866 315728 74898
rect 346128 75454 346448 75486
rect 346128 75218 346170 75454
rect 346406 75218 346448 75454
rect 346128 75134 346448 75218
rect 346128 74898 346170 75134
rect 346406 74898 346448 75134
rect 346128 74866 346448 74898
rect 376848 75454 377168 75486
rect 376848 75218 376890 75454
rect 377126 75218 377168 75454
rect 376848 75134 377168 75218
rect 376848 74898 376890 75134
rect 377126 74898 377168 75134
rect 376848 74866 377168 74898
rect 407568 75454 407888 75486
rect 407568 75218 407610 75454
rect 407846 75218 407888 75454
rect 407568 75134 407888 75218
rect 407568 74898 407610 75134
rect 407846 74898 407888 75134
rect 407568 74866 407888 74898
rect 438288 75454 438608 75486
rect 438288 75218 438330 75454
rect 438566 75218 438608 75454
rect 438288 75134 438608 75218
rect 438288 74898 438330 75134
rect 438566 74898 438608 75134
rect 438288 74866 438608 74898
rect 469008 75454 469328 75486
rect 469008 75218 469050 75454
rect 469286 75218 469328 75454
rect 469008 75134 469328 75218
rect 469008 74898 469050 75134
rect 469286 74898 469328 75134
rect 469008 74866 469328 74898
rect 499728 75454 500048 75486
rect 499728 75218 499770 75454
rect 500006 75218 500048 75454
rect 499728 75134 500048 75218
rect 499728 74898 499770 75134
rect 500006 74898 500048 75134
rect 499728 74866 500048 74898
rect 530448 75454 530768 75486
rect 530448 75218 530490 75454
rect 530726 75218 530768 75454
rect 530448 75134 530768 75218
rect 530448 74898 530490 75134
rect 530726 74898 530768 75134
rect 530448 74866 530768 74898
rect 561168 75454 561488 75486
rect 561168 75218 561210 75454
rect 561446 75218 561488 75454
rect 561168 75134 561488 75218
rect 561168 74898 561210 75134
rect 561446 74898 561488 75134
rect 561168 74866 561488 74898
rect 567234 64894 567854 100338
rect 567234 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 567854 64894
rect 567234 64574 567854 64658
rect 567234 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 567854 64574
rect 23568 57454 23888 57486
rect 23568 57218 23610 57454
rect 23846 57218 23888 57454
rect 23568 57134 23888 57218
rect 23568 56898 23610 57134
rect 23846 56898 23888 57134
rect 23568 56866 23888 56898
rect 54288 57454 54608 57486
rect 54288 57218 54330 57454
rect 54566 57218 54608 57454
rect 54288 57134 54608 57218
rect 54288 56898 54330 57134
rect 54566 56898 54608 57134
rect 54288 56866 54608 56898
rect 85008 57454 85328 57486
rect 85008 57218 85050 57454
rect 85286 57218 85328 57454
rect 85008 57134 85328 57218
rect 85008 56898 85050 57134
rect 85286 56898 85328 57134
rect 85008 56866 85328 56898
rect 115728 57454 116048 57486
rect 115728 57218 115770 57454
rect 116006 57218 116048 57454
rect 115728 57134 116048 57218
rect 115728 56898 115770 57134
rect 116006 56898 116048 57134
rect 115728 56866 116048 56898
rect 146448 57454 146768 57486
rect 146448 57218 146490 57454
rect 146726 57218 146768 57454
rect 146448 57134 146768 57218
rect 146448 56898 146490 57134
rect 146726 56898 146768 57134
rect 146448 56866 146768 56898
rect 177168 57454 177488 57486
rect 177168 57218 177210 57454
rect 177446 57218 177488 57454
rect 177168 57134 177488 57218
rect 177168 56898 177210 57134
rect 177446 56898 177488 57134
rect 177168 56866 177488 56898
rect 207888 57454 208208 57486
rect 207888 57218 207930 57454
rect 208166 57218 208208 57454
rect 207888 57134 208208 57218
rect 207888 56898 207930 57134
rect 208166 56898 208208 57134
rect 207888 56866 208208 56898
rect 238608 57454 238928 57486
rect 238608 57218 238650 57454
rect 238886 57218 238928 57454
rect 238608 57134 238928 57218
rect 238608 56898 238650 57134
rect 238886 56898 238928 57134
rect 238608 56866 238928 56898
rect 269328 57454 269648 57486
rect 269328 57218 269370 57454
rect 269606 57218 269648 57454
rect 269328 57134 269648 57218
rect 269328 56898 269370 57134
rect 269606 56898 269648 57134
rect 269328 56866 269648 56898
rect 300048 57454 300368 57486
rect 300048 57218 300090 57454
rect 300326 57218 300368 57454
rect 300048 57134 300368 57218
rect 300048 56898 300090 57134
rect 300326 56898 300368 57134
rect 300048 56866 300368 56898
rect 330768 57454 331088 57486
rect 330768 57218 330810 57454
rect 331046 57218 331088 57454
rect 330768 57134 331088 57218
rect 330768 56898 330810 57134
rect 331046 56898 331088 57134
rect 330768 56866 331088 56898
rect 361488 57454 361808 57486
rect 361488 57218 361530 57454
rect 361766 57218 361808 57454
rect 361488 57134 361808 57218
rect 361488 56898 361530 57134
rect 361766 56898 361808 57134
rect 361488 56866 361808 56898
rect 392208 57454 392528 57486
rect 392208 57218 392250 57454
rect 392486 57218 392528 57454
rect 392208 57134 392528 57218
rect 392208 56898 392250 57134
rect 392486 56898 392528 57134
rect 392208 56866 392528 56898
rect 422928 57454 423248 57486
rect 422928 57218 422970 57454
rect 423206 57218 423248 57454
rect 422928 57134 423248 57218
rect 422928 56898 422970 57134
rect 423206 56898 423248 57134
rect 422928 56866 423248 56898
rect 453648 57454 453968 57486
rect 453648 57218 453690 57454
rect 453926 57218 453968 57454
rect 453648 57134 453968 57218
rect 453648 56898 453690 57134
rect 453926 56898 453968 57134
rect 453648 56866 453968 56898
rect 484368 57454 484688 57486
rect 484368 57218 484410 57454
rect 484646 57218 484688 57454
rect 484368 57134 484688 57218
rect 484368 56898 484410 57134
rect 484646 56898 484688 57134
rect 484368 56866 484688 56898
rect 515088 57454 515408 57486
rect 515088 57218 515130 57454
rect 515366 57218 515408 57454
rect 515088 57134 515408 57218
rect 515088 56898 515130 57134
rect 515366 56898 515408 57134
rect 515088 56866 515408 56898
rect 545808 57454 546128 57486
rect 545808 57218 545850 57454
rect 546086 57218 546128 57454
rect 545808 57134 546128 57218
rect 545808 56898 545850 57134
rect 546086 56898 546128 57134
rect 545808 56866 546128 56898
rect -2006 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 -1386 39454
rect -2006 39134 -1386 39218
rect -2006 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 -1386 39134
rect -2006 3454 -1386 38898
rect 8208 39454 8528 39486
rect 8208 39218 8250 39454
rect 8486 39218 8528 39454
rect 8208 39134 8528 39218
rect 8208 38898 8250 39134
rect 8486 38898 8528 39134
rect 8208 38866 8528 38898
rect 38928 39454 39248 39486
rect 38928 39218 38970 39454
rect 39206 39218 39248 39454
rect 38928 39134 39248 39218
rect 38928 38898 38970 39134
rect 39206 38898 39248 39134
rect 38928 38866 39248 38898
rect 69648 39454 69968 39486
rect 69648 39218 69690 39454
rect 69926 39218 69968 39454
rect 69648 39134 69968 39218
rect 69648 38898 69690 39134
rect 69926 38898 69968 39134
rect 69648 38866 69968 38898
rect 100368 39454 100688 39486
rect 100368 39218 100410 39454
rect 100646 39218 100688 39454
rect 100368 39134 100688 39218
rect 100368 38898 100410 39134
rect 100646 38898 100688 39134
rect 100368 38866 100688 38898
rect 131088 39454 131408 39486
rect 131088 39218 131130 39454
rect 131366 39218 131408 39454
rect 131088 39134 131408 39218
rect 131088 38898 131130 39134
rect 131366 38898 131408 39134
rect 131088 38866 131408 38898
rect 161808 39454 162128 39486
rect 161808 39218 161850 39454
rect 162086 39218 162128 39454
rect 161808 39134 162128 39218
rect 161808 38898 161850 39134
rect 162086 38898 162128 39134
rect 161808 38866 162128 38898
rect 192528 39454 192848 39486
rect 192528 39218 192570 39454
rect 192806 39218 192848 39454
rect 192528 39134 192848 39218
rect 192528 38898 192570 39134
rect 192806 38898 192848 39134
rect 192528 38866 192848 38898
rect 223248 39454 223568 39486
rect 223248 39218 223290 39454
rect 223526 39218 223568 39454
rect 223248 39134 223568 39218
rect 223248 38898 223290 39134
rect 223526 38898 223568 39134
rect 223248 38866 223568 38898
rect 253968 39454 254288 39486
rect 253968 39218 254010 39454
rect 254246 39218 254288 39454
rect 253968 39134 254288 39218
rect 253968 38898 254010 39134
rect 254246 38898 254288 39134
rect 253968 38866 254288 38898
rect 284688 39454 285008 39486
rect 284688 39218 284730 39454
rect 284966 39218 285008 39454
rect 284688 39134 285008 39218
rect 284688 38898 284730 39134
rect 284966 38898 285008 39134
rect 284688 38866 285008 38898
rect 315408 39454 315728 39486
rect 315408 39218 315450 39454
rect 315686 39218 315728 39454
rect 315408 39134 315728 39218
rect 315408 38898 315450 39134
rect 315686 38898 315728 39134
rect 315408 38866 315728 38898
rect 346128 39454 346448 39486
rect 346128 39218 346170 39454
rect 346406 39218 346448 39454
rect 346128 39134 346448 39218
rect 346128 38898 346170 39134
rect 346406 38898 346448 39134
rect 346128 38866 346448 38898
rect 376848 39454 377168 39486
rect 376848 39218 376890 39454
rect 377126 39218 377168 39454
rect 376848 39134 377168 39218
rect 376848 38898 376890 39134
rect 377126 38898 377168 39134
rect 376848 38866 377168 38898
rect 407568 39454 407888 39486
rect 407568 39218 407610 39454
rect 407846 39218 407888 39454
rect 407568 39134 407888 39218
rect 407568 38898 407610 39134
rect 407846 38898 407888 39134
rect 407568 38866 407888 38898
rect 438288 39454 438608 39486
rect 438288 39218 438330 39454
rect 438566 39218 438608 39454
rect 438288 39134 438608 39218
rect 438288 38898 438330 39134
rect 438566 38898 438608 39134
rect 438288 38866 438608 38898
rect 469008 39454 469328 39486
rect 469008 39218 469050 39454
rect 469286 39218 469328 39454
rect 469008 39134 469328 39218
rect 469008 38898 469050 39134
rect 469286 38898 469328 39134
rect 469008 38866 469328 38898
rect 499728 39454 500048 39486
rect 499728 39218 499770 39454
rect 500006 39218 500048 39454
rect 499728 39134 500048 39218
rect 499728 38898 499770 39134
rect 500006 38898 500048 39134
rect 499728 38866 500048 38898
rect 530448 39454 530768 39486
rect 530448 39218 530490 39454
rect 530726 39218 530768 39454
rect 530448 39134 530768 39218
rect 530448 38898 530490 39134
rect 530726 38898 530768 39134
rect 530448 38866 530768 38898
rect 561168 39454 561488 39486
rect 561168 39218 561210 39454
rect 561446 39218 561488 39454
rect 561168 39134 561488 39218
rect 561168 38898 561210 39134
rect 561446 38898 561488 39134
rect 561168 38866 561488 38898
rect 567234 28894 567854 64338
rect 567234 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 567854 28894
rect 567234 28574 567854 28658
rect 567234 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 567854 28574
rect 23568 21454 23888 21486
rect 23568 21218 23610 21454
rect 23846 21218 23888 21454
rect 23568 21134 23888 21218
rect 23568 20898 23610 21134
rect 23846 20898 23888 21134
rect 23568 20866 23888 20898
rect 54288 21454 54608 21486
rect 54288 21218 54330 21454
rect 54566 21218 54608 21454
rect 54288 21134 54608 21218
rect 54288 20898 54330 21134
rect 54566 20898 54608 21134
rect 54288 20866 54608 20898
rect 85008 21454 85328 21486
rect 85008 21218 85050 21454
rect 85286 21218 85328 21454
rect 85008 21134 85328 21218
rect 85008 20898 85050 21134
rect 85286 20898 85328 21134
rect 85008 20866 85328 20898
rect 115728 21454 116048 21486
rect 115728 21218 115770 21454
rect 116006 21218 116048 21454
rect 115728 21134 116048 21218
rect 115728 20898 115770 21134
rect 116006 20898 116048 21134
rect 115728 20866 116048 20898
rect 146448 21454 146768 21486
rect 146448 21218 146490 21454
rect 146726 21218 146768 21454
rect 146448 21134 146768 21218
rect 146448 20898 146490 21134
rect 146726 20898 146768 21134
rect 146448 20866 146768 20898
rect 177168 21454 177488 21486
rect 177168 21218 177210 21454
rect 177446 21218 177488 21454
rect 177168 21134 177488 21218
rect 177168 20898 177210 21134
rect 177446 20898 177488 21134
rect 177168 20866 177488 20898
rect 207888 21454 208208 21486
rect 207888 21218 207930 21454
rect 208166 21218 208208 21454
rect 207888 21134 208208 21218
rect 207888 20898 207930 21134
rect 208166 20898 208208 21134
rect 207888 20866 208208 20898
rect 238608 21454 238928 21486
rect 238608 21218 238650 21454
rect 238886 21218 238928 21454
rect 238608 21134 238928 21218
rect 238608 20898 238650 21134
rect 238886 20898 238928 21134
rect 238608 20866 238928 20898
rect 269328 21454 269648 21486
rect 269328 21218 269370 21454
rect 269606 21218 269648 21454
rect 269328 21134 269648 21218
rect 269328 20898 269370 21134
rect 269606 20898 269648 21134
rect 269328 20866 269648 20898
rect 300048 21454 300368 21486
rect 300048 21218 300090 21454
rect 300326 21218 300368 21454
rect 300048 21134 300368 21218
rect 300048 20898 300090 21134
rect 300326 20898 300368 21134
rect 300048 20866 300368 20898
rect 330768 21454 331088 21486
rect 330768 21218 330810 21454
rect 331046 21218 331088 21454
rect 330768 21134 331088 21218
rect 330768 20898 330810 21134
rect 331046 20898 331088 21134
rect 330768 20866 331088 20898
rect 361488 21454 361808 21486
rect 361488 21218 361530 21454
rect 361766 21218 361808 21454
rect 361488 21134 361808 21218
rect 361488 20898 361530 21134
rect 361766 20898 361808 21134
rect 361488 20866 361808 20898
rect 392208 21454 392528 21486
rect 392208 21218 392250 21454
rect 392486 21218 392528 21454
rect 392208 21134 392528 21218
rect 392208 20898 392250 21134
rect 392486 20898 392528 21134
rect 392208 20866 392528 20898
rect 422928 21454 423248 21486
rect 422928 21218 422970 21454
rect 423206 21218 423248 21454
rect 422928 21134 423248 21218
rect 422928 20898 422970 21134
rect 423206 20898 423248 21134
rect 422928 20866 423248 20898
rect 453648 21454 453968 21486
rect 453648 21218 453690 21454
rect 453926 21218 453968 21454
rect 453648 21134 453968 21218
rect 453648 20898 453690 21134
rect 453926 20898 453968 21134
rect 453648 20866 453968 20898
rect 484368 21454 484688 21486
rect 484368 21218 484410 21454
rect 484646 21218 484688 21454
rect 484368 21134 484688 21218
rect 484368 20898 484410 21134
rect 484646 20898 484688 21134
rect 484368 20866 484688 20898
rect 515088 21454 515408 21486
rect 515088 21218 515130 21454
rect 515366 21218 515408 21454
rect 515088 21134 515408 21218
rect 515088 20898 515130 21134
rect 515366 20898 515408 21134
rect 515088 20866 515408 20898
rect 545808 21454 546128 21486
rect 545808 21218 545850 21454
rect 546086 21218 546128 21454
rect 545808 21134 546128 21218
rect 545808 20898 545850 21134
rect 546086 20898 546128 21134
rect 545808 20866 546128 20898
rect -2006 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 -1386 3454
rect -2006 3134 -1386 3218
rect -2006 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 -1386 3134
rect -2006 -346 -1386 2898
rect 8208 3454 8528 3486
rect 8208 3218 8250 3454
rect 8486 3218 8528 3454
rect 8208 3134 8528 3218
rect 8208 2898 8250 3134
rect 8486 2898 8528 3134
rect 8208 2866 8528 2898
rect 38928 3454 39248 3486
rect 38928 3218 38970 3454
rect 39206 3218 39248 3454
rect 38928 3134 39248 3218
rect 38928 2898 38970 3134
rect 39206 2898 39248 3134
rect 38928 2866 39248 2898
rect 69648 3454 69968 3486
rect 69648 3218 69690 3454
rect 69926 3218 69968 3454
rect 69648 3134 69968 3218
rect 69648 2898 69690 3134
rect 69926 2898 69968 3134
rect 69648 2866 69968 2898
rect 100368 3454 100688 3486
rect 100368 3218 100410 3454
rect 100646 3218 100688 3454
rect 100368 3134 100688 3218
rect 100368 2898 100410 3134
rect 100646 2898 100688 3134
rect 100368 2866 100688 2898
rect 131088 3454 131408 3486
rect 131088 3218 131130 3454
rect 131366 3218 131408 3454
rect 131088 3134 131408 3218
rect 131088 2898 131130 3134
rect 131366 2898 131408 3134
rect 131088 2866 131408 2898
rect 161808 3454 162128 3486
rect 161808 3218 161850 3454
rect 162086 3218 162128 3454
rect 161808 3134 162128 3218
rect 161808 2898 161850 3134
rect 162086 2898 162128 3134
rect 161808 2866 162128 2898
rect 192528 3454 192848 3486
rect 192528 3218 192570 3454
rect 192806 3218 192848 3454
rect 192528 3134 192848 3218
rect 192528 2898 192570 3134
rect 192806 2898 192848 3134
rect 192528 2866 192848 2898
rect 223248 3454 223568 3486
rect 223248 3218 223290 3454
rect 223526 3218 223568 3454
rect 223248 3134 223568 3218
rect 223248 2898 223290 3134
rect 223526 2898 223568 3134
rect 223248 2866 223568 2898
rect 253968 3454 254288 3486
rect 253968 3218 254010 3454
rect 254246 3218 254288 3454
rect 253968 3134 254288 3218
rect 253968 2898 254010 3134
rect 254246 2898 254288 3134
rect 253968 2866 254288 2898
rect 284688 3454 285008 3486
rect 284688 3218 284730 3454
rect 284966 3218 285008 3454
rect 284688 3134 285008 3218
rect 284688 2898 284730 3134
rect 284966 2898 285008 3134
rect 284688 2866 285008 2898
rect 315408 3454 315728 3486
rect 315408 3218 315450 3454
rect 315686 3218 315728 3454
rect 315408 3134 315728 3218
rect 315408 2898 315450 3134
rect 315686 2898 315728 3134
rect 315408 2866 315728 2898
rect 346128 3454 346448 3486
rect 346128 3218 346170 3454
rect 346406 3218 346448 3454
rect 346128 3134 346448 3218
rect 346128 2898 346170 3134
rect 346406 2898 346448 3134
rect 346128 2866 346448 2898
rect 376848 3454 377168 3486
rect 376848 3218 376890 3454
rect 377126 3218 377168 3454
rect 376848 3134 377168 3218
rect 376848 2898 376890 3134
rect 377126 2898 377168 3134
rect 376848 2866 377168 2898
rect 407568 3454 407888 3486
rect 407568 3218 407610 3454
rect 407846 3218 407888 3454
rect 407568 3134 407888 3218
rect 407568 2898 407610 3134
rect 407846 2898 407888 3134
rect 407568 2866 407888 2898
rect 438288 3454 438608 3486
rect 438288 3218 438330 3454
rect 438566 3218 438608 3454
rect 438288 3134 438608 3218
rect 438288 2898 438330 3134
rect 438566 2898 438608 3134
rect 438288 2866 438608 2898
rect 469008 3454 469328 3486
rect 469008 3218 469050 3454
rect 469286 3218 469328 3454
rect 469008 3134 469328 3218
rect 469008 2898 469050 3134
rect 469286 2898 469328 3134
rect 469008 2866 469328 2898
rect 499728 3454 500048 3486
rect 499728 3218 499770 3454
rect 500006 3218 500048 3454
rect 499728 3134 500048 3218
rect 499728 2898 499770 3134
rect 500006 2898 500048 3134
rect 499728 2866 500048 2898
rect 530448 3454 530768 3486
rect 530448 3218 530490 3454
rect 530726 3218 530768 3454
rect 530448 3134 530768 3218
rect 530448 2898 530490 3134
rect 530726 2898 530768 3134
rect 530448 2866 530768 2898
rect 561168 3454 561488 3486
rect 561168 3218 561210 3454
rect 561446 3218 561488 3454
rect 561168 3134 561488 3218
rect 561168 2898 561210 3134
rect 561446 2898 561488 3134
rect 561168 2866 561488 2898
rect 531083 1460 531149 1461
rect 531083 1396 531084 1460
rect 531148 1396 531149 1460
rect 531083 1395 531149 1396
rect 205587 508 205653 509
rect 205587 444 205588 508
rect 205652 444 205653 508
rect 205587 443 205653 444
rect 205590 237 205650 443
rect 531086 237 531146 1395
rect 542859 1188 542925 1189
rect 542859 1124 542860 1188
rect 542924 1124 542925 1188
rect 542859 1123 542925 1124
rect 542491 916 542557 917
rect 542491 852 542492 916
rect 542556 852 542557 916
rect 542491 851 542557 852
rect 542494 509 542554 851
rect 542862 509 542922 1123
rect 551139 780 551205 781
rect 551139 716 551140 780
rect 551204 716 551205 780
rect 551139 715 551205 716
rect 542491 508 542557 509
rect 542491 444 542492 508
rect 542556 444 542557 508
rect 542491 443 542557 444
rect 542859 508 542925 509
rect 542859 444 542860 508
rect 542924 444 542925 508
rect 542859 443 542925 444
rect 551142 373 551202 715
rect 551139 372 551205 373
rect 551139 308 551140 372
rect 551204 308 551205 372
rect 551139 307 551205 308
rect 205587 236 205653 237
rect 205587 172 205588 236
rect 205652 172 205653 236
rect 205587 171 205653 172
rect 531083 236 531149 237
rect 531083 172 531084 236
rect 531148 172 531149 236
rect 531083 171 531149 172
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 -1386 -346
rect -2006 -666 -1386 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 -1386 -666
rect -2006 -934 -1386 -902
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 -2346 -1306
rect -2966 -1626 -2346 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 -2346 -1626
rect -2966 -1894 -2346 -1862
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 -3306 -2266
rect -3926 -2586 -3306 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 -3306 -2586
rect -3926 -2854 -3306 -2822
rect 5514 -2266 6134 -2000
rect 5514 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 6134 -2266
rect 5514 -2586 6134 -2502
rect 5514 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 6134 -2586
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 -4266 -3226
rect -4886 -3546 -4266 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 -4266 -3546
rect -4886 -3814 -4266 -3782
rect 5514 -3814 6134 -2822
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 -5226 -4186
rect -5846 -4506 -5226 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 -5226 -4506
rect -5846 -4774 -5226 -4742
rect 9234 -4186 9854 -2000
rect 9234 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 9854 -4186
rect 9234 -4506 9854 -4422
rect 9234 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 9854 -4506
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 -6186 -5146
rect -6806 -5466 -6186 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 -6186 -5466
rect -6806 -5734 -6186 -5702
rect 9234 -5734 9854 -4742
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 -7146 -6106
rect -7766 -6426 -7146 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 -7146 -6426
rect -7766 -6694 -7146 -6662
rect 12954 -6106 13574 -2000
rect 23514 -3226 24134 -2000
rect 23514 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 24134 -3226
rect 23514 -3546 24134 -3462
rect 23514 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 24134 -3546
rect 23514 -3814 24134 -3782
rect 27234 -5146 27854 -2000
rect 27234 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 27854 -5146
rect 27234 -5466 27854 -5382
rect 27234 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 27854 -5466
rect 27234 -5734 27854 -5702
rect 12954 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 13574 -6106
rect 12954 -6426 13574 -6342
rect 12954 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 13574 -6426
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 -8106 -7066
rect -8726 -7386 -8106 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 -8106 -7386
rect -8726 -7654 -8106 -7622
rect 12954 -7654 13574 -6662
rect 30954 -7066 31574 -2000
rect 41514 -2266 42134 -2000
rect 41514 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 42134 -2266
rect 41514 -2586 42134 -2502
rect 41514 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 42134 -2586
rect 41514 -3814 42134 -2822
rect 45234 -4186 45854 -2000
rect 45234 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 45854 -4186
rect 45234 -4506 45854 -4422
rect 45234 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 45854 -4506
rect 45234 -5734 45854 -4742
rect 30954 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 31574 -7066
rect 30954 -7386 31574 -7302
rect 30954 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 31574 -7386
rect 30954 -7654 31574 -7622
rect 48954 -6106 49574 -2000
rect 59514 -3226 60134 -2000
rect 59514 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 60134 -3226
rect 59514 -3546 60134 -3462
rect 59514 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 60134 -3546
rect 59514 -3814 60134 -3782
rect 63234 -5146 63854 -2000
rect 63234 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 63854 -5146
rect 63234 -5466 63854 -5382
rect 63234 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 63854 -5466
rect 63234 -5734 63854 -5702
rect 48954 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 49574 -6106
rect 48954 -6426 49574 -6342
rect 48954 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 49574 -6426
rect 48954 -7654 49574 -6662
rect 66954 -7066 67574 -2000
rect 77514 -2266 78134 -2000
rect 77514 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 78134 -2266
rect 77514 -2586 78134 -2502
rect 77514 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 78134 -2586
rect 77514 -3814 78134 -2822
rect 81234 -4186 81854 -2000
rect 81234 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 81854 -4186
rect 81234 -4506 81854 -4422
rect 81234 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 81854 -4506
rect 81234 -5734 81854 -4742
rect 66954 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 67574 -7066
rect 66954 -7386 67574 -7302
rect 66954 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 67574 -7386
rect 66954 -7654 67574 -7622
rect 84954 -6106 85574 -2000
rect 95514 -3226 96134 -2000
rect 95514 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 96134 -3226
rect 95514 -3546 96134 -3462
rect 95514 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 96134 -3546
rect 95514 -3814 96134 -3782
rect 99234 -5146 99854 -2000
rect 99234 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 99854 -5146
rect 99234 -5466 99854 -5382
rect 99234 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 99854 -5466
rect 99234 -5734 99854 -5702
rect 84954 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 85574 -6106
rect 84954 -6426 85574 -6342
rect 84954 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 85574 -6426
rect 84954 -7654 85574 -6662
rect 102954 -7066 103574 -2000
rect 113514 -2266 114134 -2000
rect 113514 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 114134 -2266
rect 113514 -2586 114134 -2502
rect 113514 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 114134 -2586
rect 113514 -3814 114134 -2822
rect 117234 -4186 117854 -2000
rect 117234 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 117854 -4186
rect 117234 -4506 117854 -4422
rect 117234 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 117854 -4506
rect 117234 -5734 117854 -4742
rect 102954 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 103574 -7066
rect 102954 -7386 103574 -7302
rect 102954 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 103574 -7386
rect 102954 -7654 103574 -7622
rect 120954 -6106 121574 -2000
rect 131514 -3226 132134 -2000
rect 131514 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 132134 -3226
rect 131514 -3546 132134 -3462
rect 131514 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 132134 -3546
rect 131514 -3814 132134 -3782
rect 135234 -5146 135854 -2000
rect 135234 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 135854 -5146
rect 135234 -5466 135854 -5382
rect 135234 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 135854 -5466
rect 135234 -5734 135854 -5702
rect 120954 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 121574 -6106
rect 120954 -6426 121574 -6342
rect 120954 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 121574 -6426
rect 120954 -7654 121574 -6662
rect 138954 -7066 139574 -2000
rect 149514 -2266 150134 -2000
rect 149514 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 150134 -2266
rect 149514 -2586 150134 -2502
rect 149514 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 150134 -2586
rect 149514 -3814 150134 -2822
rect 153234 -4186 153854 -2000
rect 153234 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 153854 -4186
rect 153234 -4506 153854 -4422
rect 153234 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 153854 -4506
rect 153234 -5734 153854 -4742
rect 138954 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 139574 -7066
rect 138954 -7386 139574 -7302
rect 138954 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 139574 -7386
rect 138954 -7654 139574 -7622
rect 156954 -6106 157574 -2000
rect 167514 -3226 168134 -2000
rect 167514 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 168134 -3226
rect 167514 -3546 168134 -3462
rect 167514 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 168134 -3546
rect 167514 -3814 168134 -3782
rect 171234 -5146 171854 -2000
rect 171234 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 171854 -5146
rect 171234 -5466 171854 -5382
rect 171234 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 171854 -5466
rect 171234 -5734 171854 -5702
rect 156954 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 157574 -6106
rect 156954 -6426 157574 -6342
rect 156954 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 157574 -6426
rect 156954 -7654 157574 -6662
rect 174954 -7066 175574 -2000
rect 185514 -2266 186134 -2000
rect 185514 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 186134 -2266
rect 185514 -2586 186134 -2502
rect 185514 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 186134 -2586
rect 185514 -3814 186134 -2822
rect 189234 -4186 189854 -2000
rect 189234 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 189854 -4186
rect 189234 -4506 189854 -4422
rect 189234 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 189854 -4506
rect 189234 -5734 189854 -4742
rect 174954 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 175574 -7066
rect 174954 -7386 175574 -7302
rect 174954 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 175574 -7386
rect 174954 -7654 175574 -7622
rect 192954 -6106 193574 -2000
rect 203514 -3226 204134 -2000
rect 203514 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 204134 -3226
rect 203514 -3546 204134 -3462
rect 203514 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 204134 -3546
rect 203514 -3814 204134 -3782
rect 207234 -5146 207854 -2000
rect 207234 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 207854 -5146
rect 207234 -5466 207854 -5382
rect 207234 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 207854 -5466
rect 207234 -5734 207854 -5702
rect 192954 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 193574 -6106
rect 192954 -6426 193574 -6342
rect 192954 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 193574 -6426
rect 192954 -7654 193574 -6662
rect 210954 -7066 211574 -2000
rect 221514 -2266 222134 -2000
rect 221514 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 222134 -2266
rect 221514 -2586 222134 -2502
rect 221514 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 222134 -2586
rect 221514 -3814 222134 -2822
rect 225234 -4186 225854 -2000
rect 225234 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 225854 -4186
rect 225234 -4506 225854 -4422
rect 225234 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 225854 -4506
rect 225234 -5734 225854 -4742
rect 210954 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 211574 -7066
rect 210954 -7386 211574 -7302
rect 210954 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 211574 -7386
rect 210954 -7654 211574 -7622
rect 228954 -6106 229574 -2000
rect 239514 -3226 240134 -2000
rect 239514 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 240134 -3226
rect 239514 -3546 240134 -3462
rect 239514 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 240134 -3546
rect 239514 -3814 240134 -3782
rect 243234 -5146 243854 -2000
rect 243234 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 243854 -5146
rect 243234 -5466 243854 -5382
rect 243234 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 243854 -5466
rect 243234 -5734 243854 -5702
rect 228954 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 229574 -6106
rect 228954 -6426 229574 -6342
rect 228954 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 229574 -6426
rect 228954 -7654 229574 -6662
rect 246954 -7066 247574 -2000
rect 257514 -2266 258134 -2000
rect 257514 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 258134 -2266
rect 257514 -2586 258134 -2502
rect 257514 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 258134 -2586
rect 257514 -3814 258134 -2822
rect 261234 -4186 261854 -2000
rect 261234 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 261854 -4186
rect 261234 -4506 261854 -4422
rect 261234 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 261854 -4506
rect 261234 -5734 261854 -4742
rect 246954 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 247574 -7066
rect 246954 -7386 247574 -7302
rect 246954 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 247574 -7386
rect 246954 -7654 247574 -7622
rect 264954 -6106 265574 -2000
rect 275514 -3226 276134 -2000
rect 275514 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 276134 -3226
rect 275514 -3546 276134 -3462
rect 275514 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 276134 -3546
rect 275514 -3814 276134 -3782
rect 279234 -5146 279854 -2000
rect 279234 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 279854 -5146
rect 279234 -5466 279854 -5382
rect 279234 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 279854 -5466
rect 279234 -5734 279854 -5702
rect 264954 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 265574 -6106
rect 264954 -6426 265574 -6342
rect 264954 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 265574 -6426
rect 264954 -7654 265574 -6662
rect 282954 -7066 283574 -2000
rect 293514 -2266 294134 -2000
rect 293514 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 294134 -2266
rect 293514 -2586 294134 -2502
rect 293514 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 294134 -2586
rect 293514 -3814 294134 -2822
rect 297234 -4186 297854 -2000
rect 297234 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 297854 -4186
rect 297234 -4506 297854 -4422
rect 297234 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 297854 -4506
rect 297234 -5734 297854 -4742
rect 282954 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 283574 -7066
rect 282954 -7386 283574 -7302
rect 282954 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 283574 -7386
rect 282954 -7654 283574 -7622
rect 300954 -6106 301574 -2000
rect 311514 -3226 312134 -2000
rect 311514 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 312134 -3226
rect 311514 -3546 312134 -3462
rect 311514 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 312134 -3546
rect 311514 -3814 312134 -3782
rect 315234 -5146 315854 -2000
rect 315234 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 315854 -5146
rect 315234 -5466 315854 -5382
rect 315234 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 315854 -5466
rect 315234 -5734 315854 -5702
rect 300954 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 301574 -6106
rect 300954 -6426 301574 -6342
rect 300954 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 301574 -6426
rect 300954 -7654 301574 -6662
rect 318954 -7066 319574 -2000
rect 329514 -2266 330134 -2000
rect 329514 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 330134 -2266
rect 329514 -2586 330134 -2502
rect 329514 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 330134 -2586
rect 329514 -3814 330134 -2822
rect 333234 -4186 333854 -2000
rect 333234 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 333854 -4186
rect 333234 -4506 333854 -4422
rect 333234 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 333854 -4506
rect 333234 -5734 333854 -4742
rect 318954 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 319574 -7066
rect 318954 -7386 319574 -7302
rect 318954 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 319574 -7386
rect 318954 -7654 319574 -7622
rect 336954 -6106 337574 -2000
rect 347514 -3226 348134 -2000
rect 347514 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 348134 -3226
rect 347514 -3546 348134 -3462
rect 347514 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 348134 -3546
rect 347514 -3814 348134 -3782
rect 351234 -5146 351854 -2000
rect 351234 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 351854 -5146
rect 351234 -5466 351854 -5382
rect 351234 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 351854 -5466
rect 351234 -5734 351854 -5702
rect 336954 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 337574 -6106
rect 336954 -6426 337574 -6342
rect 336954 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 337574 -6426
rect 336954 -7654 337574 -6662
rect 354954 -7066 355574 -2000
rect 365514 -2266 366134 -2000
rect 365514 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 366134 -2266
rect 365514 -2586 366134 -2502
rect 365514 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 366134 -2586
rect 365514 -3814 366134 -2822
rect 369234 -4186 369854 -2000
rect 369234 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 369854 -4186
rect 369234 -4506 369854 -4422
rect 369234 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 369854 -4506
rect 369234 -5734 369854 -4742
rect 354954 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 355574 -7066
rect 354954 -7386 355574 -7302
rect 354954 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 355574 -7386
rect 354954 -7654 355574 -7622
rect 372954 -6106 373574 -2000
rect 383514 -3226 384134 -2000
rect 383514 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 384134 -3226
rect 383514 -3546 384134 -3462
rect 383514 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 384134 -3546
rect 383514 -3814 384134 -3782
rect 387234 -5146 387854 -2000
rect 387234 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 387854 -5146
rect 387234 -5466 387854 -5382
rect 387234 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 387854 -5466
rect 387234 -5734 387854 -5702
rect 372954 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 373574 -6106
rect 372954 -6426 373574 -6342
rect 372954 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 373574 -6426
rect 372954 -7654 373574 -6662
rect 390954 -7066 391574 -2000
rect 401514 -2266 402134 -2000
rect 401514 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 402134 -2266
rect 401514 -2586 402134 -2502
rect 401514 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 402134 -2586
rect 401514 -3814 402134 -2822
rect 405234 -4186 405854 -2000
rect 405234 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 405854 -4186
rect 405234 -4506 405854 -4422
rect 405234 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 405854 -4506
rect 405234 -5734 405854 -4742
rect 390954 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 391574 -7066
rect 390954 -7386 391574 -7302
rect 390954 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 391574 -7386
rect 390954 -7654 391574 -7622
rect 408954 -6106 409574 -2000
rect 419514 -3226 420134 -2000
rect 419514 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 420134 -3226
rect 419514 -3546 420134 -3462
rect 419514 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 420134 -3546
rect 419514 -3814 420134 -3782
rect 423234 -5146 423854 -2000
rect 423234 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 423854 -5146
rect 423234 -5466 423854 -5382
rect 423234 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 423854 -5466
rect 423234 -5734 423854 -5702
rect 408954 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 409574 -6106
rect 408954 -6426 409574 -6342
rect 408954 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 409574 -6426
rect 408954 -7654 409574 -6662
rect 426954 -7066 427574 -2000
rect 437514 -2266 438134 -2000
rect 437514 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 438134 -2266
rect 437514 -2586 438134 -2502
rect 437514 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 438134 -2586
rect 437514 -3814 438134 -2822
rect 441234 -4186 441854 -2000
rect 441234 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 441854 -4186
rect 441234 -4506 441854 -4422
rect 441234 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 441854 -4506
rect 441234 -5734 441854 -4742
rect 426954 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 427574 -7066
rect 426954 -7386 427574 -7302
rect 426954 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 427574 -7386
rect 426954 -7654 427574 -7622
rect 444954 -6106 445574 -2000
rect 455514 -3226 456134 -2000
rect 455514 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 456134 -3226
rect 455514 -3546 456134 -3462
rect 455514 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 456134 -3546
rect 455514 -3814 456134 -3782
rect 459234 -5146 459854 -2000
rect 459234 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 459854 -5146
rect 459234 -5466 459854 -5382
rect 459234 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 459854 -5466
rect 459234 -5734 459854 -5702
rect 444954 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 445574 -6106
rect 444954 -6426 445574 -6342
rect 444954 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 445574 -6426
rect 444954 -7654 445574 -6662
rect 462954 -7066 463574 -2000
rect 473514 -2266 474134 -2000
rect 473514 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 474134 -2266
rect 473514 -2586 474134 -2502
rect 473514 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 474134 -2586
rect 473514 -3814 474134 -2822
rect 477234 -4186 477854 -2000
rect 477234 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 477854 -4186
rect 477234 -4506 477854 -4422
rect 477234 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 477854 -4506
rect 477234 -5734 477854 -4742
rect 462954 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 463574 -7066
rect 462954 -7386 463574 -7302
rect 462954 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 463574 -7386
rect 462954 -7654 463574 -7622
rect 480954 -6106 481574 -2000
rect 491514 -3226 492134 -2000
rect 491514 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 492134 -3226
rect 491514 -3546 492134 -3462
rect 491514 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 492134 -3546
rect 491514 -3814 492134 -3782
rect 495234 -5146 495854 -2000
rect 495234 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 495854 -5146
rect 495234 -5466 495854 -5382
rect 495234 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 495854 -5466
rect 495234 -5734 495854 -5702
rect 480954 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 481574 -6106
rect 480954 -6426 481574 -6342
rect 480954 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 481574 -6426
rect 480954 -7654 481574 -6662
rect 498954 -7066 499574 -2000
rect 509514 -2266 510134 -2000
rect 509514 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 510134 -2266
rect 509514 -2586 510134 -2502
rect 509514 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 510134 -2586
rect 509514 -3814 510134 -2822
rect 513234 -4186 513854 -2000
rect 513234 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 513854 -4186
rect 513234 -4506 513854 -4422
rect 513234 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 513854 -4506
rect 513234 -5734 513854 -4742
rect 498954 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 499574 -7066
rect 498954 -7386 499574 -7302
rect 498954 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 499574 -7386
rect 498954 -7654 499574 -7622
rect 516954 -6106 517574 -2000
rect 527514 -3226 528134 -2000
rect 527514 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 528134 -3226
rect 527514 -3546 528134 -3462
rect 527514 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 528134 -3546
rect 527514 -3814 528134 -3782
rect 531234 -5146 531854 -2000
rect 531234 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 531854 -5146
rect 531234 -5466 531854 -5382
rect 531234 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 531854 -5466
rect 531234 -5734 531854 -5702
rect 516954 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 517574 -6106
rect 516954 -6426 517574 -6342
rect 516954 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 517574 -6426
rect 516954 -7654 517574 -6662
rect 534954 -7066 535574 -2000
rect 545514 -2266 546134 -2000
rect 545514 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 546134 -2266
rect 545514 -2586 546134 -2502
rect 545514 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 546134 -2586
rect 545514 -3814 546134 -2822
rect 549234 -4186 549854 -2000
rect 549234 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 549854 -4186
rect 549234 -4506 549854 -4422
rect 549234 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 549854 -4506
rect 549234 -5734 549854 -4742
rect 534954 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 535574 -7066
rect 534954 -7386 535574 -7302
rect 534954 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 535574 -7386
rect 534954 -7654 535574 -7622
rect 552954 -6106 553574 -2000
rect 563514 -3226 564134 -2000
rect 563514 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 564134 -3226
rect 563514 -3546 564134 -3462
rect 563514 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 564134 -3546
rect 563514 -3814 564134 -3782
rect 567234 -5146 567854 28338
rect 567234 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 567854 -5146
rect 567234 -5466 567854 -5382
rect 567234 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 567854 -5466
rect 567234 -5734 567854 -5702
rect 570954 680614 571574 711002
rect 592030 711558 592650 711590
rect 592030 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect 592030 711238 592650 711322
rect 592030 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect 591070 710598 591690 710630
rect 591070 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect 591070 710278 591690 710362
rect 591070 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect 590110 709638 590730 709670
rect 590110 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect 590110 709318 590730 709402
rect 590110 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect 589150 708678 589770 708710
rect 589150 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect 589150 708358 589770 708442
rect 589150 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect 581514 706758 582134 707750
rect 588190 707718 588810 707750
rect 588190 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect 588190 707398 588810 707482
rect 588190 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect 581514 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 582134 706758
rect 581514 706438 582134 706522
rect 581514 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 582134 706438
rect 570954 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 571574 680614
rect 570954 680294 571574 680378
rect 570954 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 571574 680294
rect 570954 644614 571574 680058
rect 570954 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 571574 644614
rect 570954 644294 571574 644378
rect 570954 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 571574 644294
rect 570954 608614 571574 644058
rect 570954 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 571574 608614
rect 570954 608294 571574 608378
rect 570954 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 571574 608294
rect 570954 572614 571574 608058
rect 570954 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 571574 572614
rect 570954 572294 571574 572378
rect 570954 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 571574 572294
rect 570954 536614 571574 572058
rect 570954 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 571574 536614
rect 570954 536294 571574 536378
rect 570954 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 571574 536294
rect 570954 500614 571574 536058
rect 570954 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 571574 500614
rect 570954 500294 571574 500378
rect 570954 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 571574 500294
rect 570954 464614 571574 500058
rect 570954 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 571574 464614
rect 570954 464294 571574 464378
rect 570954 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 571574 464294
rect 570954 428614 571574 464058
rect 570954 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 571574 428614
rect 570954 428294 571574 428378
rect 570954 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 571574 428294
rect 570954 392614 571574 428058
rect 570954 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 571574 392614
rect 570954 392294 571574 392378
rect 570954 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 571574 392294
rect 570954 356614 571574 392058
rect 570954 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 571574 356614
rect 570954 356294 571574 356378
rect 570954 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 571574 356294
rect 570954 320614 571574 356058
rect 570954 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 571574 320614
rect 570954 320294 571574 320378
rect 570954 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 571574 320294
rect 570954 284614 571574 320058
rect 570954 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 571574 284614
rect 570954 284294 571574 284378
rect 570954 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 571574 284294
rect 570954 248614 571574 284058
rect 570954 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 571574 248614
rect 570954 248294 571574 248378
rect 570954 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 571574 248294
rect 570954 212614 571574 248058
rect 570954 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 571574 212614
rect 570954 212294 571574 212378
rect 570954 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 571574 212294
rect 570954 176614 571574 212058
rect 570954 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 571574 176614
rect 570954 176294 571574 176378
rect 570954 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 571574 176294
rect 570954 140614 571574 176058
rect 570954 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 571574 140614
rect 570954 140294 571574 140378
rect 570954 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 571574 140294
rect 570954 104614 571574 140058
rect 570954 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 571574 104614
rect 570954 104294 571574 104378
rect 570954 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 571574 104294
rect 570954 68614 571574 104058
rect 570954 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 571574 68614
rect 570954 68294 571574 68378
rect 570954 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 571574 68294
rect 570954 32614 571574 68058
rect 570954 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 571574 32614
rect 570954 32294 571574 32378
rect 570954 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 571574 32294
rect 552954 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 553574 -6106
rect 552954 -6426 553574 -6342
rect 552954 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 553574 -6426
rect 552954 -7654 553574 -6662
rect 570954 -7066 571574 32058
rect 577794 704838 578414 705830
rect 577794 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 578414 704838
rect 577794 704518 578414 704602
rect 577794 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 578414 704518
rect 577794 687454 578414 704282
rect 577794 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 578414 687454
rect 577794 687134 578414 687218
rect 577794 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 578414 687134
rect 577794 651454 578414 686898
rect 577794 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 578414 651454
rect 577794 651134 578414 651218
rect 577794 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 578414 651134
rect 577794 615454 578414 650898
rect 577794 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 578414 615454
rect 577794 615134 578414 615218
rect 577794 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 578414 615134
rect 577794 579454 578414 614898
rect 577794 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 578414 579454
rect 577794 579134 578414 579218
rect 577794 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 578414 579134
rect 577794 543454 578414 578898
rect 577794 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 578414 543454
rect 577794 543134 578414 543218
rect 577794 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 578414 543134
rect 577794 507454 578414 542898
rect 577794 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 578414 507454
rect 577794 507134 578414 507218
rect 577794 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 578414 507134
rect 577794 471454 578414 506898
rect 577794 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 578414 471454
rect 577794 471134 578414 471218
rect 577794 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 578414 471134
rect 577794 435454 578414 470898
rect 577794 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 578414 435454
rect 577794 435134 578414 435218
rect 577794 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 578414 435134
rect 577794 399454 578414 434898
rect 577794 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 578414 399454
rect 577794 399134 578414 399218
rect 577794 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 578414 399134
rect 577794 363454 578414 398898
rect 577794 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 578414 363454
rect 577794 363134 578414 363218
rect 577794 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 578414 363134
rect 577794 327454 578414 362898
rect 577794 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 578414 327454
rect 577794 327134 578414 327218
rect 577794 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 578414 327134
rect 577794 291454 578414 326898
rect 577794 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 578414 291454
rect 577794 291134 578414 291218
rect 577794 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 578414 291134
rect 577794 255454 578414 290898
rect 577794 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 578414 255454
rect 577794 255134 578414 255218
rect 577794 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 578414 255134
rect 577794 219454 578414 254898
rect 577794 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 578414 219454
rect 577794 219134 578414 219218
rect 577794 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 578414 219134
rect 577794 183454 578414 218898
rect 577794 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 578414 183454
rect 577794 183134 578414 183218
rect 577794 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 578414 183134
rect 577794 147454 578414 182898
rect 577794 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 578414 147454
rect 577794 147134 578414 147218
rect 577794 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 578414 147134
rect 577794 111454 578414 146898
rect 577794 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 578414 111454
rect 577794 111134 578414 111218
rect 577794 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 578414 111134
rect 577794 75454 578414 110898
rect 577794 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 578414 75454
rect 577794 75134 578414 75218
rect 577794 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 578414 75134
rect 577794 39454 578414 74898
rect 577794 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 578414 39454
rect 577794 39134 578414 39218
rect 577794 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 578414 39134
rect 577794 3454 578414 38898
rect 577794 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 578414 3454
rect 577794 3134 578414 3218
rect 577794 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 578414 3134
rect 577794 -346 578414 2898
rect 577794 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 578414 -346
rect 577794 -666 578414 -582
rect 577794 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 578414 -666
rect 577794 -1894 578414 -902
rect 581514 691174 582134 706202
rect 587230 706758 587850 706790
rect 587230 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect 587230 706438 587850 706522
rect 587230 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect 586270 705798 586890 705830
rect 586270 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect 586270 705478 586890 705562
rect 586270 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect 581514 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 582134 691174
rect 581514 690854 582134 690938
rect 581514 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 582134 690854
rect 581514 655174 582134 690618
rect 581514 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 582134 655174
rect 581514 654854 582134 654938
rect 581514 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 582134 654854
rect 581514 619174 582134 654618
rect 581514 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 582134 619174
rect 581514 618854 582134 618938
rect 581514 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 582134 618854
rect 581514 583174 582134 618618
rect 581514 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 582134 583174
rect 581514 582854 582134 582938
rect 581514 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 582134 582854
rect 581514 547174 582134 582618
rect 581514 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 582134 547174
rect 581514 546854 582134 546938
rect 581514 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 582134 546854
rect 581514 511174 582134 546618
rect 581514 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 582134 511174
rect 581514 510854 582134 510938
rect 581514 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 582134 510854
rect 581514 475174 582134 510618
rect 581514 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 582134 475174
rect 581514 474854 582134 474938
rect 581514 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 582134 474854
rect 581514 439174 582134 474618
rect 581514 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 582134 439174
rect 581514 438854 582134 438938
rect 581514 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 582134 438854
rect 581514 403174 582134 438618
rect 581514 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 582134 403174
rect 581514 402854 582134 402938
rect 581514 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 582134 402854
rect 581514 367174 582134 402618
rect 581514 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 582134 367174
rect 581514 366854 582134 366938
rect 581514 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 582134 366854
rect 581514 331174 582134 366618
rect 581514 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 582134 331174
rect 581514 330854 582134 330938
rect 581514 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 582134 330854
rect 581514 295174 582134 330618
rect 581514 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 582134 295174
rect 581514 294854 582134 294938
rect 581514 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 582134 294854
rect 581514 259174 582134 294618
rect 581514 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 582134 259174
rect 581514 258854 582134 258938
rect 581514 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 582134 258854
rect 581514 223174 582134 258618
rect 581514 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 582134 223174
rect 581514 222854 582134 222938
rect 581514 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 582134 222854
rect 581514 187174 582134 222618
rect 581514 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 582134 187174
rect 581514 186854 582134 186938
rect 581514 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 582134 186854
rect 581514 151174 582134 186618
rect 581514 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 582134 151174
rect 581514 150854 582134 150938
rect 581514 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 582134 150854
rect 581514 115174 582134 150618
rect 581514 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 582134 115174
rect 581514 114854 582134 114938
rect 581514 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 582134 114854
rect 581514 79174 582134 114618
rect 581514 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 582134 79174
rect 581514 78854 582134 78938
rect 581514 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 582134 78854
rect 581514 43174 582134 78618
rect 581514 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 582134 43174
rect 581514 42854 582134 42938
rect 581514 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 582134 42854
rect 581514 7174 582134 42618
rect 581514 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 582134 7174
rect 581514 6854 582134 6938
rect 581514 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 582134 6854
rect 581514 -2266 582134 6618
rect 585310 704838 585930 704870
rect 585310 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect 585310 704518 585930 704602
rect 585310 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect 585310 687454 585930 704282
rect 585310 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 585930 687454
rect 585310 687134 585930 687218
rect 585310 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 585930 687134
rect 585310 651454 585930 686898
rect 585310 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 585930 651454
rect 585310 651134 585930 651218
rect 585310 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 585930 651134
rect 585310 615454 585930 650898
rect 585310 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 585930 615454
rect 585310 615134 585930 615218
rect 585310 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 585930 615134
rect 585310 579454 585930 614898
rect 585310 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 585930 579454
rect 585310 579134 585930 579218
rect 585310 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 585930 579134
rect 585310 543454 585930 578898
rect 585310 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 585930 543454
rect 585310 543134 585930 543218
rect 585310 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 585930 543134
rect 585310 507454 585930 542898
rect 585310 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 585930 507454
rect 585310 507134 585930 507218
rect 585310 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 585930 507134
rect 585310 471454 585930 506898
rect 585310 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 585930 471454
rect 585310 471134 585930 471218
rect 585310 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 585930 471134
rect 585310 435454 585930 470898
rect 585310 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 585930 435454
rect 585310 435134 585930 435218
rect 585310 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 585930 435134
rect 585310 399454 585930 434898
rect 585310 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 585930 399454
rect 585310 399134 585930 399218
rect 585310 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 585930 399134
rect 585310 363454 585930 398898
rect 585310 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 585930 363454
rect 585310 363134 585930 363218
rect 585310 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 585930 363134
rect 585310 327454 585930 362898
rect 585310 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 585930 327454
rect 585310 327134 585930 327218
rect 585310 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 585930 327134
rect 585310 291454 585930 326898
rect 585310 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 585930 291454
rect 585310 291134 585930 291218
rect 585310 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 585930 291134
rect 585310 255454 585930 290898
rect 585310 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 585930 255454
rect 585310 255134 585930 255218
rect 585310 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 585930 255134
rect 585310 219454 585930 254898
rect 585310 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 585930 219454
rect 585310 219134 585930 219218
rect 585310 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 585930 219134
rect 585310 183454 585930 218898
rect 585310 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 585930 183454
rect 585310 183134 585930 183218
rect 585310 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 585930 183134
rect 585310 147454 585930 182898
rect 585310 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 585930 147454
rect 585310 147134 585930 147218
rect 585310 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 585930 147134
rect 585310 111454 585930 146898
rect 585310 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 585930 111454
rect 585310 111134 585930 111218
rect 585310 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 585930 111134
rect 585310 75454 585930 110898
rect 585310 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 585930 75454
rect 585310 75134 585930 75218
rect 585310 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 585930 75134
rect 585310 39454 585930 74898
rect 585310 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 585930 39454
rect 585310 39134 585930 39218
rect 585310 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 585930 39134
rect 585310 3454 585930 38898
rect 585310 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 585930 3454
rect 585310 3134 585930 3218
rect 585310 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 585930 3134
rect 585310 -346 585930 2898
rect 585310 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect 585310 -666 585930 -582
rect 585310 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect 585310 -934 585930 -902
rect 586270 669454 586890 705242
rect 586270 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect 586270 669134 586890 669218
rect 586270 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect 586270 633454 586890 668898
rect 586270 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect 586270 633134 586890 633218
rect 586270 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect 586270 597454 586890 632898
rect 586270 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect 586270 597134 586890 597218
rect 586270 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect 586270 561454 586890 596898
rect 586270 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect 586270 561134 586890 561218
rect 586270 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect 586270 525454 586890 560898
rect 586270 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect 586270 525134 586890 525218
rect 586270 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect 586270 489454 586890 524898
rect 586270 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect 586270 489134 586890 489218
rect 586270 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect 586270 453454 586890 488898
rect 586270 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect 586270 453134 586890 453218
rect 586270 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect 586270 417454 586890 452898
rect 586270 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect 586270 417134 586890 417218
rect 586270 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect 586270 381454 586890 416898
rect 586270 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect 586270 381134 586890 381218
rect 586270 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect 586270 345454 586890 380898
rect 586270 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect 586270 345134 586890 345218
rect 586270 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect 586270 309454 586890 344898
rect 586270 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect 586270 309134 586890 309218
rect 586270 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect 586270 273454 586890 308898
rect 586270 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect 586270 273134 586890 273218
rect 586270 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect 586270 237454 586890 272898
rect 586270 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect 586270 237134 586890 237218
rect 586270 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect 586270 201454 586890 236898
rect 586270 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect 586270 201134 586890 201218
rect 586270 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect 586270 165454 586890 200898
rect 586270 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect 586270 165134 586890 165218
rect 586270 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect 586270 129454 586890 164898
rect 586270 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect 586270 129134 586890 129218
rect 586270 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect 586270 93454 586890 128898
rect 586270 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect 586270 93134 586890 93218
rect 586270 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect 586270 57454 586890 92898
rect 586270 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect 586270 57134 586890 57218
rect 586270 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect 586270 21454 586890 56898
rect 586270 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect 586270 21134 586890 21218
rect 586270 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect 586270 -1306 586890 20898
rect 586270 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect 586270 -1626 586890 -1542
rect 586270 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect 586270 -1894 586890 -1862
rect 587230 691174 587850 706202
rect 587230 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 587850 691174
rect 587230 690854 587850 690938
rect 587230 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 587850 690854
rect 587230 655174 587850 690618
rect 587230 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 587850 655174
rect 587230 654854 587850 654938
rect 587230 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 587850 654854
rect 587230 619174 587850 654618
rect 587230 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 587850 619174
rect 587230 618854 587850 618938
rect 587230 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 587850 618854
rect 587230 583174 587850 618618
rect 587230 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 587850 583174
rect 587230 582854 587850 582938
rect 587230 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 587850 582854
rect 587230 547174 587850 582618
rect 587230 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 587850 547174
rect 587230 546854 587850 546938
rect 587230 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 587850 546854
rect 587230 511174 587850 546618
rect 587230 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 587850 511174
rect 587230 510854 587850 510938
rect 587230 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 587850 510854
rect 587230 475174 587850 510618
rect 587230 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 587850 475174
rect 587230 474854 587850 474938
rect 587230 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 587850 474854
rect 587230 439174 587850 474618
rect 587230 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 587850 439174
rect 587230 438854 587850 438938
rect 587230 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 587850 438854
rect 587230 403174 587850 438618
rect 587230 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 587850 403174
rect 587230 402854 587850 402938
rect 587230 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 587850 402854
rect 587230 367174 587850 402618
rect 587230 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 587850 367174
rect 587230 366854 587850 366938
rect 587230 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 587850 366854
rect 587230 331174 587850 366618
rect 587230 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 587850 331174
rect 587230 330854 587850 330938
rect 587230 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 587850 330854
rect 587230 295174 587850 330618
rect 587230 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 587850 295174
rect 587230 294854 587850 294938
rect 587230 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 587850 294854
rect 587230 259174 587850 294618
rect 587230 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 587850 259174
rect 587230 258854 587850 258938
rect 587230 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 587850 258854
rect 587230 223174 587850 258618
rect 587230 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 587850 223174
rect 587230 222854 587850 222938
rect 587230 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 587850 222854
rect 587230 187174 587850 222618
rect 587230 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 587850 187174
rect 587230 186854 587850 186938
rect 587230 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 587850 186854
rect 587230 151174 587850 186618
rect 587230 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 587850 151174
rect 587230 150854 587850 150938
rect 587230 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 587850 150854
rect 587230 115174 587850 150618
rect 587230 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 587850 115174
rect 587230 114854 587850 114938
rect 587230 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 587850 114854
rect 587230 79174 587850 114618
rect 587230 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 587850 79174
rect 587230 78854 587850 78938
rect 587230 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 587850 78854
rect 587230 43174 587850 78618
rect 587230 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 587850 43174
rect 587230 42854 587850 42938
rect 587230 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 587850 42854
rect 587230 7174 587850 42618
rect 587230 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 587850 7174
rect 587230 6854 587850 6938
rect 587230 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 587850 6854
rect 581514 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 582134 -2266
rect 581514 -2586 582134 -2502
rect 581514 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 582134 -2586
rect 581514 -3814 582134 -2822
rect 587230 -2266 587850 6618
rect 587230 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect 587230 -2586 587850 -2502
rect 587230 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect 587230 -2854 587850 -2822
rect 588190 673174 588810 707162
rect 588190 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect 588190 672854 588810 672938
rect 588190 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect 588190 637174 588810 672618
rect 588190 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect 588190 636854 588810 636938
rect 588190 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect 588190 601174 588810 636618
rect 588190 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect 588190 600854 588810 600938
rect 588190 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect 588190 565174 588810 600618
rect 588190 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect 588190 564854 588810 564938
rect 588190 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect 588190 529174 588810 564618
rect 588190 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect 588190 528854 588810 528938
rect 588190 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect 588190 493174 588810 528618
rect 588190 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect 588190 492854 588810 492938
rect 588190 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect 588190 457174 588810 492618
rect 588190 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect 588190 456854 588810 456938
rect 588190 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect 588190 421174 588810 456618
rect 588190 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect 588190 420854 588810 420938
rect 588190 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect 588190 385174 588810 420618
rect 588190 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect 588190 384854 588810 384938
rect 588190 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect 588190 349174 588810 384618
rect 588190 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect 588190 348854 588810 348938
rect 588190 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect 588190 313174 588810 348618
rect 588190 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect 588190 312854 588810 312938
rect 588190 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect 588190 277174 588810 312618
rect 588190 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect 588190 276854 588810 276938
rect 588190 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect 588190 241174 588810 276618
rect 588190 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect 588190 240854 588810 240938
rect 588190 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect 588190 205174 588810 240618
rect 588190 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect 588190 204854 588810 204938
rect 588190 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect 588190 169174 588810 204618
rect 588190 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect 588190 168854 588810 168938
rect 588190 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect 588190 133174 588810 168618
rect 588190 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect 588190 132854 588810 132938
rect 588190 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect 588190 97174 588810 132618
rect 588190 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect 588190 96854 588810 96938
rect 588190 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect 588190 61174 588810 96618
rect 588190 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect 588190 60854 588810 60938
rect 588190 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect 588190 25174 588810 60618
rect 588190 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect 588190 24854 588810 24938
rect 588190 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect 588190 -3226 588810 24618
rect 588190 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect 588190 -3546 588810 -3462
rect 588190 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect 588190 -3814 588810 -3782
rect 589150 694894 589770 708122
rect 589150 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 589770 694894
rect 589150 694574 589770 694658
rect 589150 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 589770 694574
rect 589150 658894 589770 694338
rect 589150 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 589770 658894
rect 589150 658574 589770 658658
rect 589150 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 589770 658574
rect 589150 622894 589770 658338
rect 589150 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 589770 622894
rect 589150 622574 589770 622658
rect 589150 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 589770 622574
rect 589150 586894 589770 622338
rect 589150 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 589770 586894
rect 589150 586574 589770 586658
rect 589150 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 589770 586574
rect 589150 550894 589770 586338
rect 589150 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 589770 550894
rect 589150 550574 589770 550658
rect 589150 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 589770 550574
rect 589150 514894 589770 550338
rect 589150 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 589770 514894
rect 589150 514574 589770 514658
rect 589150 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 589770 514574
rect 589150 478894 589770 514338
rect 589150 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 589770 478894
rect 589150 478574 589770 478658
rect 589150 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 589770 478574
rect 589150 442894 589770 478338
rect 589150 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 589770 442894
rect 589150 442574 589770 442658
rect 589150 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 589770 442574
rect 589150 406894 589770 442338
rect 589150 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 589770 406894
rect 589150 406574 589770 406658
rect 589150 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 589770 406574
rect 589150 370894 589770 406338
rect 589150 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 589770 370894
rect 589150 370574 589770 370658
rect 589150 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 589770 370574
rect 589150 334894 589770 370338
rect 589150 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 589770 334894
rect 589150 334574 589770 334658
rect 589150 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 589770 334574
rect 589150 298894 589770 334338
rect 589150 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 589770 298894
rect 589150 298574 589770 298658
rect 589150 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 589770 298574
rect 589150 262894 589770 298338
rect 589150 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 589770 262894
rect 589150 262574 589770 262658
rect 589150 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 589770 262574
rect 589150 226894 589770 262338
rect 589150 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 589770 226894
rect 589150 226574 589770 226658
rect 589150 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 589770 226574
rect 589150 190894 589770 226338
rect 589150 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 589770 190894
rect 589150 190574 589770 190658
rect 589150 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 589770 190574
rect 589150 154894 589770 190338
rect 589150 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 589770 154894
rect 589150 154574 589770 154658
rect 589150 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 589770 154574
rect 589150 118894 589770 154338
rect 589150 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 589770 118894
rect 589150 118574 589770 118658
rect 589150 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 589770 118574
rect 589150 82894 589770 118338
rect 589150 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 589770 82894
rect 589150 82574 589770 82658
rect 589150 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 589770 82574
rect 589150 46894 589770 82338
rect 589150 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 589770 46894
rect 589150 46574 589770 46658
rect 589150 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 589770 46574
rect 589150 10894 589770 46338
rect 589150 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 589770 10894
rect 589150 10574 589770 10658
rect 589150 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 589770 10574
rect 589150 -4186 589770 10338
rect 589150 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect 589150 -4506 589770 -4422
rect 589150 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect 589150 -4774 589770 -4742
rect 590110 676894 590730 709082
rect 590110 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect 590110 676574 590730 676658
rect 590110 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect 590110 640894 590730 676338
rect 590110 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect 590110 640574 590730 640658
rect 590110 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect 590110 604894 590730 640338
rect 590110 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect 590110 604574 590730 604658
rect 590110 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect 590110 568894 590730 604338
rect 590110 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect 590110 568574 590730 568658
rect 590110 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect 590110 532894 590730 568338
rect 590110 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect 590110 532574 590730 532658
rect 590110 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect 590110 496894 590730 532338
rect 590110 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect 590110 496574 590730 496658
rect 590110 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect 590110 460894 590730 496338
rect 590110 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect 590110 460574 590730 460658
rect 590110 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect 590110 424894 590730 460338
rect 590110 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect 590110 424574 590730 424658
rect 590110 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect 590110 388894 590730 424338
rect 590110 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect 590110 388574 590730 388658
rect 590110 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect 590110 352894 590730 388338
rect 590110 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect 590110 352574 590730 352658
rect 590110 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect 590110 316894 590730 352338
rect 590110 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect 590110 316574 590730 316658
rect 590110 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect 590110 280894 590730 316338
rect 590110 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect 590110 280574 590730 280658
rect 590110 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect 590110 244894 590730 280338
rect 590110 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect 590110 244574 590730 244658
rect 590110 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect 590110 208894 590730 244338
rect 590110 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect 590110 208574 590730 208658
rect 590110 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect 590110 172894 590730 208338
rect 590110 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect 590110 172574 590730 172658
rect 590110 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect 590110 136894 590730 172338
rect 590110 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect 590110 136574 590730 136658
rect 590110 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect 590110 100894 590730 136338
rect 590110 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect 590110 100574 590730 100658
rect 590110 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect 590110 64894 590730 100338
rect 590110 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect 590110 64574 590730 64658
rect 590110 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect 590110 28894 590730 64338
rect 590110 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect 590110 28574 590730 28658
rect 590110 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect 590110 -5146 590730 28338
rect 590110 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect 590110 -5466 590730 -5382
rect 590110 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect 590110 -5734 590730 -5702
rect 591070 698614 591690 710042
rect 591070 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 591690 698614
rect 591070 698294 591690 698378
rect 591070 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 591690 698294
rect 591070 662614 591690 698058
rect 591070 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 591690 662614
rect 591070 662294 591690 662378
rect 591070 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 591690 662294
rect 591070 626614 591690 662058
rect 591070 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 591690 626614
rect 591070 626294 591690 626378
rect 591070 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 591690 626294
rect 591070 590614 591690 626058
rect 591070 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 591690 590614
rect 591070 590294 591690 590378
rect 591070 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 591690 590294
rect 591070 554614 591690 590058
rect 591070 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 591690 554614
rect 591070 554294 591690 554378
rect 591070 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 591690 554294
rect 591070 518614 591690 554058
rect 591070 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 591690 518614
rect 591070 518294 591690 518378
rect 591070 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 591690 518294
rect 591070 482614 591690 518058
rect 591070 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 591690 482614
rect 591070 482294 591690 482378
rect 591070 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 591690 482294
rect 591070 446614 591690 482058
rect 591070 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 591690 446614
rect 591070 446294 591690 446378
rect 591070 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 591690 446294
rect 591070 410614 591690 446058
rect 591070 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 591690 410614
rect 591070 410294 591690 410378
rect 591070 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 591690 410294
rect 591070 374614 591690 410058
rect 591070 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 591690 374614
rect 591070 374294 591690 374378
rect 591070 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 591690 374294
rect 591070 338614 591690 374058
rect 591070 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 591690 338614
rect 591070 338294 591690 338378
rect 591070 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 591690 338294
rect 591070 302614 591690 338058
rect 591070 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 591690 302614
rect 591070 302294 591690 302378
rect 591070 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 591690 302294
rect 591070 266614 591690 302058
rect 591070 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 591690 266614
rect 591070 266294 591690 266378
rect 591070 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 591690 266294
rect 591070 230614 591690 266058
rect 591070 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 591690 230614
rect 591070 230294 591690 230378
rect 591070 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 591690 230294
rect 591070 194614 591690 230058
rect 591070 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 591690 194614
rect 591070 194294 591690 194378
rect 591070 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 591690 194294
rect 591070 158614 591690 194058
rect 591070 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 591690 158614
rect 591070 158294 591690 158378
rect 591070 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 591690 158294
rect 591070 122614 591690 158058
rect 591070 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 591690 122614
rect 591070 122294 591690 122378
rect 591070 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 591690 122294
rect 591070 86614 591690 122058
rect 591070 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 591690 86614
rect 591070 86294 591690 86378
rect 591070 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 591690 86294
rect 591070 50614 591690 86058
rect 591070 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 591690 50614
rect 591070 50294 591690 50378
rect 591070 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 591690 50294
rect 591070 14614 591690 50058
rect 591070 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 591690 14614
rect 591070 14294 591690 14378
rect 591070 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 591690 14294
rect 591070 -6106 591690 14058
rect 591070 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect 591070 -6426 591690 -6342
rect 591070 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect 591070 -6694 591690 -6662
rect 592030 680614 592650 711002
rect 592030 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect 592030 680294 592650 680378
rect 592030 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect 592030 644614 592650 680058
rect 592030 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect 592030 644294 592650 644378
rect 592030 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect 592030 608614 592650 644058
rect 592030 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect 592030 608294 592650 608378
rect 592030 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect 592030 572614 592650 608058
rect 592030 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect 592030 572294 592650 572378
rect 592030 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect 592030 536614 592650 572058
rect 592030 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect 592030 536294 592650 536378
rect 592030 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect 592030 500614 592650 536058
rect 592030 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect 592030 500294 592650 500378
rect 592030 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect 592030 464614 592650 500058
rect 592030 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect 592030 464294 592650 464378
rect 592030 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect 592030 428614 592650 464058
rect 592030 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect 592030 428294 592650 428378
rect 592030 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect 592030 392614 592650 428058
rect 592030 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect 592030 392294 592650 392378
rect 592030 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect 592030 356614 592650 392058
rect 592030 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect 592030 356294 592650 356378
rect 592030 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect 592030 320614 592650 356058
rect 592030 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect 592030 320294 592650 320378
rect 592030 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect 592030 284614 592650 320058
rect 592030 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect 592030 284294 592650 284378
rect 592030 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect 592030 248614 592650 284058
rect 592030 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect 592030 248294 592650 248378
rect 592030 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect 592030 212614 592650 248058
rect 592030 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect 592030 212294 592650 212378
rect 592030 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect 592030 176614 592650 212058
rect 592030 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect 592030 176294 592650 176378
rect 592030 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect 592030 140614 592650 176058
rect 592030 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect 592030 140294 592650 140378
rect 592030 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect 592030 104614 592650 140058
rect 592030 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect 592030 104294 592650 104378
rect 592030 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect 592030 68614 592650 104058
rect 592030 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect 592030 68294 592650 68378
rect 592030 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect 592030 32614 592650 68058
rect 592030 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect 592030 32294 592650 32378
rect 592030 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect 570954 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 571574 -7066
rect 570954 -7386 571574 -7302
rect 570954 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 571574 -7386
rect 570954 -7654 571574 -7622
rect 592030 -7066 592650 32058
rect 592030 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect 592030 -7386 592650 -7302
rect 592030 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect 592030 -7654 592650 -7622
<< via4 >>
rect -8694 711322 -8458 711558
rect -8374 711322 -8138 711558
rect -8694 711002 -8458 711238
rect -8374 711002 -8138 711238
rect -8694 680378 -8458 680614
rect -8374 680378 -8138 680614
rect -8694 680058 -8458 680294
rect -8374 680058 -8138 680294
rect -8694 644378 -8458 644614
rect -8374 644378 -8138 644614
rect -8694 644058 -8458 644294
rect -8374 644058 -8138 644294
rect -8694 608378 -8458 608614
rect -8374 608378 -8138 608614
rect -8694 608058 -8458 608294
rect -8374 608058 -8138 608294
rect -8694 572378 -8458 572614
rect -8374 572378 -8138 572614
rect -8694 572058 -8458 572294
rect -8374 572058 -8138 572294
rect -8694 536378 -8458 536614
rect -8374 536378 -8138 536614
rect -8694 536058 -8458 536294
rect -8374 536058 -8138 536294
rect -8694 500378 -8458 500614
rect -8374 500378 -8138 500614
rect -8694 500058 -8458 500294
rect -8374 500058 -8138 500294
rect -8694 464378 -8458 464614
rect -8374 464378 -8138 464614
rect -8694 464058 -8458 464294
rect -8374 464058 -8138 464294
rect -8694 428378 -8458 428614
rect -8374 428378 -8138 428614
rect -8694 428058 -8458 428294
rect -8374 428058 -8138 428294
rect -8694 392378 -8458 392614
rect -8374 392378 -8138 392614
rect -8694 392058 -8458 392294
rect -8374 392058 -8138 392294
rect -8694 356378 -8458 356614
rect -8374 356378 -8138 356614
rect -8694 356058 -8458 356294
rect -8374 356058 -8138 356294
rect -8694 320378 -8458 320614
rect -8374 320378 -8138 320614
rect -8694 320058 -8458 320294
rect -8374 320058 -8138 320294
rect -8694 284378 -8458 284614
rect -8374 284378 -8138 284614
rect -8694 284058 -8458 284294
rect -8374 284058 -8138 284294
rect -8694 248378 -8458 248614
rect -8374 248378 -8138 248614
rect -8694 248058 -8458 248294
rect -8374 248058 -8138 248294
rect -8694 212378 -8458 212614
rect -8374 212378 -8138 212614
rect -8694 212058 -8458 212294
rect -8374 212058 -8138 212294
rect -8694 176378 -8458 176614
rect -8374 176378 -8138 176614
rect -8694 176058 -8458 176294
rect -8374 176058 -8138 176294
rect -8694 140378 -8458 140614
rect -8374 140378 -8138 140614
rect -8694 140058 -8458 140294
rect -8374 140058 -8138 140294
rect -8694 104378 -8458 104614
rect -8374 104378 -8138 104614
rect -8694 104058 -8458 104294
rect -8374 104058 -8138 104294
rect -8694 68378 -8458 68614
rect -8374 68378 -8138 68614
rect -8694 68058 -8458 68294
rect -8374 68058 -8138 68294
rect -8694 32378 -8458 32614
rect -8374 32378 -8138 32614
rect -8694 32058 -8458 32294
rect -8374 32058 -8138 32294
rect -7734 710362 -7498 710598
rect -7414 710362 -7178 710598
rect -7734 710042 -7498 710278
rect -7414 710042 -7178 710278
rect 12986 710362 13222 710598
rect 13306 710362 13542 710598
rect 12986 710042 13222 710278
rect 13306 710042 13542 710278
rect -7734 698378 -7498 698614
rect -7414 698378 -7178 698614
rect -7734 698058 -7498 698294
rect -7414 698058 -7178 698294
rect -7734 662378 -7498 662614
rect -7414 662378 -7178 662614
rect -7734 662058 -7498 662294
rect -7414 662058 -7178 662294
rect -7734 626378 -7498 626614
rect -7414 626378 -7178 626614
rect -7734 626058 -7498 626294
rect -7414 626058 -7178 626294
rect -7734 590378 -7498 590614
rect -7414 590378 -7178 590614
rect -7734 590058 -7498 590294
rect -7414 590058 -7178 590294
rect -7734 554378 -7498 554614
rect -7414 554378 -7178 554614
rect -7734 554058 -7498 554294
rect -7414 554058 -7178 554294
rect -7734 518378 -7498 518614
rect -7414 518378 -7178 518614
rect -7734 518058 -7498 518294
rect -7414 518058 -7178 518294
rect -7734 482378 -7498 482614
rect -7414 482378 -7178 482614
rect -7734 482058 -7498 482294
rect -7414 482058 -7178 482294
rect -7734 446378 -7498 446614
rect -7414 446378 -7178 446614
rect -7734 446058 -7498 446294
rect -7414 446058 -7178 446294
rect -7734 410378 -7498 410614
rect -7414 410378 -7178 410614
rect -7734 410058 -7498 410294
rect -7414 410058 -7178 410294
rect -7734 374378 -7498 374614
rect -7414 374378 -7178 374614
rect -7734 374058 -7498 374294
rect -7414 374058 -7178 374294
rect -7734 338378 -7498 338614
rect -7414 338378 -7178 338614
rect -7734 338058 -7498 338294
rect -7414 338058 -7178 338294
rect -7734 302378 -7498 302614
rect -7414 302378 -7178 302614
rect -7734 302058 -7498 302294
rect -7414 302058 -7178 302294
rect -7734 266378 -7498 266614
rect -7414 266378 -7178 266614
rect -7734 266058 -7498 266294
rect -7414 266058 -7178 266294
rect -7734 230378 -7498 230614
rect -7414 230378 -7178 230614
rect -7734 230058 -7498 230294
rect -7414 230058 -7178 230294
rect -7734 194378 -7498 194614
rect -7414 194378 -7178 194614
rect -7734 194058 -7498 194294
rect -7414 194058 -7178 194294
rect -7734 158378 -7498 158614
rect -7414 158378 -7178 158614
rect -7734 158058 -7498 158294
rect -7414 158058 -7178 158294
rect -7734 122378 -7498 122614
rect -7414 122378 -7178 122614
rect -7734 122058 -7498 122294
rect -7414 122058 -7178 122294
rect -7734 86378 -7498 86614
rect -7414 86378 -7178 86614
rect -7734 86058 -7498 86294
rect -7414 86058 -7178 86294
rect -7734 50378 -7498 50614
rect -7414 50378 -7178 50614
rect -7734 50058 -7498 50294
rect -7414 50058 -7178 50294
rect -7734 14378 -7498 14614
rect -7414 14378 -7178 14614
rect -7734 14058 -7498 14294
rect -7414 14058 -7178 14294
rect -6774 709402 -6538 709638
rect -6454 709402 -6218 709638
rect -6774 709082 -6538 709318
rect -6454 709082 -6218 709318
rect -6774 676658 -6538 676894
rect -6454 676658 -6218 676894
rect -6774 676338 -6538 676574
rect -6454 676338 -6218 676574
rect -6774 640658 -6538 640894
rect -6454 640658 -6218 640894
rect -6774 640338 -6538 640574
rect -6454 640338 -6218 640574
rect -6774 604658 -6538 604894
rect -6454 604658 -6218 604894
rect -6774 604338 -6538 604574
rect -6454 604338 -6218 604574
rect -6774 568658 -6538 568894
rect -6454 568658 -6218 568894
rect -6774 568338 -6538 568574
rect -6454 568338 -6218 568574
rect -6774 532658 -6538 532894
rect -6454 532658 -6218 532894
rect -6774 532338 -6538 532574
rect -6454 532338 -6218 532574
rect -6774 496658 -6538 496894
rect -6454 496658 -6218 496894
rect -6774 496338 -6538 496574
rect -6454 496338 -6218 496574
rect -6774 460658 -6538 460894
rect -6454 460658 -6218 460894
rect -6774 460338 -6538 460574
rect -6454 460338 -6218 460574
rect -6774 424658 -6538 424894
rect -6454 424658 -6218 424894
rect -6774 424338 -6538 424574
rect -6454 424338 -6218 424574
rect -6774 388658 -6538 388894
rect -6454 388658 -6218 388894
rect -6774 388338 -6538 388574
rect -6454 388338 -6218 388574
rect -6774 352658 -6538 352894
rect -6454 352658 -6218 352894
rect -6774 352338 -6538 352574
rect -6454 352338 -6218 352574
rect -6774 316658 -6538 316894
rect -6454 316658 -6218 316894
rect -6774 316338 -6538 316574
rect -6454 316338 -6218 316574
rect -6774 280658 -6538 280894
rect -6454 280658 -6218 280894
rect -6774 280338 -6538 280574
rect -6454 280338 -6218 280574
rect -6774 244658 -6538 244894
rect -6454 244658 -6218 244894
rect -6774 244338 -6538 244574
rect -6454 244338 -6218 244574
rect -6774 208658 -6538 208894
rect -6454 208658 -6218 208894
rect -6774 208338 -6538 208574
rect -6454 208338 -6218 208574
rect -6774 172658 -6538 172894
rect -6454 172658 -6218 172894
rect -6774 172338 -6538 172574
rect -6454 172338 -6218 172574
rect -6774 136658 -6538 136894
rect -6454 136658 -6218 136894
rect -6774 136338 -6538 136574
rect -6454 136338 -6218 136574
rect -6774 100658 -6538 100894
rect -6454 100658 -6218 100894
rect -6774 100338 -6538 100574
rect -6454 100338 -6218 100574
rect -6774 64658 -6538 64894
rect -6454 64658 -6218 64894
rect -6774 64338 -6538 64574
rect -6454 64338 -6218 64574
rect -6774 28658 -6538 28894
rect -6454 28658 -6218 28894
rect -6774 28338 -6538 28574
rect -6454 28338 -6218 28574
rect -5814 708442 -5578 708678
rect -5494 708442 -5258 708678
rect -5814 708122 -5578 708358
rect -5494 708122 -5258 708358
rect 9266 708442 9502 708678
rect 9586 708442 9822 708678
rect 9266 708122 9502 708358
rect 9586 708122 9822 708358
rect -5814 694658 -5578 694894
rect -5494 694658 -5258 694894
rect -5814 694338 -5578 694574
rect -5494 694338 -5258 694574
rect -5814 658658 -5578 658894
rect -5494 658658 -5258 658894
rect -5814 658338 -5578 658574
rect -5494 658338 -5258 658574
rect -5814 622658 -5578 622894
rect -5494 622658 -5258 622894
rect -5814 622338 -5578 622574
rect -5494 622338 -5258 622574
rect -5814 586658 -5578 586894
rect -5494 586658 -5258 586894
rect -5814 586338 -5578 586574
rect -5494 586338 -5258 586574
rect -5814 550658 -5578 550894
rect -5494 550658 -5258 550894
rect -5814 550338 -5578 550574
rect -5494 550338 -5258 550574
rect -5814 514658 -5578 514894
rect -5494 514658 -5258 514894
rect -5814 514338 -5578 514574
rect -5494 514338 -5258 514574
rect -5814 478658 -5578 478894
rect -5494 478658 -5258 478894
rect -5814 478338 -5578 478574
rect -5494 478338 -5258 478574
rect -5814 442658 -5578 442894
rect -5494 442658 -5258 442894
rect -5814 442338 -5578 442574
rect -5494 442338 -5258 442574
rect -5814 406658 -5578 406894
rect -5494 406658 -5258 406894
rect -5814 406338 -5578 406574
rect -5494 406338 -5258 406574
rect -5814 370658 -5578 370894
rect -5494 370658 -5258 370894
rect -5814 370338 -5578 370574
rect -5494 370338 -5258 370574
rect -5814 334658 -5578 334894
rect -5494 334658 -5258 334894
rect -5814 334338 -5578 334574
rect -5494 334338 -5258 334574
rect -5814 298658 -5578 298894
rect -5494 298658 -5258 298894
rect -5814 298338 -5578 298574
rect -5494 298338 -5258 298574
rect -5814 262658 -5578 262894
rect -5494 262658 -5258 262894
rect -5814 262338 -5578 262574
rect -5494 262338 -5258 262574
rect -5814 226658 -5578 226894
rect -5494 226658 -5258 226894
rect -5814 226338 -5578 226574
rect -5494 226338 -5258 226574
rect -5814 190658 -5578 190894
rect -5494 190658 -5258 190894
rect -5814 190338 -5578 190574
rect -5494 190338 -5258 190574
rect -5814 154658 -5578 154894
rect -5494 154658 -5258 154894
rect -5814 154338 -5578 154574
rect -5494 154338 -5258 154574
rect -5814 118658 -5578 118894
rect -5494 118658 -5258 118894
rect -5814 118338 -5578 118574
rect -5494 118338 -5258 118574
rect -5814 82658 -5578 82894
rect -5494 82658 -5258 82894
rect -5814 82338 -5578 82574
rect -5494 82338 -5258 82574
rect -5814 46658 -5578 46894
rect -5494 46658 -5258 46894
rect -5814 46338 -5578 46574
rect -5494 46338 -5258 46574
rect -5814 10658 -5578 10894
rect -5494 10658 -5258 10894
rect -5814 10338 -5578 10574
rect -5494 10338 -5258 10574
rect -4854 707482 -4618 707718
rect -4534 707482 -4298 707718
rect -4854 707162 -4618 707398
rect -4534 707162 -4298 707398
rect -4854 672938 -4618 673174
rect -4534 672938 -4298 673174
rect -4854 672618 -4618 672854
rect -4534 672618 -4298 672854
rect -4854 636938 -4618 637174
rect -4534 636938 -4298 637174
rect -4854 636618 -4618 636854
rect -4534 636618 -4298 636854
rect -4854 600938 -4618 601174
rect -4534 600938 -4298 601174
rect -4854 600618 -4618 600854
rect -4534 600618 -4298 600854
rect -4854 564938 -4618 565174
rect -4534 564938 -4298 565174
rect -4854 564618 -4618 564854
rect -4534 564618 -4298 564854
rect -4854 528938 -4618 529174
rect -4534 528938 -4298 529174
rect -4854 528618 -4618 528854
rect -4534 528618 -4298 528854
rect -4854 492938 -4618 493174
rect -4534 492938 -4298 493174
rect -4854 492618 -4618 492854
rect -4534 492618 -4298 492854
rect -4854 456938 -4618 457174
rect -4534 456938 -4298 457174
rect -4854 456618 -4618 456854
rect -4534 456618 -4298 456854
rect -4854 420938 -4618 421174
rect -4534 420938 -4298 421174
rect -4854 420618 -4618 420854
rect -4534 420618 -4298 420854
rect -4854 384938 -4618 385174
rect -4534 384938 -4298 385174
rect -4854 384618 -4618 384854
rect -4534 384618 -4298 384854
rect -4854 348938 -4618 349174
rect -4534 348938 -4298 349174
rect -4854 348618 -4618 348854
rect -4534 348618 -4298 348854
rect -4854 312938 -4618 313174
rect -4534 312938 -4298 313174
rect -4854 312618 -4618 312854
rect -4534 312618 -4298 312854
rect -4854 276938 -4618 277174
rect -4534 276938 -4298 277174
rect -4854 276618 -4618 276854
rect -4534 276618 -4298 276854
rect -4854 240938 -4618 241174
rect -4534 240938 -4298 241174
rect -4854 240618 -4618 240854
rect -4534 240618 -4298 240854
rect -4854 204938 -4618 205174
rect -4534 204938 -4298 205174
rect -4854 204618 -4618 204854
rect -4534 204618 -4298 204854
rect -4854 168938 -4618 169174
rect -4534 168938 -4298 169174
rect -4854 168618 -4618 168854
rect -4534 168618 -4298 168854
rect -4854 132938 -4618 133174
rect -4534 132938 -4298 133174
rect -4854 132618 -4618 132854
rect -4534 132618 -4298 132854
rect -4854 96938 -4618 97174
rect -4534 96938 -4298 97174
rect -4854 96618 -4618 96854
rect -4534 96618 -4298 96854
rect -4854 60938 -4618 61174
rect -4534 60938 -4298 61174
rect -4854 60618 -4618 60854
rect -4534 60618 -4298 60854
rect -4854 24938 -4618 25174
rect -4534 24938 -4298 25174
rect -4854 24618 -4618 24854
rect -4534 24618 -4298 24854
rect -3894 706522 -3658 706758
rect -3574 706522 -3338 706758
rect -3894 706202 -3658 706438
rect -3574 706202 -3338 706438
rect 5546 706522 5782 706758
rect 5866 706522 6102 706758
rect 5546 706202 5782 706438
rect 5866 706202 6102 706438
rect -3894 690938 -3658 691174
rect -3574 690938 -3338 691174
rect -3894 690618 -3658 690854
rect -3574 690618 -3338 690854
rect -3894 654938 -3658 655174
rect -3574 654938 -3338 655174
rect -3894 654618 -3658 654854
rect -3574 654618 -3338 654854
rect -3894 618938 -3658 619174
rect -3574 618938 -3338 619174
rect -3894 618618 -3658 618854
rect -3574 618618 -3338 618854
rect -3894 582938 -3658 583174
rect -3574 582938 -3338 583174
rect -3894 582618 -3658 582854
rect -3574 582618 -3338 582854
rect -3894 546938 -3658 547174
rect -3574 546938 -3338 547174
rect -3894 546618 -3658 546854
rect -3574 546618 -3338 546854
rect -3894 510938 -3658 511174
rect -3574 510938 -3338 511174
rect -3894 510618 -3658 510854
rect -3574 510618 -3338 510854
rect -3894 474938 -3658 475174
rect -3574 474938 -3338 475174
rect -3894 474618 -3658 474854
rect -3574 474618 -3338 474854
rect -3894 438938 -3658 439174
rect -3574 438938 -3338 439174
rect -3894 438618 -3658 438854
rect -3574 438618 -3338 438854
rect -3894 402938 -3658 403174
rect -3574 402938 -3338 403174
rect -3894 402618 -3658 402854
rect -3574 402618 -3338 402854
rect -3894 366938 -3658 367174
rect -3574 366938 -3338 367174
rect -3894 366618 -3658 366854
rect -3574 366618 -3338 366854
rect -3894 330938 -3658 331174
rect -3574 330938 -3338 331174
rect -3894 330618 -3658 330854
rect -3574 330618 -3338 330854
rect -3894 294938 -3658 295174
rect -3574 294938 -3338 295174
rect -3894 294618 -3658 294854
rect -3574 294618 -3338 294854
rect -3894 258938 -3658 259174
rect -3574 258938 -3338 259174
rect -3894 258618 -3658 258854
rect -3574 258618 -3338 258854
rect -3894 222938 -3658 223174
rect -3574 222938 -3338 223174
rect -3894 222618 -3658 222854
rect -3574 222618 -3338 222854
rect -3894 186938 -3658 187174
rect -3574 186938 -3338 187174
rect -3894 186618 -3658 186854
rect -3574 186618 -3338 186854
rect -3894 150938 -3658 151174
rect -3574 150938 -3338 151174
rect -3894 150618 -3658 150854
rect -3574 150618 -3338 150854
rect -3894 114938 -3658 115174
rect -3574 114938 -3338 115174
rect -3894 114618 -3658 114854
rect -3574 114618 -3338 114854
rect -3894 78938 -3658 79174
rect -3574 78938 -3338 79174
rect -3894 78618 -3658 78854
rect -3574 78618 -3338 78854
rect -3894 42938 -3658 43174
rect -3574 42938 -3338 43174
rect -3894 42618 -3658 42854
rect -3574 42618 -3338 42854
rect -3894 6938 -3658 7174
rect -3574 6938 -3338 7174
rect -3894 6618 -3658 6854
rect -3574 6618 -3338 6854
rect -2934 705562 -2698 705798
rect -2614 705562 -2378 705798
rect -2934 705242 -2698 705478
rect -2614 705242 -2378 705478
rect -2934 669218 -2698 669454
rect -2614 669218 -2378 669454
rect -2934 668898 -2698 669134
rect -2614 668898 -2378 669134
rect -2934 633218 -2698 633454
rect -2614 633218 -2378 633454
rect -2934 632898 -2698 633134
rect -2614 632898 -2378 633134
rect -2934 597218 -2698 597454
rect -2614 597218 -2378 597454
rect -2934 596898 -2698 597134
rect -2614 596898 -2378 597134
rect -2934 561218 -2698 561454
rect -2614 561218 -2378 561454
rect -2934 560898 -2698 561134
rect -2614 560898 -2378 561134
rect -2934 525218 -2698 525454
rect -2614 525218 -2378 525454
rect -2934 524898 -2698 525134
rect -2614 524898 -2378 525134
rect -2934 489218 -2698 489454
rect -2614 489218 -2378 489454
rect -2934 488898 -2698 489134
rect -2614 488898 -2378 489134
rect -2934 453218 -2698 453454
rect -2614 453218 -2378 453454
rect -2934 452898 -2698 453134
rect -2614 452898 -2378 453134
rect -2934 417218 -2698 417454
rect -2614 417218 -2378 417454
rect -2934 416898 -2698 417134
rect -2614 416898 -2378 417134
rect -2934 381218 -2698 381454
rect -2614 381218 -2378 381454
rect -2934 380898 -2698 381134
rect -2614 380898 -2378 381134
rect -2934 345218 -2698 345454
rect -2614 345218 -2378 345454
rect -2934 344898 -2698 345134
rect -2614 344898 -2378 345134
rect -2934 309218 -2698 309454
rect -2614 309218 -2378 309454
rect -2934 308898 -2698 309134
rect -2614 308898 -2378 309134
rect -2934 273218 -2698 273454
rect -2614 273218 -2378 273454
rect -2934 272898 -2698 273134
rect -2614 272898 -2378 273134
rect -2934 237218 -2698 237454
rect -2614 237218 -2378 237454
rect -2934 236898 -2698 237134
rect -2614 236898 -2378 237134
rect -2934 201218 -2698 201454
rect -2614 201218 -2378 201454
rect -2934 200898 -2698 201134
rect -2614 200898 -2378 201134
rect -2934 165218 -2698 165454
rect -2614 165218 -2378 165454
rect -2934 164898 -2698 165134
rect -2614 164898 -2378 165134
rect -2934 129218 -2698 129454
rect -2614 129218 -2378 129454
rect -2934 128898 -2698 129134
rect -2614 128898 -2378 129134
rect -2934 93218 -2698 93454
rect -2614 93218 -2378 93454
rect -2934 92898 -2698 93134
rect -2614 92898 -2378 93134
rect -2934 57218 -2698 57454
rect -2614 57218 -2378 57454
rect -2934 56898 -2698 57134
rect -2614 56898 -2378 57134
rect -2934 21218 -2698 21454
rect -2614 21218 -2378 21454
rect -2934 20898 -2698 21134
rect -2614 20898 -2378 21134
rect -1974 704602 -1738 704838
rect -1654 704602 -1418 704838
rect -1974 704282 -1738 704518
rect -1654 704282 -1418 704518
rect 1826 704602 2062 704838
rect 2146 704602 2382 704838
rect 1826 704282 2062 704518
rect 2146 704282 2382 704518
rect 30986 711322 31222 711558
rect 31306 711322 31542 711558
rect 30986 711002 31222 711238
rect 31306 711002 31542 711238
rect 27266 709402 27502 709638
rect 27586 709402 27822 709638
rect 27266 709082 27502 709318
rect 27586 709082 27822 709318
rect 23546 707482 23782 707718
rect 23866 707482 24102 707718
rect 23546 707162 23782 707398
rect 23866 707162 24102 707398
rect 19826 705562 20062 705798
rect 20146 705562 20382 705798
rect 19826 705242 20062 705478
rect 20146 705242 20382 705478
rect 48986 710362 49222 710598
rect 49306 710362 49542 710598
rect 48986 710042 49222 710278
rect 49306 710042 49542 710278
rect 45266 708442 45502 708678
rect 45586 708442 45822 708678
rect 45266 708122 45502 708358
rect 45586 708122 45822 708358
rect 41546 706522 41782 706758
rect 41866 706522 42102 706758
rect 41546 706202 41782 706438
rect 41866 706202 42102 706438
rect 37826 704602 38062 704838
rect 38146 704602 38382 704838
rect 37826 704282 38062 704518
rect 38146 704282 38382 704518
rect 66986 711322 67222 711558
rect 67306 711322 67542 711558
rect 66986 711002 67222 711238
rect 67306 711002 67542 711238
rect 63266 709402 63502 709638
rect 63586 709402 63822 709638
rect 63266 709082 63502 709318
rect 63586 709082 63822 709318
rect 59546 707482 59782 707718
rect 59866 707482 60102 707718
rect 59546 707162 59782 707398
rect 59866 707162 60102 707398
rect 55826 705562 56062 705798
rect 56146 705562 56382 705798
rect 55826 705242 56062 705478
rect 56146 705242 56382 705478
rect 84986 710362 85222 710598
rect 85306 710362 85542 710598
rect 84986 710042 85222 710278
rect 85306 710042 85542 710278
rect 81266 708442 81502 708678
rect 81586 708442 81822 708678
rect 81266 708122 81502 708358
rect 81586 708122 81822 708358
rect 77546 706522 77782 706758
rect 77866 706522 78102 706758
rect 77546 706202 77782 706438
rect 77866 706202 78102 706438
rect 73826 704602 74062 704838
rect 74146 704602 74382 704838
rect 73826 704282 74062 704518
rect 74146 704282 74382 704518
rect 102986 711322 103222 711558
rect 103306 711322 103542 711558
rect 102986 711002 103222 711238
rect 103306 711002 103542 711238
rect 99266 709402 99502 709638
rect 99586 709402 99822 709638
rect 99266 709082 99502 709318
rect 99586 709082 99822 709318
rect 95546 707482 95782 707718
rect 95866 707482 96102 707718
rect 95546 707162 95782 707398
rect 95866 707162 96102 707398
rect 91826 705562 92062 705798
rect 92146 705562 92382 705798
rect 91826 705242 92062 705478
rect 92146 705242 92382 705478
rect 120986 710362 121222 710598
rect 121306 710362 121542 710598
rect 120986 710042 121222 710278
rect 121306 710042 121542 710278
rect 117266 708442 117502 708678
rect 117586 708442 117822 708678
rect 117266 708122 117502 708358
rect 117586 708122 117822 708358
rect 113546 706522 113782 706758
rect 113866 706522 114102 706758
rect 113546 706202 113782 706438
rect 113866 706202 114102 706438
rect 109826 704602 110062 704838
rect 110146 704602 110382 704838
rect 109826 704282 110062 704518
rect 110146 704282 110382 704518
rect 138986 711322 139222 711558
rect 139306 711322 139542 711558
rect 138986 711002 139222 711238
rect 139306 711002 139542 711238
rect 135266 709402 135502 709638
rect 135586 709402 135822 709638
rect 135266 709082 135502 709318
rect 135586 709082 135822 709318
rect 131546 707482 131782 707718
rect 131866 707482 132102 707718
rect 131546 707162 131782 707398
rect 131866 707162 132102 707398
rect 127826 705562 128062 705798
rect 128146 705562 128382 705798
rect 127826 705242 128062 705478
rect 128146 705242 128382 705478
rect 156986 710362 157222 710598
rect 157306 710362 157542 710598
rect 156986 710042 157222 710278
rect 157306 710042 157542 710278
rect 153266 708442 153502 708678
rect 153586 708442 153822 708678
rect 153266 708122 153502 708358
rect 153586 708122 153822 708358
rect 149546 706522 149782 706758
rect 149866 706522 150102 706758
rect 149546 706202 149782 706438
rect 149866 706202 150102 706438
rect 145826 704602 146062 704838
rect 146146 704602 146382 704838
rect 145826 704282 146062 704518
rect 146146 704282 146382 704518
rect 174986 711322 175222 711558
rect 175306 711322 175542 711558
rect 174986 711002 175222 711238
rect 175306 711002 175542 711238
rect 171266 709402 171502 709638
rect 171586 709402 171822 709638
rect 171266 709082 171502 709318
rect 171586 709082 171822 709318
rect 167546 707482 167782 707718
rect 167866 707482 168102 707718
rect 167546 707162 167782 707398
rect 167866 707162 168102 707398
rect 163826 705562 164062 705798
rect 164146 705562 164382 705798
rect 163826 705242 164062 705478
rect 164146 705242 164382 705478
rect 192986 710362 193222 710598
rect 193306 710362 193542 710598
rect 192986 710042 193222 710278
rect 193306 710042 193542 710278
rect 189266 708442 189502 708678
rect 189586 708442 189822 708678
rect 189266 708122 189502 708358
rect 189586 708122 189822 708358
rect 185546 706522 185782 706758
rect 185866 706522 186102 706758
rect 185546 706202 185782 706438
rect 185866 706202 186102 706438
rect 181826 704602 182062 704838
rect 182146 704602 182382 704838
rect 181826 704282 182062 704518
rect 182146 704282 182382 704518
rect 210986 711322 211222 711558
rect 211306 711322 211542 711558
rect 210986 711002 211222 711238
rect 211306 711002 211542 711238
rect 207266 709402 207502 709638
rect 207586 709402 207822 709638
rect 207266 709082 207502 709318
rect 207586 709082 207822 709318
rect 203546 707482 203782 707718
rect 203866 707482 204102 707718
rect 203546 707162 203782 707398
rect 203866 707162 204102 707398
rect 199826 705562 200062 705798
rect 200146 705562 200382 705798
rect 199826 705242 200062 705478
rect 200146 705242 200382 705478
rect 228986 710362 229222 710598
rect 229306 710362 229542 710598
rect 228986 710042 229222 710278
rect 229306 710042 229542 710278
rect 225266 708442 225502 708678
rect 225586 708442 225822 708678
rect 225266 708122 225502 708358
rect 225586 708122 225822 708358
rect 221546 706522 221782 706758
rect 221866 706522 222102 706758
rect 221546 706202 221782 706438
rect 221866 706202 222102 706438
rect 217826 704602 218062 704838
rect 218146 704602 218382 704838
rect 217826 704282 218062 704518
rect 218146 704282 218382 704518
rect 246986 711322 247222 711558
rect 247306 711322 247542 711558
rect 246986 711002 247222 711238
rect 247306 711002 247542 711238
rect 243266 709402 243502 709638
rect 243586 709402 243822 709638
rect 243266 709082 243502 709318
rect 243586 709082 243822 709318
rect 239546 707482 239782 707718
rect 239866 707482 240102 707718
rect 239546 707162 239782 707398
rect 239866 707162 240102 707398
rect 235826 705562 236062 705798
rect 236146 705562 236382 705798
rect 235826 705242 236062 705478
rect 236146 705242 236382 705478
rect 264986 710362 265222 710598
rect 265306 710362 265542 710598
rect 264986 710042 265222 710278
rect 265306 710042 265542 710278
rect 261266 708442 261502 708678
rect 261586 708442 261822 708678
rect 261266 708122 261502 708358
rect 261586 708122 261822 708358
rect 257546 706522 257782 706758
rect 257866 706522 258102 706758
rect 257546 706202 257782 706438
rect 257866 706202 258102 706438
rect 253826 704602 254062 704838
rect 254146 704602 254382 704838
rect 253826 704282 254062 704518
rect 254146 704282 254382 704518
rect 282986 711322 283222 711558
rect 283306 711322 283542 711558
rect 282986 711002 283222 711238
rect 283306 711002 283542 711238
rect 279266 709402 279502 709638
rect 279586 709402 279822 709638
rect 279266 709082 279502 709318
rect 279586 709082 279822 709318
rect 275546 707482 275782 707718
rect 275866 707482 276102 707718
rect 275546 707162 275782 707398
rect 275866 707162 276102 707398
rect 271826 705562 272062 705798
rect 272146 705562 272382 705798
rect 271826 705242 272062 705478
rect 272146 705242 272382 705478
rect 300986 710362 301222 710598
rect 301306 710362 301542 710598
rect 300986 710042 301222 710278
rect 301306 710042 301542 710278
rect 297266 708442 297502 708678
rect 297586 708442 297822 708678
rect 297266 708122 297502 708358
rect 297586 708122 297822 708358
rect 293546 706522 293782 706758
rect 293866 706522 294102 706758
rect 293546 706202 293782 706438
rect 293866 706202 294102 706438
rect 289826 704602 290062 704838
rect 290146 704602 290382 704838
rect 289826 704282 290062 704518
rect 290146 704282 290382 704518
rect 318986 711322 319222 711558
rect 319306 711322 319542 711558
rect 318986 711002 319222 711238
rect 319306 711002 319542 711238
rect 315266 709402 315502 709638
rect 315586 709402 315822 709638
rect 315266 709082 315502 709318
rect 315586 709082 315822 709318
rect 311546 707482 311782 707718
rect 311866 707482 312102 707718
rect 311546 707162 311782 707398
rect 311866 707162 312102 707398
rect 307826 705562 308062 705798
rect 308146 705562 308382 705798
rect 307826 705242 308062 705478
rect 308146 705242 308382 705478
rect 336986 710362 337222 710598
rect 337306 710362 337542 710598
rect 336986 710042 337222 710278
rect 337306 710042 337542 710278
rect 333266 708442 333502 708678
rect 333586 708442 333822 708678
rect 333266 708122 333502 708358
rect 333586 708122 333822 708358
rect 329546 706522 329782 706758
rect 329866 706522 330102 706758
rect 329546 706202 329782 706438
rect 329866 706202 330102 706438
rect 325826 704602 326062 704838
rect 326146 704602 326382 704838
rect 325826 704282 326062 704518
rect 326146 704282 326382 704518
rect 354986 711322 355222 711558
rect 355306 711322 355542 711558
rect 354986 711002 355222 711238
rect 355306 711002 355542 711238
rect 351266 709402 351502 709638
rect 351586 709402 351822 709638
rect 351266 709082 351502 709318
rect 351586 709082 351822 709318
rect 347546 707482 347782 707718
rect 347866 707482 348102 707718
rect 347546 707162 347782 707398
rect 347866 707162 348102 707398
rect 343826 705562 344062 705798
rect 344146 705562 344382 705798
rect 343826 705242 344062 705478
rect 344146 705242 344382 705478
rect 372986 710362 373222 710598
rect 373306 710362 373542 710598
rect 372986 710042 373222 710278
rect 373306 710042 373542 710278
rect 369266 708442 369502 708678
rect 369586 708442 369822 708678
rect 369266 708122 369502 708358
rect 369586 708122 369822 708358
rect 365546 706522 365782 706758
rect 365866 706522 366102 706758
rect 365546 706202 365782 706438
rect 365866 706202 366102 706438
rect 361826 704602 362062 704838
rect 362146 704602 362382 704838
rect 361826 704282 362062 704518
rect 362146 704282 362382 704518
rect 390986 711322 391222 711558
rect 391306 711322 391542 711558
rect 390986 711002 391222 711238
rect 391306 711002 391542 711238
rect 387266 709402 387502 709638
rect 387586 709402 387822 709638
rect 387266 709082 387502 709318
rect 387586 709082 387822 709318
rect 383546 707482 383782 707718
rect 383866 707482 384102 707718
rect 383546 707162 383782 707398
rect 383866 707162 384102 707398
rect 379826 705562 380062 705798
rect 380146 705562 380382 705798
rect 379826 705242 380062 705478
rect 380146 705242 380382 705478
rect 408986 710362 409222 710598
rect 409306 710362 409542 710598
rect 408986 710042 409222 710278
rect 409306 710042 409542 710278
rect 405266 708442 405502 708678
rect 405586 708442 405822 708678
rect 405266 708122 405502 708358
rect 405586 708122 405822 708358
rect 401546 706522 401782 706758
rect 401866 706522 402102 706758
rect 401546 706202 401782 706438
rect 401866 706202 402102 706438
rect 397826 704602 398062 704838
rect 398146 704602 398382 704838
rect 397826 704282 398062 704518
rect 398146 704282 398382 704518
rect 426986 711322 427222 711558
rect 427306 711322 427542 711558
rect 426986 711002 427222 711238
rect 427306 711002 427542 711238
rect 423266 709402 423502 709638
rect 423586 709402 423822 709638
rect 423266 709082 423502 709318
rect 423586 709082 423822 709318
rect 419546 707482 419782 707718
rect 419866 707482 420102 707718
rect 419546 707162 419782 707398
rect 419866 707162 420102 707398
rect 415826 705562 416062 705798
rect 416146 705562 416382 705798
rect 415826 705242 416062 705478
rect 416146 705242 416382 705478
rect 444986 710362 445222 710598
rect 445306 710362 445542 710598
rect 444986 710042 445222 710278
rect 445306 710042 445542 710278
rect 441266 708442 441502 708678
rect 441586 708442 441822 708678
rect 441266 708122 441502 708358
rect 441586 708122 441822 708358
rect 437546 706522 437782 706758
rect 437866 706522 438102 706758
rect 437546 706202 437782 706438
rect 437866 706202 438102 706438
rect 433826 704602 434062 704838
rect 434146 704602 434382 704838
rect 433826 704282 434062 704518
rect 434146 704282 434382 704518
rect 462986 711322 463222 711558
rect 463306 711322 463542 711558
rect 462986 711002 463222 711238
rect 463306 711002 463542 711238
rect 459266 709402 459502 709638
rect 459586 709402 459822 709638
rect 459266 709082 459502 709318
rect 459586 709082 459822 709318
rect 455546 707482 455782 707718
rect 455866 707482 456102 707718
rect 455546 707162 455782 707398
rect 455866 707162 456102 707398
rect 451826 705562 452062 705798
rect 452146 705562 452382 705798
rect 451826 705242 452062 705478
rect 452146 705242 452382 705478
rect 480986 710362 481222 710598
rect 481306 710362 481542 710598
rect 480986 710042 481222 710278
rect 481306 710042 481542 710278
rect 477266 708442 477502 708678
rect 477586 708442 477822 708678
rect 477266 708122 477502 708358
rect 477586 708122 477822 708358
rect 473546 706522 473782 706758
rect 473866 706522 474102 706758
rect 473546 706202 473782 706438
rect 473866 706202 474102 706438
rect 469826 704602 470062 704838
rect 470146 704602 470382 704838
rect 469826 704282 470062 704518
rect 470146 704282 470382 704518
rect 498986 711322 499222 711558
rect 499306 711322 499542 711558
rect 498986 711002 499222 711238
rect 499306 711002 499542 711238
rect 495266 709402 495502 709638
rect 495586 709402 495822 709638
rect 495266 709082 495502 709318
rect 495586 709082 495822 709318
rect 491546 707482 491782 707718
rect 491866 707482 492102 707718
rect 491546 707162 491782 707398
rect 491866 707162 492102 707398
rect 487826 705562 488062 705798
rect 488146 705562 488382 705798
rect 487826 705242 488062 705478
rect 488146 705242 488382 705478
rect 516986 710362 517222 710598
rect 517306 710362 517542 710598
rect 516986 710042 517222 710278
rect 517306 710042 517542 710278
rect 513266 708442 513502 708678
rect 513586 708442 513822 708678
rect 513266 708122 513502 708358
rect 513586 708122 513822 708358
rect 509546 706522 509782 706758
rect 509866 706522 510102 706758
rect 509546 706202 509782 706438
rect 509866 706202 510102 706438
rect 505826 704602 506062 704838
rect 506146 704602 506382 704838
rect 505826 704282 506062 704518
rect 506146 704282 506382 704518
rect 534986 711322 535222 711558
rect 535306 711322 535542 711558
rect 534986 711002 535222 711238
rect 535306 711002 535542 711238
rect 531266 709402 531502 709638
rect 531586 709402 531822 709638
rect 531266 709082 531502 709318
rect 531586 709082 531822 709318
rect 527546 707482 527782 707718
rect 527866 707482 528102 707718
rect 527546 707162 527782 707398
rect 527866 707162 528102 707398
rect 523826 705562 524062 705798
rect 524146 705562 524382 705798
rect 523826 705242 524062 705478
rect 524146 705242 524382 705478
rect 552986 710362 553222 710598
rect 553306 710362 553542 710598
rect 552986 710042 553222 710278
rect 553306 710042 553542 710278
rect 549266 708442 549502 708678
rect 549586 708442 549822 708678
rect 549266 708122 549502 708358
rect 549586 708122 549822 708358
rect 545546 706522 545782 706758
rect 545866 706522 546102 706758
rect 545546 706202 545782 706438
rect 545866 706202 546102 706438
rect 541826 704602 542062 704838
rect 542146 704602 542382 704838
rect 541826 704282 542062 704518
rect 542146 704282 542382 704518
rect 570986 711322 571222 711558
rect 571306 711322 571542 711558
rect 570986 711002 571222 711238
rect 571306 711002 571542 711238
rect 567266 709402 567502 709638
rect 567586 709402 567822 709638
rect 567266 709082 567502 709318
rect 567586 709082 567822 709318
rect 563546 707482 563782 707718
rect 563866 707482 564102 707718
rect 563546 707162 563782 707398
rect 563866 707162 564102 707398
rect 559826 705562 560062 705798
rect 560146 705562 560382 705798
rect 559826 705242 560062 705478
rect 560146 705242 560382 705478
rect -1974 687218 -1738 687454
rect -1654 687218 -1418 687454
rect -1974 686898 -1738 687134
rect -1654 686898 -1418 687134
rect 8250 687218 8486 687454
rect 8250 686898 8486 687134
rect 38970 687218 39206 687454
rect 38970 686898 39206 687134
rect 69690 687218 69926 687454
rect 69690 686898 69926 687134
rect 100410 687218 100646 687454
rect 100410 686898 100646 687134
rect 131130 687218 131366 687454
rect 131130 686898 131366 687134
rect 161850 687218 162086 687454
rect 161850 686898 162086 687134
rect 192570 687218 192806 687454
rect 192570 686898 192806 687134
rect 223290 687218 223526 687454
rect 223290 686898 223526 687134
rect 254010 687218 254246 687454
rect 254010 686898 254246 687134
rect 284730 687218 284966 687454
rect 284730 686898 284966 687134
rect 315450 687218 315686 687454
rect 315450 686898 315686 687134
rect 346170 687218 346406 687454
rect 346170 686898 346406 687134
rect 376890 687218 377126 687454
rect 376890 686898 377126 687134
rect 407610 687218 407846 687454
rect 407610 686898 407846 687134
rect 438330 687218 438566 687454
rect 438330 686898 438566 687134
rect 469050 687218 469286 687454
rect 469050 686898 469286 687134
rect 499770 687218 500006 687454
rect 499770 686898 500006 687134
rect 530490 687218 530726 687454
rect 530490 686898 530726 687134
rect 561210 687218 561446 687454
rect 561210 686898 561446 687134
rect 567266 676658 567502 676894
rect 567586 676658 567822 676894
rect 567266 676338 567502 676574
rect 567586 676338 567822 676574
rect 23610 669218 23846 669454
rect 23610 668898 23846 669134
rect 54330 669218 54566 669454
rect 54330 668898 54566 669134
rect 85050 669218 85286 669454
rect 85050 668898 85286 669134
rect 115770 669218 116006 669454
rect 115770 668898 116006 669134
rect 146490 669218 146726 669454
rect 146490 668898 146726 669134
rect 177210 669218 177446 669454
rect 177210 668898 177446 669134
rect 207930 669218 208166 669454
rect 207930 668898 208166 669134
rect 238650 669218 238886 669454
rect 238650 668898 238886 669134
rect 269370 669218 269606 669454
rect 269370 668898 269606 669134
rect 300090 669218 300326 669454
rect 300090 668898 300326 669134
rect 330810 669218 331046 669454
rect 330810 668898 331046 669134
rect 361530 669218 361766 669454
rect 361530 668898 361766 669134
rect 392250 669218 392486 669454
rect 392250 668898 392486 669134
rect 422970 669218 423206 669454
rect 422970 668898 423206 669134
rect 453690 669218 453926 669454
rect 453690 668898 453926 669134
rect 484410 669218 484646 669454
rect 484410 668898 484646 669134
rect 515130 669218 515366 669454
rect 515130 668898 515366 669134
rect 545850 669218 546086 669454
rect 545850 668898 546086 669134
rect -1974 651218 -1738 651454
rect -1654 651218 -1418 651454
rect -1974 650898 -1738 651134
rect -1654 650898 -1418 651134
rect 8250 651218 8486 651454
rect 8250 650898 8486 651134
rect 38970 651218 39206 651454
rect 38970 650898 39206 651134
rect 69690 651218 69926 651454
rect 69690 650898 69926 651134
rect 100410 651218 100646 651454
rect 100410 650898 100646 651134
rect 131130 651218 131366 651454
rect 131130 650898 131366 651134
rect 161850 651218 162086 651454
rect 161850 650898 162086 651134
rect 192570 651218 192806 651454
rect 192570 650898 192806 651134
rect 223290 651218 223526 651454
rect 223290 650898 223526 651134
rect 254010 651218 254246 651454
rect 254010 650898 254246 651134
rect 284730 651218 284966 651454
rect 284730 650898 284966 651134
rect 315450 651218 315686 651454
rect 315450 650898 315686 651134
rect 346170 651218 346406 651454
rect 346170 650898 346406 651134
rect 376890 651218 377126 651454
rect 376890 650898 377126 651134
rect 407610 651218 407846 651454
rect 407610 650898 407846 651134
rect 438330 651218 438566 651454
rect 438330 650898 438566 651134
rect 469050 651218 469286 651454
rect 469050 650898 469286 651134
rect 499770 651218 500006 651454
rect 499770 650898 500006 651134
rect 530490 651218 530726 651454
rect 530490 650898 530726 651134
rect 561210 651218 561446 651454
rect 561210 650898 561446 651134
rect 567266 640658 567502 640894
rect 567586 640658 567822 640894
rect 567266 640338 567502 640574
rect 567586 640338 567822 640574
rect 23610 633218 23846 633454
rect 23610 632898 23846 633134
rect 54330 633218 54566 633454
rect 54330 632898 54566 633134
rect 85050 633218 85286 633454
rect 85050 632898 85286 633134
rect 115770 633218 116006 633454
rect 115770 632898 116006 633134
rect 146490 633218 146726 633454
rect 146490 632898 146726 633134
rect 177210 633218 177446 633454
rect 177210 632898 177446 633134
rect 207930 633218 208166 633454
rect 207930 632898 208166 633134
rect 238650 633218 238886 633454
rect 238650 632898 238886 633134
rect 269370 633218 269606 633454
rect 269370 632898 269606 633134
rect 300090 633218 300326 633454
rect 300090 632898 300326 633134
rect 330810 633218 331046 633454
rect 330810 632898 331046 633134
rect 361530 633218 361766 633454
rect 361530 632898 361766 633134
rect 392250 633218 392486 633454
rect 392250 632898 392486 633134
rect 422970 633218 423206 633454
rect 422970 632898 423206 633134
rect 453690 633218 453926 633454
rect 453690 632898 453926 633134
rect 484410 633218 484646 633454
rect 484410 632898 484646 633134
rect 515130 633218 515366 633454
rect 515130 632898 515366 633134
rect 545850 633218 546086 633454
rect 545850 632898 546086 633134
rect -1974 615218 -1738 615454
rect -1654 615218 -1418 615454
rect -1974 614898 -1738 615134
rect -1654 614898 -1418 615134
rect 8250 615218 8486 615454
rect 8250 614898 8486 615134
rect 38970 615218 39206 615454
rect 38970 614898 39206 615134
rect 69690 615218 69926 615454
rect 69690 614898 69926 615134
rect 100410 615218 100646 615454
rect 100410 614898 100646 615134
rect 131130 615218 131366 615454
rect 131130 614898 131366 615134
rect 161850 615218 162086 615454
rect 161850 614898 162086 615134
rect 192570 615218 192806 615454
rect 192570 614898 192806 615134
rect 223290 615218 223526 615454
rect 223290 614898 223526 615134
rect 254010 615218 254246 615454
rect 254010 614898 254246 615134
rect 284730 615218 284966 615454
rect 284730 614898 284966 615134
rect 315450 615218 315686 615454
rect 315450 614898 315686 615134
rect 346170 615218 346406 615454
rect 346170 614898 346406 615134
rect 376890 615218 377126 615454
rect 376890 614898 377126 615134
rect 407610 615218 407846 615454
rect 407610 614898 407846 615134
rect 438330 615218 438566 615454
rect 438330 614898 438566 615134
rect 469050 615218 469286 615454
rect 469050 614898 469286 615134
rect 499770 615218 500006 615454
rect 499770 614898 500006 615134
rect 530490 615218 530726 615454
rect 530490 614898 530726 615134
rect 561210 615218 561446 615454
rect 561210 614898 561446 615134
rect 567266 604658 567502 604894
rect 567586 604658 567822 604894
rect 567266 604338 567502 604574
rect 567586 604338 567822 604574
rect 23610 597218 23846 597454
rect 23610 596898 23846 597134
rect 54330 597218 54566 597454
rect 54330 596898 54566 597134
rect 85050 597218 85286 597454
rect 85050 596898 85286 597134
rect 115770 597218 116006 597454
rect 115770 596898 116006 597134
rect 146490 597218 146726 597454
rect 146490 596898 146726 597134
rect 177210 597218 177446 597454
rect 177210 596898 177446 597134
rect 207930 597218 208166 597454
rect 207930 596898 208166 597134
rect 238650 597218 238886 597454
rect 238650 596898 238886 597134
rect 269370 597218 269606 597454
rect 269370 596898 269606 597134
rect 300090 597218 300326 597454
rect 300090 596898 300326 597134
rect 330810 597218 331046 597454
rect 330810 596898 331046 597134
rect 361530 597218 361766 597454
rect 361530 596898 361766 597134
rect 392250 597218 392486 597454
rect 392250 596898 392486 597134
rect 422970 597218 423206 597454
rect 422970 596898 423206 597134
rect 453690 597218 453926 597454
rect 453690 596898 453926 597134
rect 484410 597218 484646 597454
rect 484410 596898 484646 597134
rect 515130 597218 515366 597454
rect 515130 596898 515366 597134
rect 545850 597218 546086 597454
rect 545850 596898 546086 597134
rect -1974 579218 -1738 579454
rect -1654 579218 -1418 579454
rect -1974 578898 -1738 579134
rect -1654 578898 -1418 579134
rect 8250 579218 8486 579454
rect 8250 578898 8486 579134
rect 38970 579218 39206 579454
rect 38970 578898 39206 579134
rect 69690 579218 69926 579454
rect 69690 578898 69926 579134
rect 100410 579218 100646 579454
rect 100410 578898 100646 579134
rect 131130 579218 131366 579454
rect 131130 578898 131366 579134
rect 161850 579218 162086 579454
rect 161850 578898 162086 579134
rect 192570 579218 192806 579454
rect 192570 578898 192806 579134
rect 223290 579218 223526 579454
rect 223290 578898 223526 579134
rect 254010 579218 254246 579454
rect 254010 578898 254246 579134
rect 284730 579218 284966 579454
rect 284730 578898 284966 579134
rect 315450 579218 315686 579454
rect 315450 578898 315686 579134
rect 346170 579218 346406 579454
rect 346170 578898 346406 579134
rect 376890 579218 377126 579454
rect 376890 578898 377126 579134
rect 407610 579218 407846 579454
rect 407610 578898 407846 579134
rect 438330 579218 438566 579454
rect 438330 578898 438566 579134
rect 469050 579218 469286 579454
rect 469050 578898 469286 579134
rect 499770 579218 500006 579454
rect 499770 578898 500006 579134
rect 530490 579218 530726 579454
rect 530490 578898 530726 579134
rect 561210 579218 561446 579454
rect 561210 578898 561446 579134
rect 567266 568658 567502 568894
rect 567586 568658 567822 568894
rect 567266 568338 567502 568574
rect 567586 568338 567822 568574
rect 23610 561218 23846 561454
rect 23610 560898 23846 561134
rect 54330 561218 54566 561454
rect 54330 560898 54566 561134
rect 85050 561218 85286 561454
rect 85050 560898 85286 561134
rect 115770 561218 116006 561454
rect 115770 560898 116006 561134
rect 146490 561218 146726 561454
rect 146490 560898 146726 561134
rect 177210 561218 177446 561454
rect 177210 560898 177446 561134
rect 207930 561218 208166 561454
rect 207930 560898 208166 561134
rect 238650 561218 238886 561454
rect 238650 560898 238886 561134
rect 269370 561218 269606 561454
rect 269370 560898 269606 561134
rect 300090 561218 300326 561454
rect 300090 560898 300326 561134
rect 330810 561218 331046 561454
rect 330810 560898 331046 561134
rect 361530 561218 361766 561454
rect 361530 560898 361766 561134
rect 392250 561218 392486 561454
rect 392250 560898 392486 561134
rect 422970 561218 423206 561454
rect 422970 560898 423206 561134
rect 453690 561218 453926 561454
rect 453690 560898 453926 561134
rect 484410 561218 484646 561454
rect 484410 560898 484646 561134
rect 515130 561218 515366 561454
rect 515130 560898 515366 561134
rect 545850 561218 546086 561454
rect 545850 560898 546086 561134
rect -1974 543218 -1738 543454
rect -1654 543218 -1418 543454
rect -1974 542898 -1738 543134
rect -1654 542898 -1418 543134
rect 8250 543218 8486 543454
rect 8250 542898 8486 543134
rect 38970 543218 39206 543454
rect 38970 542898 39206 543134
rect 69690 543218 69926 543454
rect 69690 542898 69926 543134
rect 100410 543218 100646 543454
rect 100410 542898 100646 543134
rect 131130 543218 131366 543454
rect 131130 542898 131366 543134
rect 161850 543218 162086 543454
rect 161850 542898 162086 543134
rect 192570 543218 192806 543454
rect 192570 542898 192806 543134
rect 223290 543218 223526 543454
rect 223290 542898 223526 543134
rect 254010 543218 254246 543454
rect 254010 542898 254246 543134
rect 284730 543218 284966 543454
rect 284730 542898 284966 543134
rect 315450 543218 315686 543454
rect 315450 542898 315686 543134
rect 346170 543218 346406 543454
rect 346170 542898 346406 543134
rect 376890 543218 377126 543454
rect 376890 542898 377126 543134
rect 407610 543218 407846 543454
rect 407610 542898 407846 543134
rect 438330 543218 438566 543454
rect 438330 542898 438566 543134
rect 469050 543218 469286 543454
rect 469050 542898 469286 543134
rect 499770 543218 500006 543454
rect 499770 542898 500006 543134
rect 530490 543218 530726 543454
rect 530490 542898 530726 543134
rect 561210 543218 561446 543454
rect 561210 542898 561446 543134
rect 567266 532658 567502 532894
rect 567586 532658 567822 532894
rect 567266 532338 567502 532574
rect 567586 532338 567822 532574
rect 23610 525218 23846 525454
rect 23610 524898 23846 525134
rect 54330 525218 54566 525454
rect 54330 524898 54566 525134
rect 85050 525218 85286 525454
rect 85050 524898 85286 525134
rect 115770 525218 116006 525454
rect 115770 524898 116006 525134
rect 146490 525218 146726 525454
rect 146490 524898 146726 525134
rect 177210 525218 177446 525454
rect 177210 524898 177446 525134
rect 207930 525218 208166 525454
rect 207930 524898 208166 525134
rect 238650 525218 238886 525454
rect 238650 524898 238886 525134
rect 269370 525218 269606 525454
rect 269370 524898 269606 525134
rect 300090 525218 300326 525454
rect 300090 524898 300326 525134
rect 330810 525218 331046 525454
rect 330810 524898 331046 525134
rect 361530 525218 361766 525454
rect 361530 524898 361766 525134
rect 392250 525218 392486 525454
rect 392250 524898 392486 525134
rect 422970 525218 423206 525454
rect 422970 524898 423206 525134
rect 453690 525218 453926 525454
rect 453690 524898 453926 525134
rect 484410 525218 484646 525454
rect 484410 524898 484646 525134
rect 515130 525218 515366 525454
rect 515130 524898 515366 525134
rect 545850 525218 546086 525454
rect 545850 524898 546086 525134
rect -1974 507218 -1738 507454
rect -1654 507218 -1418 507454
rect -1974 506898 -1738 507134
rect -1654 506898 -1418 507134
rect 8250 507218 8486 507454
rect 8250 506898 8486 507134
rect 38970 507218 39206 507454
rect 38970 506898 39206 507134
rect 69690 507218 69926 507454
rect 69690 506898 69926 507134
rect 100410 507218 100646 507454
rect 100410 506898 100646 507134
rect 131130 507218 131366 507454
rect 131130 506898 131366 507134
rect 161850 507218 162086 507454
rect 161850 506898 162086 507134
rect 192570 507218 192806 507454
rect 192570 506898 192806 507134
rect 223290 507218 223526 507454
rect 223290 506898 223526 507134
rect 254010 507218 254246 507454
rect 254010 506898 254246 507134
rect 284730 507218 284966 507454
rect 284730 506898 284966 507134
rect 315450 507218 315686 507454
rect 315450 506898 315686 507134
rect 346170 507218 346406 507454
rect 346170 506898 346406 507134
rect 376890 507218 377126 507454
rect 376890 506898 377126 507134
rect 407610 507218 407846 507454
rect 407610 506898 407846 507134
rect 438330 507218 438566 507454
rect 438330 506898 438566 507134
rect 469050 507218 469286 507454
rect 469050 506898 469286 507134
rect 499770 507218 500006 507454
rect 499770 506898 500006 507134
rect 530490 507218 530726 507454
rect 530490 506898 530726 507134
rect 561210 507218 561446 507454
rect 561210 506898 561446 507134
rect 567266 496658 567502 496894
rect 567586 496658 567822 496894
rect 567266 496338 567502 496574
rect 567586 496338 567822 496574
rect 23610 489218 23846 489454
rect 23610 488898 23846 489134
rect 54330 489218 54566 489454
rect 54330 488898 54566 489134
rect 85050 489218 85286 489454
rect 85050 488898 85286 489134
rect 115770 489218 116006 489454
rect 115770 488898 116006 489134
rect 146490 489218 146726 489454
rect 146490 488898 146726 489134
rect 177210 489218 177446 489454
rect 177210 488898 177446 489134
rect 207930 489218 208166 489454
rect 207930 488898 208166 489134
rect 238650 489218 238886 489454
rect 238650 488898 238886 489134
rect 269370 489218 269606 489454
rect 269370 488898 269606 489134
rect 300090 489218 300326 489454
rect 300090 488898 300326 489134
rect 330810 489218 331046 489454
rect 330810 488898 331046 489134
rect 361530 489218 361766 489454
rect 361530 488898 361766 489134
rect 392250 489218 392486 489454
rect 392250 488898 392486 489134
rect 422970 489218 423206 489454
rect 422970 488898 423206 489134
rect 453690 489218 453926 489454
rect 453690 488898 453926 489134
rect 484410 489218 484646 489454
rect 484410 488898 484646 489134
rect 515130 489218 515366 489454
rect 515130 488898 515366 489134
rect 545850 489218 546086 489454
rect 545850 488898 546086 489134
rect -1974 471218 -1738 471454
rect -1654 471218 -1418 471454
rect -1974 470898 -1738 471134
rect -1654 470898 -1418 471134
rect 8250 471218 8486 471454
rect 8250 470898 8486 471134
rect 38970 471218 39206 471454
rect 38970 470898 39206 471134
rect 69690 471218 69926 471454
rect 69690 470898 69926 471134
rect 100410 471218 100646 471454
rect 100410 470898 100646 471134
rect 131130 471218 131366 471454
rect 131130 470898 131366 471134
rect 161850 471218 162086 471454
rect 161850 470898 162086 471134
rect 192570 471218 192806 471454
rect 192570 470898 192806 471134
rect 223290 471218 223526 471454
rect 223290 470898 223526 471134
rect 254010 471218 254246 471454
rect 254010 470898 254246 471134
rect 284730 471218 284966 471454
rect 284730 470898 284966 471134
rect 315450 471218 315686 471454
rect 315450 470898 315686 471134
rect 346170 471218 346406 471454
rect 346170 470898 346406 471134
rect 376890 471218 377126 471454
rect 376890 470898 377126 471134
rect 407610 471218 407846 471454
rect 407610 470898 407846 471134
rect 438330 471218 438566 471454
rect 438330 470898 438566 471134
rect 469050 471218 469286 471454
rect 469050 470898 469286 471134
rect 499770 471218 500006 471454
rect 499770 470898 500006 471134
rect 530490 471218 530726 471454
rect 530490 470898 530726 471134
rect 561210 471218 561446 471454
rect 561210 470898 561446 471134
rect 567266 460658 567502 460894
rect 567586 460658 567822 460894
rect 567266 460338 567502 460574
rect 567586 460338 567822 460574
rect 23610 453218 23846 453454
rect 23610 452898 23846 453134
rect 54330 453218 54566 453454
rect 54330 452898 54566 453134
rect 85050 453218 85286 453454
rect 85050 452898 85286 453134
rect 115770 453218 116006 453454
rect 115770 452898 116006 453134
rect 146490 453218 146726 453454
rect 146490 452898 146726 453134
rect 177210 453218 177446 453454
rect 177210 452898 177446 453134
rect 207930 453218 208166 453454
rect 207930 452898 208166 453134
rect 238650 453218 238886 453454
rect 238650 452898 238886 453134
rect 269370 453218 269606 453454
rect 269370 452898 269606 453134
rect 300090 453218 300326 453454
rect 300090 452898 300326 453134
rect 330810 453218 331046 453454
rect 330810 452898 331046 453134
rect 361530 453218 361766 453454
rect 361530 452898 361766 453134
rect 392250 453218 392486 453454
rect 392250 452898 392486 453134
rect 422970 453218 423206 453454
rect 422970 452898 423206 453134
rect 453690 453218 453926 453454
rect 453690 452898 453926 453134
rect 484410 453218 484646 453454
rect 484410 452898 484646 453134
rect 515130 453218 515366 453454
rect 515130 452898 515366 453134
rect 545850 453218 546086 453454
rect 545850 452898 546086 453134
rect -1974 435218 -1738 435454
rect -1654 435218 -1418 435454
rect -1974 434898 -1738 435134
rect -1654 434898 -1418 435134
rect 8250 435218 8486 435454
rect 8250 434898 8486 435134
rect 38970 435218 39206 435454
rect 38970 434898 39206 435134
rect 69690 435218 69926 435454
rect 69690 434898 69926 435134
rect 100410 435218 100646 435454
rect 100410 434898 100646 435134
rect 131130 435218 131366 435454
rect 131130 434898 131366 435134
rect 161850 435218 162086 435454
rect 161850 434898 162086 435134
rect 192570 435218 192806 435454
rect 192570 434898 192806 435134
rect 223290 435218 223526 435454
rect 223290 434898 223526 435134
rect 254010 435218 254246 435454
rect 254010 434898 254246 435134
rect 284730 435218 284966 435454
rect 284730 434898 284966 435134
rect 315450 435218 315686 435454
rect 315450 434898 315686 435134
rect 346170 435218 346406 435454
rect 346170 434898 346406 435134
rect 376890 435218 377126 435454
rect 376890 434898 377126 435134
rect 407610 435218 407846 435454
rect 407610 434898 407846 435134
rect 438330 435218 438566 435454
rect 438330 434898 438566 435134
rect 469050 435218 469286 435454
rect 469050 434898 469286 435134
rect 499770 435218 500006 435454
rect 499770 434898 500006 435134
rect 530490 435218 530726 435454
rect 530490 434898 530726 435134
rect 561210 435218 561446 435454
rect 561210 434898 561446 435134
rect 567266 424658 567502 424894
rect 567586 424658 567822 424894
rect 567266 424338 567502 424574
rect 567586 424338 567822 424574
rect 23610 417218 23846 417454
rect 23610 416898 23846 417134
rect 54330 417218 54566 417454
rect 54330 416898 54566 417134
rect 85050 417218 85286 417454
rect 85050 416898 85286 417134
rect 115770 417218 116006 417454
rect 115770 416898 116006 417134
rect 146490 417218 146726 417454
rect 146490 416898 146726 417134
rect 177210 417218 177446 417454
rect 177210 416898 177446 417134
rect 207930 417218 208166 417454
rect 207930 416898 208166 417134
rect 238650 417218 238886 417454
rect 238650 416898 238886 417134
rect 269370 417218 269606 417454
rect 269370 416898 269606 417134
rect 300090 417218 300326 417454
rect 300090 416898 300326 417134
rect 330810 417218 331046 417454
rect 330810 416898 331046 417134
rect 361530 417218 361766 417454
rect 361530 416898 361766 417134
rect 392250 417218 392486 417454
rect 392250 416898 392486 417134
rect 422970 417218 423206 417454
rect 422970 416898 423206 417134
rect 453690 417218 453926 417454
rect 453690 416898 453926 417134
rect 484410 417218 484646 417454
rect 484410 416898 484646 417134
rect 515130 417218 515366 417454
rect 515130 416898 515366 417134
rect 545850 417218 546086 417454
rect 545850 416898 546086 417134
rect -1974 399218 -1738 399454
rect -1654 399218 -1418 399454
rect -1974 398898 -1738 399134
rect -1654 398898 -1418 399134
rect 8250 399218 8486 399454
rect 8250 398898 8486 399134
rect 38970 399218 39206 399454
rect 38970 398898 39206 399134
rect 69690 399218 69926 399454
rect 69690 398898 69926 399134
rect 100410 399218 100646 399454
rect 100410 398898 100646 399134
rect 131130 399218 131366 399454
rect 131130 398898 131366 399134
rect 161850 399218 162086 399454
rect 161850 398898 162086 399134
rect 192570 399218 192806 399454
rect 192570 398898 192806 399134
rect 223290 399218 223526 399454
rect 223290 398898 223526 399134
rect 254010 399218 254246 399454
rect 254010 398898 254246 399134
rect 284730 399218 284966 399454
rect 284730 398898 284966 399134
rect 315450 399218 315686 399454
rect 315450 398898 315686 399134
rect 346170 399218 346406 399454
rect 346170 398898 346406 399134
rect 376890 399218 377126 399454
rect 376890 398898 377126 399134
rect 407610 399218 407846 399454
rect 407610 398898 407846 399134
rect 438330 399218 438566 399454
rect 438330 398898 438566 399134
rect 469050 399218 469286 399454
rect 469050 398898 469286 399134
rect 499770 399218 500006 399454
rect 499770 398898 500006 399134
rect 530490 399218 530726 399454
rect 530490 398898 530726 399134
rect 561210 399218 561446 399454
rect 561210 398898 561446 399134
rect 567266 388658 567502 388894
rect 567586 388658 567822 388894
rect 567266 388338 567502 388574
rect 567586 388338 567822 388574
rect 23610 381218 23846 381454
rect 23610 380898 23846 381134
rect 54330 381218 54566 381454
rect 54330 380898 54566 381134
rect 85050 381218 85286 381454
rect 85050 380898 85286 381134
rect 115770 381218 116006 381454
rect 115770 380898 116006 381134
rect 146490 381218 146726 381454
rect 146490 380898 146726 381134
rect 177210 381218 177446 381454
rect 177210 380898 177446 381134
rect 207930 381218 208166 381454
rect 207930 380898 208166 381134
rect 238650 381218 238886 381454
rect 238650 380898 238886 381134
rect 269370 381218 269606 381454
rect 269370 380898 269606 381134
rect 300090 381218 300326 381454
rect 300090 380898 300326 381134
rect 330810 381218 331046 381454
rect 330810 380898 331046 381134
rect 361530 381218 361766 381454
rect 361530 380898 361766 381134
rect 392250 381218 392486 381454
rect 392250 380898 392486 381134
rect 422970 381218 423206 381454
rect 422970 380898 423206 381134
rect 453690 381218 453926 381454
rect 453690 380898 453926 381134
rect 484410 381218 484646 381454
rect 484410 380898 484646 381134
rect 515130 381218 515366 381454
rect 515130 380898 515366 381134
rect 545850 381218 546086 381454
rect 545850 380898 546086 381134
rect -1974 363218 -1738 363454
rect -1654 363218 -1418 363454
rect -1974 362898 -1738 363134
rect -1654 362898 -1418 363134
rect 8250 363218 8486 363454
rect 8250 362898 8486 363134
rect 38970 363218 39206 363454
rect 38970 362898 39206 363134
rect 69690 363218 69926 363454
rect 69690 362898 69926 363134
rect 100410 363218 100646 363454
rect 100410 362898 100646 363134
rect 131130 363218 131366 363454
rect 131130 362898 131366 363134
rect 161850 363218 162086 363454
rect 161850 362898 162086 363134
rect 192570 363218 192806 363454
rect 192570 362898 192806 363134
rect 223290 363218 223526 363454
rect 223290 362898 223526 363134
rect 254010 363218 254246 363454
rect 254010 362898 254246 363134
rect 284730 363218 284966 363454
rect 284730 362898 284966 363134
rect 315450 363218 315686 363454
rect 315450 362898 315686 363134
rect 346170 363218 346406 363454
rect 346170 362898 346406 363134
rect 376890 363218 377126 363454
rect 376890 362898 377126 363134
rect 407610 363218 407846 363454
rect 407610 362898 407846 363134
rect 438330 363218 438566 363454
rect 438330 362898 438566 363134
rect 469050 363218 469286 363454
rect 469050 362898 469286 363134
rect 499770 363218 500006 363454
rect 499770 362898 500006 363134
rect 530490 363218 530726 363454
rect 530490 362898 530726 363134
rect 561210 363218 561446 363454
rect 561210 362898 561446 363134
rect 567266 352658 567502 352894
rect 567586 352658 567822 352894
rect 567266 352338 567502 352574
rect 567586 352338 567822 352574
rect 23610 345218 23846 345454
rect 23610 344898 23846 345134
rect 54330 345218 54566 345454
rect 54330 344898 54566 345134
rect 85050 345218 85286 345454
rect 85050 344898 85286 345134
rect 115770 345218 116006 345454
rect 115770 344898 116006 345134
rect 146490 345218 146726 345454
rect 146490 344898 146726 345134
rect 177210 345218 177446 345454
rect 177210 344898 177446 345134
rect 207930 345218 208166 345454
rect 207930 344898 208166 345134
rect 238650 345218 238886 345454
rect 238650 344898 238886 345134
rect 269370 345218 269606 345454
rect 269370 344898 269606 345134
rect 300090 345218 300326 345454
rect 300090 344898 300326 345134
rect 330810 345218 331046 345454
rect 330810 344898 331046 345134
rect 361530 345218 361766 345454
rect 361530 344898 361766 345134
rect 392250 345218 392486 345454
rect 392250 344898 392486 345134
rect 422970 345218 423206 345454
rect 422970 344898 423206 345134
rect 453690 345218 453926 345454
rect 453690 344898 453926 345134
rect 484410 345218 484646 345454
rect 484410 344898 484646 345134
rect 515130 345218 515366 345454
rect 515130 344898 515366 345134
rect 545850 345218 546086 345454
rect 545850 344898 546086 345134
rect -1974 327218 -1738 327454
rect -1654 327218 -1418 327454
rect -1974 326898 -1738 327134
rect -1654 326898 -1418 327134
rect 8250 327218 8486 327454
rect 8250 326898 8486 327134
rect 38970 327218 39206 327454
rect 38970 326898 39206 327134
rect 69690 327218 69926 327454
rect 69690 326898 69926 327134
rect 100410 327218 100646 327454
rect 100410 326898 100646 327134
rect 131130 327218 131366 327454
rect 131130 326898 131366 327134
rect 161850 327218 162086 327454
rect 161850 326898 162086 327134
rect 192570 327218 192806 327454
rect 192570 326898 192806 327134
rect 223290 327218 223526 327454
rect 223290 326898 223526 327134
rect 254010 327218 254246 327454
rect 254010 326898 254246 327134
rect 284730 327218 284966 327454
rect 284730 326898 284966 327134
rect 315450 327218 315686 327454
rect 315450 326898 315686 327134
rect 346170 327218 346406 327454
rect 346170 326898 346406 327134
rect 376890 327218 377126 327454
rect 376890 326898 377126 327134
rect 407610 327218 407846 327454
rect 407610 326898 407846 327134
rect 438330 327218 438566 327454
rect 438330 326898 438566 327134
rect 469050 327218 469286 327454
rect 469050 326898 469286 327134
rect 499770 327218 500006 327454
rect 499770 326898 500006 327134
rect 530490 327218 530726 327454
rect 530490 326898 530726 327134
rect 561210 327218 561446 327454
rect 561210 326898 561446 327134
rect 567266 316658 567502 316894
rect 567586 316658 567822 316894
rect 567266 316338 567502 316574
rect 567586 316338 567822 316574
rect 23610 309218 23846 309454
rect 23610 308898 23846 309134
rect 54330 309218 54566 309454
rect 54330 308898 54566 309134
rect 85050 309218 85286 309454
rect 85050 308898 85286 309134
rect 115770 309218 116006 309454
rect 115770 308898 116006 309134
rect 146490 309218 146726 309454
rect 146490 308898 146726 309134
rect 177210 309218 177446 309454
rect 177210 308898 177446 309134
rect 207930 309218 208166 309454
rect 207930 308898 208166 309134
rect 238650 309218 238886 309454
rect 238650 308898 238886 309134
rect 269370 309218 269606 309454
rect 269370 308898 269606 309134
rect 300090 309218 300326 309454
rect 300090 308898 300326 309134
rect 330810 309218 331046 309454
rect 330810 308898 331046 309134
rect 361530 309218 361766 309454
rect 361530 308898 361766 309134
rect 392250 309218 392486 309454
rect 392250 308898 392486 309134
rect 422970 309218 423206 309454
rect 422970 308898 423206 309134
rect 453690 309218 453926 309454
rect 453690 308898 453926 309134
rect 484410 309218 484646 309454
rect 484410 308898 484646 309134
rect 515130 309218 515366 309454
rect 515130 308898 515366 309134
rect 545850 309218 546086 309454
rect 545850 308898 546086 309134
rect -1974 291218 -1738 291454
rect -1654 291218 -1418 291454
rect -1974 290898 -1738 291134
rect -1654 290898 -1418 291134
rect 8250 291218 8486 291454
rect 8250 290898 8486 291134
rect 38970 291218 39206 291454
rect 38970 290898 39206 291134
rect 69690 291218 69926 291454
rect 69690 290898 69926 291134
rect 100410 291218 100646 291454
rect 100410 290898 100646 291134
rect 131130 291218 131366 291454
rect 131130 290898 131366 291134
rect 161850 291218 162086 291454
rect 161850 290898 162086 291134
rect 192570 291218 192806 291454
rect 192570 290898 192806 291134
rect 223290 291218 223526 291454
rect 223290 290898 223526 291134
rect 254010 291218 254246 291454
rect 254010 290898 254246 291134
rect 284730 291218 284966 291454
rect 284730 290898 284966 291134
rect 315450 291218 315686 291454
rect 315450 290898 315686 291134
rect 346170 291218 346406 291454
rect 346170 290898 346406 291134
rect 376890 291218 377126 291454
rect 376890 290898 377126 291134
rect 407610 291218 407846 291454
rect 407610 290898 407846 291134
rect 438330 291218 438566 291454
rect 438330 290898 438566 291134
rect 469050 291218 469286 291454
rect 469050 290898 469286 291134
rect 499770 291218 500006 291454
rect 499770 290898 500006 291134
rect 530490 291218 530726 291454
rect 530490 290898 530726 291134
rect 561210 291218 561446 291454
rect 561210 290898 561446 291134
rect 567266 280658 567502 280894
rect 567586 280658 567822 280894
rect 567266 280338 567502 280574
rect 567586 280338 567822 280574
rect 23610 273218 23846 273454
rect 23610 272898 23846 273134
rect 54330 273218 54566 273454
rect 54330 272898 54566 273134
rect 85050 273218 85286 273454
rect 85050 272898 85286 273134
rect 115770 273218 116006 273454
rect 115770 272898 116006 273134
rect 146490 273218 146726 273454
rect 146490 272898 146726 273134
rect 177210 273218 177446 273454
rect 177210 272898 177446 273134
rect 207930 273218 208166 273454
rect 207930 272898 208166 273134
rect 238650 273218 238886 273454
rect 238650 272898 238886 273134
rect 269370 273218 269606 273454
rect 269370 272898 269606 273134
rect 300090 273218 300326 273454
rect 300090 272898 300326 273134
rect 330810 273218 331046 273454
rect 330810 272898 331046 273134
rect 361530 273218 361766 273454
rect 361530 272898 361766 273134
rect 392250 273218 392486 273454
rect 392250 272898 392486 273134
rect 422970 273218 423206 273454
rect 422970 272898 423206 273134
rect 453690 273218 453926 273454
rect 453690 272898 453926 273134
rect 484410 273218 484646 273454
rect 484410 272898 484646 273134
rect 515130 273218 515366 273454
rect 515130 272898 515366 273134
rect 545850 273218 546086 273454
rect 545850 272898 546086 273134
rect -1974 255218 -1738 255454
rect -1654 255218 -1418 255454
rect -1974 254898 -1738 255134
rect -1654 254898 -1418 255134
rect 8250 255218 8486 255454
rect 8250 254898 8486 255134
rect 38970 255218 39206 255454
rect 38970 254898 39206 255134
rect 69690 255218 69926 255454
rect 69690 254898 69926 255134
rect 100410 255218 100646 255454
rect 100410 254898 100646 255134
rect 131130 255218 131366 255454
rect 131130 254898 131366 255134
rect 161850 255218 162086 255454
rect 161850 254898 162086 255134
rect 192570 255218 192806 255454
rect 192570 254898 192806 255134
rect 223290 255218 223526 255454
rect 223290 254898 223526 255134
rect 254010 255218 254246 255454
rect 254010 254898 254246 255134
rect 284730 255218 284966 255454
rect 284730 254898 284966 255134
rect 315450 255218 315686 255454
rect 315450 254898 315686 255134
rect 346170 255218 346406 255454
rect 346170 254898 346406 255134
rect 376890 255218 377126 255454
rect 376890 254898 377126 255134
rect 407610 255218 407846 255454
rect 407610 254898 407846 255134
rect 438330 255218 438566 255454
rect 438330 254898 438566 255134
rect 469050 255218 469286 255454
rect 469050 254898 469286 255134
rect 499770 255218 500006 255454
rect 499770 254898 500006 255134
rect 530490 255218 530726 255454
rect 530490 254898 530726 255134
rect 561210 255218 561446 255454
rect 561210 254898 561446 255134
rect 567266 244658 567502 244894
rect 567586 244658 567822 244894
rect 567266 244338 567502 244574
rect 567586 244338 567822 244574
rect 23610 237218 23846 237454
rect 23610 236898 23846 237134
rect 54330 237218 54566 237454
rect 54330 236898 54566 237134
rect 85050 237218 85286 237454
rect 85050 236898 85286 237134
rect 115770 237218 116006 237454
rect 115770 236898 116006 237134
rect 146490 237218 146726 237454
rect 146490 236898 146726 237134
rect 177210 237218 177446 237454
rect 177210 236898 177446 237134
rect 207930 237218 208166 237454
rect 207930 236898 208166 237134
rect 238650 237218 238886 237454
rect 238650 236898 238886 237134
rect 269370 237218 269606 237454
rect 269370 236898 269606 237134
rect 300090 237218 300326 237454
rect 300090 236898 300326 237134
rect 330810 237218 331046 237454
rect 330810 236898 331046 237134
rect 361530 237218 361766 237454
rect 361530 236898 361766 237134
rect 392250 237218 392486 237454
rect 392250 236898 392486 237134
rect 422970 237218 423206 237454
rect 422970 236898 423206 237134
rect 453690 237218 453926 237454
rect 453690 236898 453926 237134
rect 484410 237218 484646 237454
rect 484410 236898 484646 237134
rect 515130 237218 515366 237454
rect 515130 236898 515366 237134
rect 545850 237218 546086 237454
rect 545850 236898 546086 237134
rect -1974 219218 -1738 219454
rect -1654 219218 -1418 219454
rect -1974 218898 -1738 219134
rect -1654 218898 -1418 219134
rect 8250 219218 8486 219454
rect 8250 218898 8486 219134
rect 38970 219218 39206 219454
rect 38970 218898 39206 219134
rect 69690 219218 69926 219454
rect 69690 218898 69926 219134
rect 100410 219218 100646 219454
rect 100410 218898 100646 219134
rect 131130 219218 131366 219454
rect 131130 218898 131366 219134
rect 161850 219218 162086 219454
rect 161850 218898 162086 219134
rect 192570 219218 192806 219454
rect 192570 218898 192806 219134
rect 223290 219218 223526 219454
rect 223290 218898 223526 219134
rect 254010 219218 254246 219454
rect 254010 218898 254246 219134
rect 284730 219218 284966 219454
rect 284730 218898 284966 219134
rect 315450 219218 315686 219454
rect 315450 218898 315686 219134
rect 346170 219218 346406 219454
rect 346170 218898 346406 219134
rect 376890 219218 377126 219454
rect 376890 218898 377126 219134
rect 407610 219218 407846 219454
rect 407610 218898 407846 219134
rect 438330 219218 438566 219454
rect 438330 218898 438566 219134
rect 469050 219218 469286 219454
rect 469050 218898 469286 219134
rect 499770 219218 500006 219454
rect 499770 218898 500006 219134
rect 530490 219218 530726 219454
rect 530490 218898 530726 219134
rect 561210 219218 561446 219454
rect 561210 218898 561446 219134
rect 567266 208658 567502 208894
rect 567586 208658 567822 208894
rect 567266 208338 567502 208574
rect 567586 208338 567822 208574
rect 23610 201218 23846 201454
rect 23610 200898 23846 201134
rect 54330 201218 54566 201454
rect 54330 200898 54566 201134
rect 85050 201218 85286 201454
rect 85050 200898 85286 201134
rect 115770 201218 116006 201454
rect 115770 200898 116006 201134
rect 146490 201218 146726 201454
rect 146490 200898 146726 201134
rect 177210 201218 177446 201454
rect 177210 200898 177446 201134
rect 207930 201218 208166 201454
rect 207930 200898 208166 201134
rect 238650 201218 238886 201454
rect 238650 200898 238886 201134
rect 269370 201218 269606 201454
rect 269370 200898 269606 201134
rect 300090 201218 300326 201454
rect 300090 200898 300326 201134
rect 330810 201218 331046 201454
rect 330810 200898 331046 201134
rect 361530 201218 361766 201454
rect 361530 200898 361766 201134
rect 392250 201218 392486 201454
rect 392250 200898 392486 201134
rect 422970 201218 423206 201454
rect 422970 200898 423206 201134
rect 453690 201218 453926 201454
rect 453690 200898 453926 201134
rect 484410 201218 484646 201454
rect 484410 200898 484646 201134
rect 515130 201218 515366 201454
rect 515130 200898 515366 201134
rect 545850 201218 546086 201454
rect 545850 200898 546086 201134
rect -1974 183218 -1738 183454
rect -1654 183218 -1418 183454
rect -1974 182898 -1738 183134
rect -1654 182898 -1418 183134
rect 8250 183218 8486 183454
rect 8250 182898 8486 183134
rect 38970 183218 39206 183454
rect 38970 182898 39206 183134
rect 69690 183218 69926 183454
rect 69690 182898 69926 183134
rect 100410 183218 100646 183454
rect 100410 182898 100646 183134
rect 131130 183218 131366 183454
rect 131130 182898 131366 183134
rect 161850 183218 162086 183454
rect 161850 182898 162086 183134
rect 192570 183218 192806 183454
rect 192570 182898 192806 183134
rect 223290 183218 223526 183454
rect 223290 182898 223526 183134
rect 254010 183218 254246 183454
rect 254010 182898 254246 183134
rect 284730 183218 284966 183454
rect 284730 182898 284966 183134
rect 315450 183218 315686 183454
rect 315450 182898 315686 183134
rect 346170 183218 346406 183454
rect 346170 182898 346406 183134
rect 376890 183218 377126 183454
rect 376890 182898 377126 183134
rect 407610 183218 407846 183454
rect 407610 182898 407846 183134
rect 438330 183218 438566 183454
rect 438330 182898 438566 183134
rect 469050 183218 469286 183454
rect 469050 182898 469286 183134
rect 499770 183218 500006 183454
rect 499770 182898 500006 183134
rect 530490 183218 530726 183454
rect 530490 182898 530726 183134
rect 561210 183218 561446 183454
rect 561210 182898 561446 183134
rect 567266 172658 567502 172894
rect 567586 172658 567822 172894
rect 567266 172338 567502 172574
rect 567586 172338 567822 172574
rect 23610 165218 23846 165454
rect 23610 164898 23846 165134
rect 54330 165218 54566 165454
rect 54330 164898 54566 165134
rect 85050 165218 85286 165454
rect 85050 164898 85286 165134
rect 115770 165218 116006 165454
rect 115770 164898 116006 165134
rect 146490 165218 146726 165454
rect 146490 164898 146726 165134
rect 177210 165218 177446 165454
rect 177210 164898 177446 165134
rect 207930 165218 208166 165454
rect 207930 164898 208166 165134
rect 238650 165218 238886 165454
rect 238650 164898 238886 165134
rect 269370 165218 269606 165454
rect 269370 164898 269606 165134
rect 300090 165218 300326 165454
rect 300090 164898 300326 165134
rect 330810 165218 331046 165454
rect 330810 164898 331046 165134
rect 361530 165218 361766 165454
rect 361530 164898 361766 165134
rect 392250 165218 392486 165454
rect 392250 164898 392486 165134
rect 422970 165218 423206 165454
rect 422970 164898 423206 165134
rect 453690 165218 453926 165454
rect 453690 164898 453926 165134
rect 484410 165218 484646 165454
rect 484410 164898 484646 165134
rect 515130 165218 515366 165454
rect 515130 164898 515366 165134
rect 545850 165218 546086 165454
rect 545850 164898 546086 165134
rect -1974 147218 -1738 147454
rect -1654 147218 -1418 147454
rect -1974 146898 -1738 147134
rect -1654 146898 -1418 147134
rect 8250 147218 8486 147454
rect 8250 146898 8486 147134
rect 38970 147218 39206 147454
rect 38970 146898 39206 147134
rect 69690 147218 69926 147454
rect 69690 146898 69926 147134
rect 100410 147218 100646 147454
rect 100410 146898 100646 147134
rect 131130 147218 131366 147454
rect 131130 146898 131366 147134
rect 161850 147218 162086 147454
rect 161850 146898 162086 147134
rect 192570 147218 192806 147454
rect 192570 146898 192806 147134
rect 223290 147218 223526 147454
rect 223290 146898 223526 147134
rect 254010 147218 254246 147454
rect 254010 146898 254246 147134
rect 284730 147218 284966 147454
rect 284730 146898 284966 147134
rect 315450 147218 315686 147454
rect 315450 146898 315686 147134
rect 346170 147218 346406 147454
rect 346170 146898 346406 147134
rect 376890 147218 377126 147454
rect 376890 146898 377126 147134
rect 407610 147218 407846 147454
rect 407610 146898 407846 147134
rect 438330 147218 438566 147454
rect 438330 146898 438566 147134
rect 469050 147218 469286 147454
rect 469050 146898 469286 147134
rect 499770 147218 500006 147454
rect 499770 146898 500006 147134
rect 530490 147218 530726 147454
rect 530490 146898 530726 147134
rect 561210 147218 561446 147454
rect 561210 146898 561446 147134
rect 567266 136658 567502 136894
rect 567586 136658 567822 136894
rect 567266 136338 567502 136574
rect 567586 136338 567822 136574
rect 23610 129218 23846 129454
rect 23610 128898 23846 129134
rect 54330 129218 54566 129454
rect 54330 128898 54566 129134
rect 85050 129218 85286 129454
rect 85050 128898 85286 129134
rect 115770 129218 116006 129454
rect 115770 128898 116006 129134
rect 146490 129218 146726 129454
rect 146490 128898 146726 129134
rect 177210 129218 177446 129454
rect 177210 128898 177446 129134
rect 207930 129218 208166 129454
rect 207930 128898 208166 129134
rect 238650 129218 238886 129454
rect 238650 128898 238886 129134
rect 269370 129218 269606 129454
rect 269370 128898 269606 129134
rect 300090 129218 300326 129454
rect 300090 128898 300326 129134
rect 330810 129218 331046 129454
rect 330810 128898 331046 129134
rect 361530 129218 361766 129454
rect 361530 128898 361766 129134
rect 392250 129218 392486 129454
rect 392250 128898 392486 129134
rect 422970 129218 423206 129454
rect 422970 128898 423206 129134
rect 453690 129218 453926 129454
rect 453690 128898 453926 129134
rect 484410 129218 484646 129454
rect 484410 128898 484646 129134
rect 515130 129218 515366 129454
rect 515130 128898 515366 129134
rect 545850 129218 546086 129454
rect 545850 128898 546086 129134
rect -1974 111218 -1738 111454
rect -1654 111218 -1418 111454
rect -1974 110898 -1738 111134
rect -1654 110898 -1418 111134
rect 8250 111218 8486 111454
rect 8250 110898 8486 111134
rect 38970 111218 39206 111454
rect 38970 110898 39206 111134
rect 69690 111218 69926 111454
rect 69690 110898 69926 111134
rect 100410 111218 100646 111454
rect 100410 110898 100646 111134
rect 131130 111218 131366 111454
rect 131130 110898 131366 111134
rect 161850 111218 162086 111454
rect 161850 110898 162086 111134
rect 192570 111218 192806 111454
rect 192570 110898 192806 111134
rect 223290 111218 223526 111454
rect 223290 110898 223526 111134
rect 254010 111218 254246 111454
rect 254010 110898 254246 111134
rect 284730 111218 284966 111454
rect 284730 110898 284966 111134
rect 315450 111218 315686 111454
rect 315450 110898 315686 111134
rect 346170 111218 346406 111454
rect 346170 110898 346406 111134
rect 376890 111218 377126 111454
rect 376890 110898 377126 111134
rect 407610 111218 407846 111454
rect 407610 110898 407846 111134
rect 438330 111218 438566 111454
rect 438330 110898 438566 111134
rect 469050 111218 469286 111454
rect 469050 110898 469286 111134
rect 499770 111218 500006 111454
rect 499770 110898 500006 111134
rect 530490 111218 530726 111454
rect 530490 110898 530726 111134
rect 561210 111218 561446 111454
rect 561210 110898 561446 111134
rect 567266 100658 567502 100894
rect 567586 100658 567822 100894
rect 567266 100338 567502 100574
rect 567586 100338 567822 100574
rect 23610 93218 23846 93454
rect 23610 92898 23846 93134
rect 54330 93218 54566 93454
rect 54330 92898 54566 93134
rect 85050 93218 85286 93454
rect 85050 92898 85286 93134
rect 115770 93218 116006 93454
rect 115770 92898 116006 93134
rect 146490 93218 146726 93454
rect 146490 92898 146726 93134
rect 177210 93218 177446 93454
rect 177210 92898 177446 93134
rect 207930 93218 208166 93454
rect 207930 92898 208166 93134
rect 238650 93218 238886 93454
rect 238650 92898 238886 93134
rect 269370 93218 269606 93454
rect 269370 92898 269606 93134
rect 300090 93218 300326 93454
rect 300090 92898 300326 93134
rect 330810 93218 331046 93454
rect 330810 92898 331046 93134
rect 361530 93218 361766 93454
rect 361530 92898 361766 93134
rect 392250 93218 392486 93454
rect 392250 92898 392486 93134
rect 422970 93218 423206 93454
rect 422970 92898 423206 93134
rect 453690 93218 453926 93454
rect 453690 92898 453926 93134
rect 484410 93218 484646 93454
rect 484410 92898 484646 93134
rect 515130 93218 515366 93454
rect 515130 92898 515366 93134
rect 545850 93218 546086 93454
rect 545850 92898 546086 93134
rect -1974 75218 -1738 75454
rect -1654 75218 -1418 75454
rect -1974 74898 -1738 75134
rect -1654 74898 -1418 75134
rect 8250 75218 8486 75454
rect 8250 74898 8486 75134
rect 38970 75218 39206 75454
rect 38970 74898 39206 75134
rect 69690 75218 69926 75454
rect 69690 74898 69926 75134
rect 100410 75218 100646 75454
rect 100410 74898 100646 75134
rect 131130 75218 131366 75454
rect 131130 74898 131366 75134
rect 161850 75218 162086 75454
rect 161850 74898 162086 75134
rect 192570 75218 192806 75454
rect 192570 74898 192806 75134
rect 223290 75218 223526 75454
rect 223290 74898 223526 75134
rect 254010 75218 254246 75454
rect 254010 74898 254246 75134
rect 284730 75218 284966 75454
rect 284730 74898 284966 75134
rect 315450 75218 315686 75454
rect 315450 74898 315686 75134
rect 346170 75218 346406 75454
rect 346170 74898 346406 75134
rect 376890 75218 377126 75454
rect 376890 74898 377126 75134
rect 407610 75218 407846 75454
rect 407610 74898 407846 75134
rect 438330 75218 438566 75454
rect 438330 74898 438566 75134
rect 469050 75218 469286 75454
rect 469050 74898 469286 75134
rect 499770 75218 500006 75454
rect 499770 74898 500006 75134
rect 530490 75218 530726 75454
rect 530490 74898 530726 75134
rect 561210 75218 561446 75454
rect 561210 74898 561446 75134
rect 567266 64658 567502 64894
rect 567586 64658 567822 64894
rect 567266 64338 567502 64574
rect 567586 64338 567822 64574
rect 23610 57218 23846 57454
rect 23610 56898 23846 57134
rect 54330 57218 54566 57454
rect 54330 56898 54566 57134
rect 85050 57218 85286 57454
rect 85050 56898 85286 57134
rect 115770 57218 116006 57454
rect 115770 56898 116006 57134
rect 146490 57218 146726 57454
rect 146490 56898 146726 57134
rect 177210 57218 177446 57454
rect 177210 56898 177446 57134
rect 207930 57218 208166 57454
rect 207930 56898 208166 57134
rect 238650 57218 238886 57454
rect 238650 56898 238886 57134
rect 269370 57218 269606 57454
rect 269370 56898 269606 57134
rect 300090 57218 300326 57454
rect 300090 56898 300326 57134
rect 330810 57218 331046 57454
rect 330810 56898 331046 57134
rect 361530 57218 361766 57454
rect 361530 56898 361766 57134
rect 392250 57218 392486 57454
rect 392250 56898 392486 57134
rect 422970 57218 423206 57454
rect 422970 56898 423206 57134
rect 453690 57218 453926 57454
rect 453690 56898 453926 57134
rect 484410 57218 484646 57454
rect 484410 56898 484646 57134
rect 515130 57218 515366 57454
rect 515130 56898 515366 57134
rect 545850 57218 546086 57454
rect 545850 56898 546086 57134
rect -1974 39218 -1738 39454
rect -1654 39218 -1418 39454
rect -1974 38898 -1738 39134
rect -1654 38898 -1418 39134
rect 8250 39218 8486 39454
rect 8250 38898 8486 39134
rect 38970 39218 39206 39454
rect 38970 38898 39206 39134
rect 69690 39218 69926 39454
rect 69690 38898 69926 39134
rect 100410 39218 100646 39454
rect 100410 38898 100646 39134
rect 131130 39218 131366 39454
rect 131130 38898 131366 39134
rect 161850 39218 162086 39454
rect 161850 38898 162086 39134
rect 192570 39218 192806 39454
rect 192570 38898 192806 39134
rect 223290 39218 223526 39454
rect 223290 38898 223526 39134
rect 254010 39218 254246 39454
rect 254010 38898 254246 39134
rect 284730 39218 284966 39454
rect 284730 38898 284966 39134
rect 315450 39218 315686 39454
rect 315450 38898 315686 39134
rect 346170 39218 346406 39454
rect 346170 38898 346406 39134
rect 376890 39218 377126 39454
rect 376890 38898 377126 39134
rect 407610 39218 407846 39454
rect 407610 38898 407846 39134
rect 438330 39218 438566 39454
rect 438330 38898 438566 39134
rect 469050 39218 469286 39454
rect 469050 38898 469286 39134
rect 499770 39218 500006 39454
rect 499770 38898 500006 39134
rect 530490 39218 530726 39454
rect 530490 38898 530726 39134
rect 561210 39218 561446 39454
rect 561210 38898 561446 39134
rect 567266 28658 567502 28894
rect 567586 28658 567822 28894
rect 567266 28338 567502 28574
rect 567586 28338 567822 28574
rect 23610 21218 23846 21454
rect 23610 20898 23846 21134
rect 54330 21218 54566 21454
rect 54330 20898 54566 21134
rect 85050 21218 85286 21454
rect 85050 20898 85286 21134
rect 115770 21218 116006 21454
rect 115770 20898 116006 21134
rect 146490 21218 146726 21454
rect 146490 20898 146726 21134
rect 177210 21218 177446 21454
rect 177210 20898 177446 21134
rect 207930 21218 208166 21454
rect 207930 20898 208166 21134
rect 238650 21218 238886 21454
rect 238650 20898 238886 21134
rect 269370 21218 269606 21454
rect 269370 20898 269606 21134
rect 300090 21218 300326 21454
rect 300090 20898 300326 21134
rect 330810 21218 331046 21454
rect 330810 20898 331046 21134
rect 361530 21218 361766 21454
rect 361530 20898 361766 21134
rect 392250 21218 392486 21454
rect 392250 20898 392486 21134
rect 422970 21218 423206 21454
rect 422970 20898 423206 21134
rect 453690 21218 453926 21454
rect 453690 20898 453926 21134
rect 484410 21218 484646 21454
rect 484410 20898 484646 21134
rect 515130 21218 515366 21454
rect 515130 20898 515366 21134
rect 545850 21218 546086 21454
rect 545850 20898 546086 21134
rect -1974 3218 -1738 3454
rect -1654 3218 -1418 3454
rect -1974 2898 -1738 3134
rect -1654 2898 -1418 3134
rect 8250 3218 8486 3454
rect 8250 2898 8486 3134
rect 38970 3218 39206 3454
rect 38970 2898 39206 3134
rect 69690 3218 69926 3454
rect 69690 2898 69926 3134
rect 100410 3218 100646 3454
rect 100410 2898 100646 3134
rect 131130 3218 131366 3454
rect 131130 2898 131366 3134
rect 161850 3218 162086 3454
rect 161850 2898 162086 3134
rect 192570 3218 192806 3454
rect 192570 2898 192806 3134
rect 223290 3218 223526 3454
rect 223290 2898 223526 3134
rect 254010 3218 254246 3454
rect 254010 2898 254246 3134
rect 284730 3218 284966 3454
rect 284730 2898 284966 3134
rect 315450 3218 315686 3454
rect 315450 2898 315686 3134
rect 346170 3218 346406 3454
rect 346170 2898 346406 3134
rect 376890 3218 377126 3454
rect 376890 2898 377126 3134
rect 407610 3218 407846 3454
rect 407610 2898 407846 3134
rect 438330 3218 438566 3454
rect 438330 2898 438566 3134
rect 469050 3218 469286 3454
rect 469050 2898 469286 3134
rect 499770 3218 500006 3454
rect 499770 2898 500006 3134
rect 530490 3218 530726 3454
rect 530490 2898 530726 3134
rect 561210 3218 561446 3454
rect 561210 2898 561446 3134
rect -1974 -582 -1738 -346
rect -1654 -582 -1418 -346
rect -1974 -902 -1738 -666
rect -1654 -902 -1418 -666
rect -2934 -1542 -2698 -1306
rect -2614 -1542 -2378 -1306
rect -2934 -1862 -2698 -1626
rect -2614 -1862 -2378 -1626
rect -3894 -2502 -3658 -2266
rect -3574 -2502 -3338 -2266
rect -3894 -2822 -3658 -2586
rect -3574 -2822 -3338 -2586
rect 5546 -2502 5782 -2266
rect 5866 -2502 6102 -2266
rect 5546 -2822 5782 -2586
rect 5866 -2822 6102 -2586
rect -4854 -3462 -4618 -3226
rect -4534 -3462 -4298 -3226
rect -4854 -3782 -4618 -3546
rect -4534 -3782 -4298 -3546
rect -5814 -4422 -5578 -4186
rect -5494 -4422 -5258 -4186
rect -5814 -4742 -5578 -4506
rect -5494 -4742 -5258 -4506
rect 9266 -4422 9502 -4186
rect 9586 -4422 9822 -4186
rect 9266 -4742 9502 -4506
rect 9586 -4742 9822 -4506
rect -6774 -5382 -6538 -5146
rect -6454 -5382 -6218 -5146
rect -6774 -5702 -6538 -5466
rect -6454 -5702 -6218 -5466
rect -7734 -6342 -7498 -6106
rect -7414 -6342 -7178 -6106
rect -7734 -6662 -7498 -6426
rect -7414 -6662 -7178 -6426
rect 23546 -3462 23782 -3226
rect 23866 -3462 24102 -3226
rect 23546 -3782 23782 -3546
rect 23866 -3782 24102 -3546
rect 27266 -5382 27502 -5146
rect 27586 -5382 27822 -5146
rect 27266 -5702 27502 -5466
rect 27586 -5702 27822 -5466
rect 12986 -6342 13222 -6106
rect 13306 -6342 13542 -6106
rect 12986 -6662 13222 -6426
rect 13306 -6662 13542 -6426
rect -8694 -7302 -8458 -7066
rect -8374 -7302 -8138 -7066
rect -8694 -7622 -8458 -7386
rect -8374 -7622 -8138 -7386
rect 41546 -2502 41782 -2266
rect 41866 -2502 42102 -2266
rect 41546 -2822 41782 -2586
rect 41866 -2822 42102 -2586
rect 45266 -4422 45502 -4186
rect 45586 -4422 45822 -4186
rect 45266 -4742 45502 -4506
rect 45586 -4742 45822 -4506
rect 30986 -7302 31222 -7066
rect 31306 -7302 31542 -7066
rect 30986 -7622 31222 -7386
rect 31306 -7622 31542 -7386
rect 59546 -3462 59782 -3226
rect 59866 -3462 60102 -3226
rect 59546 -3782 59782 -3546
rect 59866 -3782 60102 -3546
rect 63266 -5382 63502 -5146
rect 63586 -5382 63822 -5146
rect 63266 -5702 63502 -5466
rect 63586 -5702 63822 -5466
rect 48986 -6342 49222 -6106
rect 49306 -6342 49542 -6106
rect 48986 -6662 49222 -6426
rect 49306 -6662 49542 -6426
rect 77546 -2502 77782 -2266
rect 77866 -2502 78102 -2266
rect 77546 -2822 77782 -2586
rect 77866 -2822 78102 -2586
rect 81266 -4422 81502 -4186
rect 81586 -4422 81822 -4186
rect 81266 -4742 81502 -4506
rect 81586 -4742 81822 -4506
rect 66986 -7302 67222 -7066
rect 67306 -7302 67542 -7066
rect 66986 -7622 67222 -7386
rect 67306 -7622 67542 -7386
rect 95546 -3462 95782 -3226
rect 95866 -3462 96102 -3226
rect 95546 -3782 95782 -3546
rect 95866 -3782 96102 -3546
rect 99266 -5382 99502 -5146
rect 99586 -5382 99822 -5146
rect 99266 -5702 99502 -5466
rect 99586 -5702 99822 -5466
rect 84986 -6342 85222 -6106
rect 85306 -6342 85542 -6106
rect 84986 -6662 85222 -6426
rect 85306 -6662 85542 -6426
rect 113546 -2502 113782 -2266
rect 113866 -2502 114102 -2266
rect 113546 -2822 113782 -2586
rect 113866 -2822 114102 -2586
rect 117266 -4422 117502 -4186
rect 117586 -4422 117822 -4186
rect 117266 -4742 117502 -4506
rect 117586 -4742 117822 -4506
rect 102986 -7302 103222 -7066
rect 103306 -7302 103542 -7066
rect 102986 -7622 103222 -7386
rect 103306 -7622 103542 -7386
rect 131546 -3462 131782 -3226
rect 131866 -3462 132102 -3226
rect 131546 -3782 131782 -3546
rect 131866 -3782 132102 -3546
rect 135266 -5382 135502 -5146
rect 135586 -5382 135822 -5146
rect 135266 -5702 135502 -5466
rect 135586 -5702 135822 -5466
rect 120986 -6342 121222 -6106
rect 121306 -6342 121542 -6106
rect 120986 -6662 121222 -6426
rect 121306 -6662 121542 -6426
rect 149546 -2502 149782 -2266
rect 149866 -2502 150102 -2266
rect 149546 -2822 149782 -2586
rect 149866 -2822 150102 -2586
rect 153266 -4422 153502 -4186
rect 153586 -4422 153822 -4186
rect 153266 -4742 153502 -4506
rect 153586 -4742 153822 -4506
rect 138986 -7302 139222 -7066
rect 139306 -7302 139542 -7066
rect 138986 -7622 139222 -7386
rect 139306 -7622 139542 -7386
rect 167546 -3462 167782 -3226
rect 167866 -3462 168102 -3226
rect 167546 -3782 167782 -3546
rect 167866 -3782 168102 -3546
rect 171266 -5382 171502 -5146
rect 171586 -5382 171822 -5146
rect 171266 -5702 171502 -5466
rect 171586 -5702 171822 -5466
rect 156986 -6342 157222 -6106
rect 157306 -6342 157542 -6106
rect 156986 -6662 157222 -6426
rect 157306 -6662 157542 -6426
rect 185546 -2502 185782 -2266
rect 185866 -2502 186102 -2266
rect 185546 -2822 185782 -2586
rect 185866 -2822 186102 -2586
rect 189266 -4422 189502 -4186
rect 189586 -4422 189822 -4186
rect 189266 -4742 189502 -4506
rect 189586 -4742 189822 -4506
rect 174986 -7302 175222 -7066
rect 175306 -7302 175542 -7066
rect 174986 -7622 175222 -7386
rect 175306 -7622 175542 -7386
rect 203546 -3462 203782 -3226
rect 203866 -3462 204102 -3226
rect 203546 -3782 203782 -3546
rect 203866 -3782 204102 -3546
rect 207266 -5382 207502 -5146
rect 207586 -5382 207822 -5146
rect 207266 -5702 207502 -5466
rect 207586 -5702 207822 -5466
rect 192986 -6342 193222 -6106
rect 193306 -6342 193542 -6106
rect 192986 -6662 193222 -6426
rect 193306 -6662 193542 -6426
rect 221546 -2502 221782 -2266
rect 221866 -2502 222102 -2266
rect 221546 -2822 221782 -2586
rect 221866 -2822 222102 -2586
rect 225266 -4422 225502 -4186
rect 225586 -4422 225822 -4186
rect 225266 -4742 225502 -4506
rect 225586 -4742 225822 -4506
rect 210986 -7302 211222 -7066
rect 211306 -7302 211542 -7066
rect 210986 -7622 211222 -7386
rect 211306 -7622 211542 -7386
rect 239546 -3462 239782 -3226
rect 239866 -3462 240102 -3226
rect 239546 -3782 239782 -3546
rect 239866 -3782 240102 -3546
rect 243266 -5382 243502 -5146
rect 243586 -5382 243822 -5146
rect 243266 -5702 243502 -5466
rect 243586 -5702 243822 -5466
rect 228986 -6342 229222 -6106
rect 229306 -6342 229542 -6106
rect 228986 -6662 229222 -6426
rect 229306 -6662 229542 -6426
rect 257546 -2502 257782 -2266
rect 257866 -2502 258102 -2266
rect 257546 -2822 257782 -2586
rect 257866 -2822 258102 -2586
rect 261266 -4422 261502 -4186
rect 261586 -4422 261822 -4186
rect 261266 -4742 261502 -4506
rect 261586 -4742 261822 -4506
rect 246986 -7302 247222 -7066
rect 247306 -7302 247542 -7066
rect 246986 -7622 247222 -7386
rect 247306 -7622 247542 -7386
rect 275546 -3462 275782 -3226
rect 275866 -3462 276102 -3226
rect 275546 -3782 275782 -3546
rect 275866 -3782 276102 -3546
rect 279266 -5382 279502 -5146
rect 279586 -5382 279822 -5146
rect 279266 -5702 279502 -5466
rect 279586 -5702 279822 -5466
rect 264986 -6342 265222 -6106
rect 265306 -6342 265542 -6106
rect 264986 -6662 265222 -6426
rect 265306 -6662 265542 -6426
rect 293546 -2502 293782 -2266
rect 293866 -2502 294102 -2266
rect 293546 -2822 293782 -2586
rect 293866 -2822 294102 -2586
rect 297266 -4422 297502 -4186
rect 297586 -4422 297822 -4186
rect 297266 -4742 297502 -4506
rect 297586 -4742 297822 -4506
rect 282986 -7302 283222 -7066
rect 283306 -7302 283542 -7066
rect 282986 -7622 283222 -7386
rect 283306 -7622 283542 -7386
rect 311546 -3462 311782 -3226
rect 311866 -3462 312102 -3226
rect 311546 -3782 311782 -3546
rect 311866 -3782 312102 -3546
rect 315266 -5382 315502 -5146
rect 315586 -5382 315822 -5146
rect 315266 -5702 315502 -5466
rect 315586 -5702 315822 -5466
rect 300986 -6342 301222 -6106
rect 301306 -6342 301542 -6106
rect 300986 -6662 301222 -6426
rect 301306 -6662 301542 -6426
rect 329546 -2502 329782 -2266
rect 329866 -2502 330102 -2266
rect 329546 -2822 329782 -2586
rect 329866 -2822 330102 -2586
rect 333266 -4422 333502 -4186
rect 333586 -4422 333822 -4186
rect 333266 -4742 333502 -4506
rect 333586 -4742 333822 -4506
rect 318986 -7302 319222 -7066
rect 319306 -7302 319542 -7066
rect 318986 -7622 319222 -7386
rect 319306 -7622 319542 -7386
rect 347546 -3462 347782 -3226
rect 347866 -3462 348102 -3226
rect 347546 -3782 347782 -3546
rect 347866 -3782 348102 -3546
rect 351266 -5382 351502 -5146
rect 351586 -5382 351822 -5146
rect 351266 -5702 351502 -5466
rect 351586 -5702 351822 -5466
rect 336986 -6342 337222 -6106
rect 337306 -6342 337542 -6106
rect 336986 -6662 337222 -6426
rect 337306 -6662 337542 -6426
rect 365546 -2502 365782 -2266
rect 365866 -2502 366102 -2266
rect 365546 -2822 365782 -2586
rect 365866 -2822 366102 -2586
rect 369266 -4422 369502 -4186
rect 369586 -4422 369822 -4186
rect 369266 -4742 369502 -4506
rect 369586 -4742 369822 -4506
rect 354986 -7302 355222 -7066
rect 355306 -7302 355542 -7066
rect 354986 -7622 355222 -7386
rect 355306 -7622 355542 -7386
rect 383546 -3462 383782 -3226
rect 383866 -3462 384102 -3226
rect 383546 -3782 383782 -3546
rect 383866 -3782 384102 -3546
rect 387266 -5382 387502 -5146
rect 387586 -5382 387822 -5146
rect 387266 -5702 387502 -5466
rect 387586 -5702 387822 -5466
rect 372986 -6342 373222 -6106
rect 373306 -6342 373542 -6106
rect 372986 -6662 373222 -6426
rect 373306 -6662 373542 -6426
rect 401546 -2502 401782 -2266
rect 401866 -2502 402102 -2266
rect 401546 -2822 401782 -2586
rect 401866 -2822 402102 -2586
rect 405266 -4422 405502 -4186
rect 405586 -4422 405822 -4186
rect 405266 -4742 405502 -4506
rect 405586 -4742 405822 -4506
rect 390986 -7302 391222 -7066
rect 391306 -7302 391542 -7066
rect 390986 -7622 391222 -7386
rect 391306 -7622 391542 -7386
rect 419546 -3462 419782 -3226
rect 419866 -3462 420102 -3226
rect 419546 -3782 419782 -3546
rect 419866 -3782 420102 -3546
rect 423266 -5382 423502 -5146
rect 423586 -5382 423822 -5146
rect 423266 -5702 423502 -5466
rect 423586 -5702 423822 -5466
rect 408986 -6342 409222 -6106
rect 409306 -6342 409542 -6106
rect 408986 -6662 409222 -6426
rect 409306 -6662 409542 -6426
rect 437546 -2502 437782 -2266
rect 437866 -2502 438102 -2266
rect 437546 -2822 437782 -2586
rect 437866 -2822 438102 -2586
rect 441266 -4422 441502 -4186
rect 441586 -4422 441822 -4186
rect 441266 -4742 441502 -4506
rect 441586 -4742 441822 -4506
rect 426986 -7302 427222 -7066
rect 427306 -7302 427542 -7066
rect 426986 -7622 427222 -7386
rect 427306 -7622 427542 -7386
rect 455546 -3462 455782 -3226
rect 455866 -3462 456102 -3226
rect 455546 -3782 455782 -3546
rect 455866 -3782 456102 -3546
rect 459266 -5382 459502 -5146
rect 459586 -5382 459822 -5146
rect 459266 -5702 459502 -5466
rect 459586 -5702 459822 -5466
rect 444986 -6342 445222 -6106
rect 445306 -6342 445542 -6106
rect 444986 -6662 445222 -6426
rect 445306 -6662 445542 -6426
rect 473546 -2502 473782 -2266
rect 473866 -2502 474102 -2266
rect 473546 -2822 473782 -2586
rect 473866 -2822 474102 -2586
rect 477266 -4422 477502 -4186
rect 477586 -4422 477822 -4186
rect 477266 -4742 477502 -4506
rect 477586 -4742 477822 -4506
rect 462986 -7302 463222 -7066
rect 463306 -7302 463542 -7066
rect 462986 -7622 463222 -7386
rect 463306 -7622 463542 -7386
rect 491546 -3462 491782 -3226
rect 491866 -3462 492102 -3226
rect 491546 -3782 491782 -3546
rect 491866 -3782 492102 -3546
rect 495266 -5382 495502 -5146
rect 495586 -5382 495822 -5146
rect 495266 -5702 495502 -5466
rect 495586 -5702 495822 -5466
rect 480986 -6342 481222 -6106
rect 481306 -6342 481542 -6106
rect 480986 -6662 481222 -6426
rect 481306 -6662 481542 -6426
rect 509546 -2502 509782 -2266
rect 509866 -2502 510102 -2266
rect 509546 -2822 509782 -2586
rect 509866 -2822 510102 -2586
rect 513266 -4422 513502 -4186
rect 513586 -4422 513822 -4186
rect 513266 -4742 513502 -4506
rect 513586 -4742 513822 -4506
rect 498986 -7302 499222 -7066
rect 499306 -7302 499542 -7066
rect 498986 -7622 499222 -7386
rect 499306 -7622 499542 -7386
rect 527546 -3462 527782 -3226
rect 527866 -3462 528102 -3226
rect 527546 -3782 527782 -3546
rect 527866 -3782 528102 -3546
rect 531266 -5382 531502 -5146
rect 531586 -5382 531822 -5146
rect 531266 -5702 531502 -5466
rect 531586 -5702 531822 -5466
rect 516986 -6342 517222 -6106
rect 517306 -6342 517542 -6106
rect 516986 -6662 517222 -6426
rect 517306 -6662 517542 -6426
rect 545546 -2502 545782 -2266
rect 545866 -2502 546102 -2266
rect 545546 -2822 545782 -2586
rect 545866 -2822 546102 -2586
rect 549266 -4422 549502 -4186
rect 549586 -4422 549822 -4186
rect 549266 -4742 549502 -4506
rect 549586 -4742 549822 -4506
rect 534986 -7302 535222 -7066
rect 535306 -7302 535542 -7066
rect 534986 -7622 535222 -7386
rect 535306 -7622 535542 -7386
rect 563546 -3462 563782 -3226
rect 563866 -3462 564102 -3226
rect 563546 -3782 563782 -3546
rect 563866 -3782 564102 -3546
rect 567266 -5382 567502 -5146
rect 567586 -5382 567822 -5146
rect 567266 -5702 567502 -5466
rect 567586 -5702 567822 -5466
rect 592062 711322 592298 711558
rect 592382 711322 592618 711558
rect 592062 711002 592298 711238
rect 592382 711002 592618 711238
rect 591102 710362 591338 710598
rect 591422 710362 591658 710598
rect 591102 710042 591338 710278
rect 591422 710042 591658 710278
rect 590142 709402 590378 709638
rect 590462 709402 590698 709638
rect 590142 709082 590378 709318
rect 590462 709082 590698 709318
rect 589182 708442 589418 708678
rect 589502 708442 589738 708678
rect 589182 708122 589418 708358
rect 589502 708122 589738 708358
rect 588222 707482 588458 707718
rect 588542 707482 588778 707718
rect 588222 707162 588458 707398
rect 588542 707162 588778 707398
rect 581546 706522 581782 706758
rect 581866 706522 582102 706758
rect 581546 706202 581782 706438
rect 581866 706202 582102 706438
rect 570986 680378 571222 680614
rect 571306 680378 571542 680614
rect 570986 680058 571222 680294
rect 571306 680058 571542 680294
rect 570986 644378 571222 644614
rect 571306 644378 571542 644614
rect 570986 644058 571222 644294
rect 571306 644058 571542 644294
rect 570986 608378 571222 608614
rect 571306 608378 571542 608614
rect 570986 608058 571222 608294
rect 571306 608058 571542 608294
rect 570986 572378 571222 572614
rect 571306 572378 571542 572614
rect 570986 572058 571222 572294
rect 571306 572058 571542 572294
rect 570986 536378 571222 536614
rect 571306 536378 571542 536614
rect 570986 536058 571222 536294
rect 571306 536058 571542 536294
rect 570986 500378 571222 500614
rect 571306 500378 571542 500614
rect 570986 500058 571222 500294
rect 571306 500058 571542 500294
rect 570986 464378 571222 464614
rect 571306 464378 571542 464614
rect 570986 464058 571222 464294
rect 571306 464058 571542 464294
rect 570986 428378 571222 428614
rect 571306 428378 571542 428614
rect 570986 428058 571222 428294
rect 571306 428058 571542 428294
rect 570986 392378 571222 392614
rect 571306 392378 571542 392614
rect 570986 392058 571222 392294
rect 571306 392058 571542 392294
rect 570986 356378 571222 356614
rect 571306 356378 571542 356614
rect 570986 356058 571222 356294
rect 571306 356058 571542 356294
rect 570986 320378 571222 320614
rect 571306 320378 571542 320614
rect 570986 320058 571222 320294
rect 571306 320058 571542 320294
rect 570986 284378 571222 284614
rect 571306 284378 571542 284614
rect 570986 284058 571222 284294
rect 571306 284058 571542 284294
rect 570986 248378 571222 248614
rect 571306 248378 571542 248614
rect 570986 248058 571222 248294
rect 571306 248058 571542 248294
rect 570986 212378 571222 212614
rect 571306 212378 571542 212614
rect 570986 212058 571222 212294
rect 571306 212058 571542 212294
rect 570986 176378 571222 176614
rect 571306 176378 571542 176614
rect 570986 176058 571222 176294
rect 571306 176058 571542 176294
rect 570986 140378 571222 140614
rect 571306 140378 571542 140614
rect 570986 140058 571222 140294
rect 571306 140058 571542 140294
rect 570986 104378 571222 104614
rect 571306 104378 571542 104614
rect 570986 104058 571222 104294
rect 571306 104058 571542 104294
rect 570986 68378 571222 68614
rect 571306 68378 571542 68614
rect 570986 68058 571222 68294
rect 571306 68058 571542 68294
rect 570986 32378 571222 32614
rect 571306 32378 571542 32614
rect 570986 32058 571222 32294
rect 571306 32058 571542 32294
rect 552986 -6342 553222 -6106
rect 553306 -6342 553542 -6106
rect 552986 -6662 553222 -6426
rect 553306 -6662 553542 -6426
rect 577826 704602 578062 704838
rect 578146 704602 578382 704838
rect 577826 704282 578062 704518
rect 578146 704282 578382 704518
rect 577826 687218 578062 687454
rect 578146 687218 578382 687454
rect 577826 686898 578062 687134
rect 578146 686898 578382 687134
rect 577826 651218 578062 651454
rect 578146 651218 578382 651454
rect 577826 650898 578062 651134
rect 578146 650898 578382 651134
rect 577826 615218 578062 615454
rect 578146 615218 578382 615454
rect 577826 614898 578062 615134
rect 578146 614898 578382 615134
rect 577826 579218 578062 579454
rect 578146 579218 578382 579454
rect 577826 578898 578062 579134
rect 578146 578898 578382 579134
rect 577826 543218 578062 543454
rect 578146 543218 578382 543454
rect 577826 542898 578062 543134
rect 578146 542898 578382 543134
rect 577826 507218 578062 507454
rect 578146 507218 578382 507454
rect 577826 506898 578062 507134
rect 578146 506898 578382 507134
rect 577826 471218 578062 471454
rect 578146 471218 578382 471454
rect 577826 470898 578062 471134
rect 578146 470898 578382 471134
rect 577826 435218 578062 435454
rect 578146 435218 578382 435454
rect 577826 434898 578062 435134
rect 578146 434898 578382 435134
rect 577826 399218 578062 399454
rect 578146 399218 578382 399454
rect 577826 398898 578062 399134
rect 578146 398898 578382 399134
rect 577826 363218 578062 363454
rect 578146 363218 578382 363454
rect 577826 362898 578062 363134
rect 578146 362898 578382 363134
rect 577826 327218 578062 327454
rect 578146 327218 578382 327454
rect 577826 326898 578062 327134
rect 578146 326898 578382 327134
rect 577826 291218 578062 291454
rect 578146 291218 578382 291454
rect 577826 290898 578062 291134
rect 578146 290898 578382 291134
rect 577826 255218 578062 255454
rect 578146 255218 578382 255454
rect 577826 254898 578062 255134
rect 578146 254898 578382 255134
rect 577826 219218 578062 219454
rect 578146 219218 578382 219454
rect 577826 218898 578062 219134
rect 578146 218898 578382 219134
rect 577826 183218 578062 183454
rect 578146 183218 578382 183454
rect 577826 182898 578062 183134
rect 578146 182898 578382 183134
rect 577826 147218 578062 147454
rect 578146 147218 578382 147454
rect 577826 146898 578062 147134
rect 578146 146898 578382 147134
rect 577826 111218 578062 111454
rect 578146 111218 578382 111454
rect 577826 110898 578062 111134
rect 578146 110898 578382 111134
rect 577826 75218 578062 75454
rect 578146 75218 578382 75454
rect 577826 74898 578062 75134
rect 578146 74898 578382 75134
rect 577826 39218 578062 39454
rect 578146 39218 578382 39454
rect 577826 38898 578062 39134
rect 578146 38898 578382 39134
rect 577826 3218 578062 3454
rect 578146 3218 578382 3454
rect 577826 2898 578062 3134
rect 578146 2898 578382 3134
rect 577826 -582 578062 -346
rect 578146 -582 578382 -346
rect 577826 -902 578062 -666
rect 578146 -902 578382 -666
rect 587262 706522 587498 706758
rect 587582 706522 587818 706758
rect 587262 706202 587498 706438
rect 587582 706202 587818 706438
rect 586302 705562 586538 705798
rect 586622 705562 586858 705798
rect 586302 705242 586538 705478
rect 586622 705242 586858 705478
rect 581546 690938 581782 691174
rect 581866 690938 582102 691174
rect 581546 690618 581782 690854
rect 581866 690618 582102 690854
rect 581546 654938 581782 655174
rect 581866 654938 582102 655174
rect 581546 654618 581782 654854
rect 581866 654618 582102 654854
rect 581546 618938 581782 619174
rect 581866 618938 582102 619174
rect 581546 618618 581782 618854
rect 581866 618618 582102 618854
rect 581546 582938 581782 583174
rect 581866 582938 582102 583174
rect 581546 582618 581782 582854
rect 581866 582618 582102 582854
rect 581546 546938 581782 547174
rect 581866 546938 582102 547174
rect 581546 546618 581782 546854
rect 581866 546618 582102 546854
rect 581546 510938 581782 511174
rect 581866 510938 582102 511174
rect 581546 510618 581782 510854
rect 581866 510618 582102 510854
rect 581546 474938 581782 475174
rect 581866 474938 582102 475174
rect 581546 474618 581782 474854
rect 581866 474618 582102 474854
rect 581546 438938 581782 439174
rect 581866 438938 582102 439174
rect 581546 438618 581782 438854
rect 581866 438618 582102 438854
rect 581546 402938 581782 403174
rect 581866 402938 582102 403174
rect 581546 402618 581782 402854
rect 581866 402618 582102 402854
rect 581546 366938 581782 367174
rect 581866 366938 582102 367174
rect 581546 366618 581782 366854
rect 581866 366618 582102 366854
rect 581546 330938 581782 331174
rect 581866 330938 582102 331174
rect 581546 330618 581782 330854
rect 581866 330618 582102 330854
rect 581546 294938 581782 295174
rect 581866 294938 582102 295174
rect 581546 294618 581782 294854
rect 581866 294618 582102 294854
rect 581546 258938 581782 259174
rect 581866 258938 582102 259174
rect 581546 258618 581782 258854
rect 581866 258618 582102 258854
rect 581546 222938 581782 223174
rect 581866 222938 582102 223174
rect 581546 222618 581782 222854
rect 581866 222618 582102 222854
rect 581546 186938 581782 187174
rect 581866 186938 582102 187174
rect 581546 186618 581782 186854
rect 581866 186618 582102 186854
rect 581546 150938 581782 151174
rect 581866 150938 582102 151174
rect 581546 150618 581782 150854
rect 581866 150618 582102 150854
rect 581546 114938 581782 115174
rect 581866 114938 582102 115174
rect 581546 114618 581782 114854
rect 581866 114618 582102 114854
rect 581546 78938 581782 79174
rect 581866 78938 582102 79174
rect 581546 78618 581782 78854
rect 581866 78618 582102 78854
rect 581546 42938 581782 43174
rect 581866 42938 582102 43174
rect 581546 42618 581782 42854
rect 581866 42618 582102 42854
rect 581546 6938 581782 7174
rect 581866 6938 582102 7174
rect 581546 6618 581782 6854
rect 581866 6618 582102 6854
rect 585342 704602 585578 704838
rect 585662 704602 585898 704838
rect 585342 704282 585578 704518
rect 585662 704282 585898 704518
rect 585342 687218 585578 687454
rect 585662 687218 585898 687454
rect 585342 686898 585578 687134
rect 585662 686898 585898 687134
rect 585342 651218 585578 651454
rect 585662 651218 585898 651454
rect 585342 650898 585578 651134
rect 585662 650898 585898 651134
rect 585342 615218 585578 615454
rect 585662 615218 585898 615454
rect 585342 614898 585578 615134
rect 585662 614898 585898 615134
rect 585342 579218 585578 579454
rect 585662 579218 585898 579454
rect 585342 578898 585578 579134
rect 585662 578898 585898 579134
rect 585342 543218 585578 543454
rect 585662 543218 585898 543454
rect 585342 542898 585578 543134
rect 585662 542898 585898 543134
rect 585342 507218 585578 507454
rect 585662 507218 585898 507454
rect 585342 506898 585578 507134
rect 585662 506898 585898 507134
rect 585342 471218 585578 471454
rect 585662 471218 585898 471454
rect 585342 470898 585578 471134
rect 585662 470898 585898 471134
rect 585342 435218 585578 435454
rect 585662 435218 585898 435454
rect 585342 434898 585578 435134
rect 585662 434898 585898 435134
rect 585342 399218 585578 399454
rect 585662 399218 585898 399454
rect 585342 398898 585578 399134
rect 585662 398898 585898 399134
rect 585342 363218 585578 363454
rect 585662 363218 585898 363454
rect 585342 362898 585578 363134
rect 585662 362898 585898 363134
rect 585342 327218 585578 327454
rect 585662 327218 585898 327454
rect 585342 326898 585578 327134
rect 585662 326898 585898 327134
rect 585342 291218 585578 291454
rect 585662 291218 585898 291454
rect 585342 290898 585578 291134
rect 585662 290898 585898 291134
rect 585342 255218 585578 255454
rect 585662 255218 585898 255454
rect 585342 254898 585578 255134
rect 585662 254898 585898 255134
rect 585342 219218 585578 219454
rect 585662 219218 585898 219454
rect 585342 218898 585578 219134
rect 585662 218898 585898 219134
rect 585342 183218 585578 183454
rect 585662 183218 585898 183454
rect 585342 182898 585578 183134
rect 585662 182898 585898 183134
rect 585342 147218 585578 147454
rect 585662 147218 585898 147454
rect 585342 146898 585578 147134
rect 585662 146898 585898 147134
rect 585342 111218 585578 111454
rect 585662 111218 585898 111454
rect 585342 110898 585578 111134
rect 585662 110898 585898 111134
rect 585342 75218 585578 75454
rect 585662 75218 585898 75454
rect 585342 74898 585578 75134
rect 585662 74898 585898 75134
rect 585342 39218 585578 39454
rect 585662 39218 585898 39454
rect 585342 38898 585578 39134
rect 585662 38898 585898 39134
rect 585342 3218 585578 3454
rect 585662 3218 585898 3454
rect 585342 2898 585578 3134
rect 585662 2898 585898 3134
rect 585342 -582 585578 -346
rect 585662 -582 585898 -346
rect 585342 -902 585578 -666
rect 585662 -902 585898 -666
rect 586302 669218 586538 669454
rect 586622 669218 586858 669454
rect 586302 668898 586538 669134
rect 586622 668898 586858 669134
rect 586302 633218 586538 633454
rect 586622 633218 586858 633454
rect 586302 632898 586538 633134
rect 586622 632898 586858 633134
rect 586302 597218 586538 597454
rect 586622 597218 586858 597454
rect 586302 596898 586538 597134
rect 586622 596898 586858 597134
rect 586302 561218 586538 561454
rect 586622 561218 586858 561454
rect 586302 560898 586538 561134
rect 586622 560898 586858 561134
rect 586302 525218 586538 525454
rect 586622 525218 586858 525454
rect 586302 524898 586538 525134
rect 586622 524898 586858 525134
rect 586302 489218 586538 489454
rect 586622 489218 586858 489454
rect 586302 488898 586538 489134
rect 586622 488898 586858 489134
rect 586302 453218 586538 453454
rect 586622 453218 586858 453454
rect 586302 452898 586538 453134
rect 586622 452898 586858 453134
rect 586302 417218 586538 417454
rect 586622 417218 586858 417454
rect 586302 416898 586538 417134
rect 586622 416898 586858 417134
rect 586302 381218 586538 381454
rect 586622 381218 586858 381454
rect 586302 380898 586538 381134
rect 586622 380898 586858 381134
rect 586302 345218 586538 345454
rect 586622 345218 586858 345454
rect 586302 344898 586538 345134
rect 586622 344898 586858 345134
rect 586302 309218 586538 309454
rect 586622 309218 586858 309454
rect 586302 308898 586538 309134
rect 586622 308898 586858 309134
rect 586302 273218 586538 273454
rect 586622 273218 586858 273454
rect 586302 272898 586538 273134
rect 586622 272898 586858 273134
rect 586302 237218 586538 237454
rect 586622 237218 586858 237454
rect 586302 236898 586538 237134
rect 586622 236898 586858 237134
rect 586302 201218 586538 201454
rect 586622 201218 586858 201454
rect 586302 200898 586538 201134
rect 586622 200898 586858 201134
rect 586302 165218 586538 165454
rect 586622 165218 586858 165454
rect 586302 164898 586538 165134
rect 586622 164898 586858 165134
rect 586302 129218 586538 129454
rect 586622 129218 586858 129454
rect 586302 128898 586538 129134
rect 586622 128898 586858 129134
rect 586302 93218 586538 93454
rect 586622 93218 586858 93454
rect 586302 92898 586538 93134
rect 586622 92898 586858 93134
rect 586302 57218 586538 57454
rect 586622 57218 586858 57454
rect 586302 56898 586538 57134
rect 586622 56898 586858 57134
rect 586302 21218 586538 21454
rect 586622 21218 586858 21454
rect 586302 20898 586538 21134
rect 586622 20898 586858 21134
rect 586302 -1542 586538 -1306
rect 586622 -1542 586858 -1306
rect 586302 -1862 586538 -1626
rect 586622 -1862 586858 -1626
rect 587262 690938 587498 691174
rect 587582 690938 587818 691174
rect 587262 690618 587498 690854
rect 587582 690618 587818 690854
rect 587262 654938 587498 655174
rect 587582 654938 587818 655174
rect 587262 654618 587498 654854
rect 587582 654618 587818 654854
rect 587262 618938 587498 619174
rect 587582 618938 587818 619174
rect 587262 618618 587498 618854
rect 587582 618618 587818 618854
rect 587262 582938 587498 583174
rect 587582 582938 587818 583174
rect 587262 582618 587498 582854
rect 587582 582618 587818 582854
rect 587262 546938 587498 547174
rect 587582 546938 587818 547174
rect 587262 546618 587498 546854
rect 587582 546618 587818 546854
rect 587262 510938 587498 511174
rect 587582 510938 587818 511174
rect 587262 510618 587498 510854
rect 587582 510618 587818 510854
rect 587262 474938 587498 475174
rect 587582 474938 587818 475174
rect 587262 474618 587498 474854
rect 587582 474618 587818 474854
rect 587262 438938 587498 439174
rect 587582 438938 587818 439174
rect 587262 438618 587498 438854
rect 587582 438618 587818 438854
rect 587262 402938 587498 403174
rect 587582 402938 587818 403174
rect 587262 402618 587498 402854
rect 587582 402618 587818 402854
rect 587262 366938 587498 367174
rect 587582 366938 587818 367174
rect 587262 366618 587498 366854
rect 587582 366618 587818 366854
rect 587262 330938 587498 331174
rect 587582 330938 587818 331174
rect 587262 330618 587498 330854
rect 587582 330618 587818 330854
rect 587262 294938 587498 295174
rect 587582 294938 587818 295174
rect 587262 294618 587498 294854
rect 587582 294618 587818 294854
rect 587262 258938 587498 259174
rect 587582 258938 587818 259174
rect 587262 258618 587498 258854
rect 587582 258618 587818 258854
rect 587262 222938 587498 223174
rect 587582 222938 587818 223174
rect 587262 222618 587498 222854
rect 587582 222618 587818 222854
rect 587262 186938 587498 187174
rect 587582 186938 587818 187174
rect 587262 186618 587498 186854
rect 587582 186618 587818 186854
rect 587262 150938 587498 151174
rect 587582 150938 587818 151174
rect 587262 150618 587498 150854
rect 587582 150618 587818 150854
rect 587262 114938 587498 115174
rect 587582 114938 587818 115174
rect 587262 114618 587498 114854
rect 587582 114618 587818 114854
rect 587262 78938 587498 79174
rect 587582 78938 587818 79174
rect 587262 78618 587498 78854
rect 587582 78618 587818 78854
rect 587262 42938 587498 43174
rect 587582 42938 587818 43174
rect 587262 42618 587498 42854
rect 587582 42618 587818 42854
rect 587262 6938 587498 7174
rect 587582 6938 587818 7174
rect 587262 6618 587498 6854
rect 587582 6618 587818 6854
rect 581546 -2502 581782 -2266
rect 581866 -2502 582102 -2266
rect 581546 -2822 581782 -2586
rect 581866 -2822 582102 -2586
rect 587262 -2502 587498 -2266
rect 587582 -2502 587818 -2266
rect 587262 -2822 587498 -2586
rect 587582 -2822 587818 -2586
rect 588222 672938 588458 673174
rect 588542 672938 588778 673174
rect 588222 672618 588458 672854
rect 588542 672618 588778 672854
rect 588222 636938 588458 637174
rect 588542 636938 588778 637174
rect 588222 636618 588458 636854
rect 588542 636618 588778 636854
rect 588222 600938 588458 601174
rect 588542 600938 588778 601174
rect 588222 600618 588458 600854
rect 588542 600618 588778 600854
rect 588222 564938 588458 565174
rect 588542 564938 588778 565174
rect 588222 564618 588458 564854
rect 588542 564618 588778 564854
rect 588222 528938 588458 529174
rect 588542 528938 588778 529174
rect 588222 528618 588458 528854
rect 588542 528618 588778 528854
rect 588222 492938 588458 493174
rect 588542 492938 588778 493174
rect 588222 492618 588458 492854
rect 588542 492618 588778 492854
rect 588222 456938 588458 457174
rect 588542 456938 588778 457174
rect 588222 456618 588458 456854
rect 588542 456618 588778 456854
rect 588222 420938 588458 421174
rect 588542 420938 588778 421174
rect 588222 420618 588458 420854
rect 588542 420618 588778 420854
rect 588222 384938 588458 385174
rect 588542 384938 588778 385174
rect 588222 384618 588458 384854
rect 588542 384618 588778 384854
rect 588222 348938 588458 349174
rect 588542 348938 588778 349174
rect 588222 348618 588458 348854
rect 588542 348618 588778 348854
rect 588222 312938 588458 313174
rect 588542 312938 588778 313174
rect 588222 312618 588458 312854
rect 588542 312618 588778 312854
rect 588222 276938 588458 277174
rect 588542 276938 588778 277174
rect 588222 276618 588458 276854
rect 588542 276618 588778 276854
rect 588222 240938 588458 241174
rect 588542 240938 588778 241174
rect 588222 240618 588458 240854
rect 588542 240618 588778 240854
rect 588222 204938 588458 205174
rect 588542 204938 588778 205174
rect 588222 204618 588458 204854
rect 588542 204618 588778 204854
rect 588222 168938 588458 169174
rect 588542 168938 588778 169174
rect 588222 168618 588458 168854
rect 588542 168618 588778 168854
rect 588222 132938 588458 133174
rect 588542 132938 588778 133174
rect 588222 132618 588458 132854
rect 588542 132618 588778 132854
rect 588222 96938 588458 97174
rect 588542 96938 588778 97174
rect 588222 96618 588458 96854
rect 588542 96618 588778 96854
rect 588222 60938 588458 61174
rect 588542 60938 588778 61174
rect 588222 60618 588458 60854
rect 588542 60618 588778 60854
rect 588222 24938 588458 25174
rect 588542 24938 588778 25174
rect 588222 24618 588458 24854
rect 588542 24618 588778 24854
rect 588222 -3462 588458 -3226
rect 588542 -3462 588778 -3226
rect 588222 -3782 588458 -3546
rect 588542 -3782 588778 -3546
rect 589182 694658 589418 694894
rect 589502 694658 589738 694894
rect 589182 694338 589418 694574
rect 589502 694338 589738 694574
rect 589182 658658 589418 658894
rect 589502 658658 589738 658894
rect 589182 658338 589418 658574
rect 589502 658338 589738 658574
rect 589182 622658 589418 622894
rect 589502 622658 589738 622894
rect 589182 622338 589418 622574
rect 589502 622338 589738 622574
rect 589182 586658 589418 586894
rect 589502 586658 589738 586894
rect 589182 586338 589418 586574
rect 589502 586338 589738 586574
rect 589182 550658 589418 550894
rect 589502 550658 589738 550894
rect 589182 550338 589418 550574
rect 589502 550338 589738 550574
rect 589182 514658 589418 514894
rect 589502 514658 589738 514894
rect 589182 514338 589418 514574
rect 589502 514338 589738 514574
rect 589182 478658 589418 478894
rect 589502 478658 589738 478894
rect 589182 478338 589418 478574
rect 589502 478338 589738 478574
rect 589182 442658 589418 442894
rect 589502 442658 589738 442894
rect 589182 442338 589418 442574
rect 589502 442338 589738 442574
rect 589182 406658 589418 406894
rect 589502 406658 589738 406894
rect 589182 406338 589418 406574
rect 589502 406338 589738 406574
rect 589182 370658 589418 370894
rect 589502 370658 589738 370894
rect 589182 370338 589418 370574
rect 589502 370338 589738 370574
rect 589182 334658 589418 334894
rect 589502 334658 589738 334894
rect 589182 334338 589418 334574
rect 589502 334338 589738 334574
rect 589182 298658 589418 298894
rect 589502 298658 589738 298894
rect 589182 298338 589418 298574
rect 589502 298338 589738 298574
rect 589182 262658 589418 262894
rect 589502 262658 589738 262894
rect 589182 262338 589418 262574
rect 589502 262338 589738 262574
rect 589182 226658 589418 226894
rect 589502 226658 589738 226894
rect 589182 226338 589418 226574
rect 589502 226338 589738 226574
rect 589182 190658 589418 190894
rect 589502 190658 589738 190894
rect 589182 190338 589418 190574
rect 589502 190338 589738 190574
rect 589182 154658 589418 154894
rect 589502 154658 589738 154894
rect 589182 154338 589418 154574
rect 589502 154338 589738 154574
rect 589182 118658 589418 118894
rect 589502 118658 589738 118894
rect 589182 118338 589418 118574
rect 589502 118338 589738 118574
rect 589182 82658 589418 82894
rect 589502 82658 589738 82894
rect 589182 82338 589418 82574
rect 589502 82338 589738 82574
rect 589182 46658 589418 46894
rect 589502 46658 589738 46894
rect 589182 46338 589418 46574
rect 589502 46338 589738 46574
rect 589182 10658 589418 10894
rect 589502 10658 589738 10894
rect 589182 10338 589418 10574
rect 589502 10338 589738 10574
rect 589182 -4422 589418 -4186
rect 589502 -4422 589738 -4186
rect 589182 -4742 589418 -4506
rect 589502 -4742 589738 -4506
rect 590142 676658 590378 676894
rect 590462 676658 590698 676894
rect 590142 676338 590378 676574
rect 590462 676338 590698 676574
rect 590142 640658 590378 640894
rect 590462 640658 590698 640894
rect 590142 640338 590378 640574
rect 590462 640338 590698 640574
rect 590142 604658 590378 604894
rect 590462 604658 590698 604894
rect 590142 604338 590378 604574
rect 590462 604338 590698 604574
rect 590142 568658 590378 568894
rect 590462 568658 590698 568894
rect 590142 568338 590378 568574
rect 590462 568338 590698 568574
rect 590142 532658 590378 532894
rect 590462 532658 590698 532894
rect 590142 532338 590378 532574
rect 590462 532338 590698 532574
rect 590142 496658 590378 496894
rect 590462 496658 590698 496894
rect 590142 496338 590378 496574
rect 590462 496338 590698 496574
rect 590142 460658 590378 460894
rect 590462 460658 590698 460894
rect 590142 460338 590378 460574
rect 590462 460338 590698 460574
rect 590142 424658 590378 424894
rect 590462 424658 590698 424894
rect 590142 424338 590378 424574
rect 590462 424338 590698 424574
rect 590142 388658 590378 388894
rect 590462 388658 590698 388894
rect 590142 388338 590378 388574
rect 590462 388338 590698 388574
rect 590142 352658 590378 352894
rect 590462 352658 590698 352894
rect 590142 352338 590378 352574
rect 590462 352338 590698 352574
rect 590142 316658 590378 316894
rect 590462 316658 590698 316894
rect 590142 316338 590378 316574
rect 590462 316338 590698 316574
rect 590142 280658 590378 280894
rect 590462 280658 590698 280894
rect 590142 280338 590378 280574
rect 590462 280338 590698 280574
rect 590142 244658 590378 244894
rect 590462 244658 590698 244894
rect 590142 244338 590378 244574
rect 590462 244338 590698 244574
rect 590142 208658 590378 208894
rect 590462 208658 590698 208894
rect 590142 208338 590378 208574
rect 590462 208338 590698 208574
rect 590142 172658 590378 172894
rect 590462 172658 590698 172894
rect 590142 172338 590378 172574
rect 590462 172338 590698 172574
rect 590142 136658 590378 136894
rect 590462 136658 590698 136894
rect 590142 136338 590378 136574
rect 590462 136338 590698 136574
rect 590142 100658 590378 100894
rect 590462 100658 590698 100894
rect 590142 100338 590378 100574
rect 590462 100338 590698 100574
rect 590142 64658 590378 64894
rect 590462 64658 590698 64894
rect 590142 64338 590378 64574
rect 590462 64338 590698 64574
rect 590142 28658 590378 28894
rect 590462 28658 590698 28894
rect 590142 28338 590378 28574
rect 590462 28338 590698 28574
rect 590142 -5382 590378 -5146
rect 590462 -5382 590698 -5146
rect 590142 -5702 590378 -5466
rect 590462 -5702 590698 -5466
rect 591102 698378 591338 698614
rect 591422 698378 591658 698614
rect 591102 698058 591338 698294
rect 591422 698058 591658 698294
rect 591102 662378 591338 662614
rect 591422 662378 591658 662614
rect 591102 662058 591338 662294
rect 591422 662058 591658 662294
rect 591102 626378 591338 626614
rect 591422 626378 591658 626614
rect 591102 626058 591338 626294
rect 591422 626058 591658 626294
rect 591102 590378 591338 590614
rect 591422 590378 591658 590614
rect 591102 590058 591338 590294
rect 591422 590058 591658 590294
rect 591102 554378 591338 554614
rect 591422 554378 591658 554614
rect 591102 554058 591338 554294
rect 591422 554058 591658 554294
rect 591102 518378 591338 518614
rect 591422 518378 591658 518614
rect 591102 518058 591338 518294
rect 591422 518058 591658 518294
rect 591102 482378 591338 482614
rect 591422 482378 591658 482614
rect 591102 482058 591338 482294
rect 591422 482058 591658 482294
rect 591102 446378 591338 446614
rect 591422 446378 591658 446614
rect 591102 446058 591338 446294
rect 591422 446058 591658 446294
rect 591102 410378 591338 410614
rect 591422 410378 591658 410614
rect 591102 410058 591338 410294
rect 591422 410058 591658 410294
rect 591102 374378 591338 374614
rect 591422 374378 591658 374614
rect 591102 374058 591338 374294
rect 591422 374058 591658 374294
rect 591102 338378 591338 338614
rect 591422 338378 591658 338614
rect 591102 338058 591338 338294
rect 591422 338058 591658 338294
rect 591102 302378 591338 302614
rect 591422 302378 591658 302614
rect 591102 302058 591338 302294
rect 591422 302058 591658 302294
rect 591102 266378 591338 266614
rect 591422 266378 591658 266614
rect 591102 266058 591338 266294
rect 591422 266058 591658 266294
rect 591102 230378 591338 230614
rect 591422 230378 591658 230614
rect 591102 230058 591338 230294
rect 591422 230058 591658 230294
rect 591102 194378 591338 194614
rect 591422 194378 591658 194614
rect 591102 194058 591338 194294
rect 591422 194058 591658 194294
rect 591102 158378 591338 158614
rect 591422 158378 591658 158614
rect 591102 158058 591338 158294
rect 591422 158058 591658 158294
rect 591102 122378 591338 122614
rect 591422 122378 591658 122614
rect 591102 122058 591338 122294
rect 591422 122058 591658 122294
rect 591102 86378 591338 86614
rect 591422 86378 591658 86614
rect 591102 86058 591338 86294
rect 591422 86058 591658 86294
rect 591102 50378 591338 50614
rect 591422 50378 591658 50614
rect 591102 50058 591338 50294
rect 591422 50058 591658 50294
rect 591102 14378 591338 14614
rect 591422 14378 591658 14614
rect 591102 14058 591338 14294
rect 591422 14058 591658 14294
rect 591102 -6342 591338 -6106
rect 591422 -6342 591658 -6106
rect 591102 -6662 591338 -6426
rect 591422 -6662 591658 -6426
rect 592062 680378 592298 680614
rect 592382 680378 592618 680614
rect 592062 680058 592298 680294
rect 592382 680058 592618 680294
rect 592062 644378 592298 644614
rect 592382 644378 592618 644614
rect 592062 644058 592298 644294
rect 592382 644058 592618 644294
rect 592062 608378 592298 608614
rect 592382 608378 592618 608614
rect 592062 608058 592298 608294
rect 592382 608058 592618 608294
rect 592062 572378 592298 572614
rect 592382 572378 592618 572614
rect 592062 572058 592298 572294
rect 592382 572058 592618 572294
rect 592062 536378 592298 536614
rect 592382 536378 592618 536614
rect 592062 536058 592298 536294
rect 592382 536058 592618 536294
rect 592062 500378 592298 500614
rect 592382 500378 592618 500614
rect 592062 500058 592298 500294
rect 592382 500058 592618 500294
rect 592062 464378 592298 464614
rect 592382 464378 592618 464614
rect 592062 464058 592298 464294
rect 592382 464058 592618 464294
rect 592062 428378 592298 428614
rect 592382 428378 592618 428614
rect 592062 428058 592298 428294
rect 592382 428058 592618 428294
rect 592062 392378 592298 392614
rect 592382 392378 592618 392614
rect 592062 392058 592298 392294
rect 592382 392058 592618 392294
rect 592062 356378 592298 356614
rect 592382 356378 592618 356614
rect 592062 356058 592298 356294
rect 592382 356058 592618 356294
rect 592062 320378 592298 320614
rect 592382 320378 592618 320614
rect 592062 320058 592298 320294
rect 592382 320058 592618 320294
rect 592062 284378 592298 284614
rect 592382 284378 592618 284614
rect 592062 284058 592298 284294
rect 592382 284058 592618 284294
rect 592062 248378 592298 248614
rect 592382 248378 592618 248614
rect 592062 248058 592298 248294
rect 592382 248058 592618 248294
rect 592062 212378 592298 212614
rect 592382 212378 592618 212614
rect 592062 212058 592298 212294
rect 592382 212058 592618 212294
rect 592062 176378 592298 176614
rect 592382 176378 592618 176614
rect 592062 176058 592298 176294
rect 592382 176058 592618 176294
rect 592062 140378 592298 140614
rect 592382 140378 592618 140614
rect 592062 140058 592298 140294
rect 592382 140058 592618 140294
rect 592062 104378 592298 104614
rect 592382 104378 592618 104614
rect 592062 104058 592298 104294
rect 592382 104058 592618 104294
rect 592062 68378 592298 68614
rect 592382 68378 592618 68614
rect 592062 68058 592298 68294
rect 592382 68058 592618 68294
rect 592062 32378 592298 32614
rect 592382 32378 592618 32614
rect 592062 32058 592298 32294
rect 592382 32058 592618 32294
rect 570986 -7302 571222 -7066
rect 571306 -7302 571542 -7066
rect 570986 -7622 571222 -7386
rect 571306 -7622 571542 -7386
rect 592062 -7302 592298 -7066
rect 592382 -7302 592618 -7066
rect 592062 -7622 592298 -7386
rect 592382 -7622 592618 -7386
<< metal5 >>
rect -8726 711558 592650 711590
rect -8726 711322 -8694 711558
rect -8458 711322 -8374 711558
rect -8138 711322 30986 711558
rect 31222 711322 31306 711558
rect 31542 711322 66986 711558
rect 67222 711322 67306 711558
rect 67542 711322 102986 711558
rect 103222 711322 103306 711558
rect 103542 711322 138986 711558
rect 139222 711322 139306 711558
rect 139542 711322 174986 711558
rect 175222 711322 175306 711558
rect 175542 711322 210986 711558
rect 211222 711322 211306 711558
rect 211542 711322 246986 711558
rect 247222 711322 247306 711558
rect 247542 711322 282986 711558
rect 283222 711322 283306 711558
rect 283542 711322 318986 711558
rect 319222 711322 319306 711558
rect 319542 711322 354986 711558
rect 355222 711322 355306 711558
rect 355542 711322 390986 711558
rect 391222 711322 391306 711558
rect 391542 711322 426986 711558
rect 427222 711322 427306 711558
rect 427542 711322 462986 711558
rect 463222 711322 463306 711558
rect 463542 711322 498986 711558
rect 499222 711322 499306 711558
rect 499542 711322 534986 711558
rect 535222 711322 535306 711558
rect 535542 711322 570986 711558
rect 571222 711322 571306 711558
rect 571542 711322 592062 711558
rect 592298 711322 592382 711558
rect 592618 711322 592650 711558
rect -8726 711238 592650 711322
rect -8726 711002 -8694 711238
rect -8458 711002 -8374 711238
rect -8138 711002 30986 711238
rect 31222 711002 31306 711238
rect 31542 711002 66986 711238
rect 67222 711002 67306 711238
rect 67542 711002 102986 711238
rect 103222 711002 103306 711238
rect 103542 711002 138986 711238
rect 139222 711002 139306 711238
rect 139542 711002 174986 711238
rect 175222 711002 175306 711238
rect 175542 711002 210986 711238
rect 211222 711002 211306 711238
rect 211542 711002 246986 711238
rect 247222 711002 247306 711238
rect 247542 711002 282986 711238
rect 283222 711002 283306 711238
rect 283542 711002 318986 711238
rect 319222 711002 319306 711238
rect 319542 711002 354986 711238
rect 355222 711002 355306 711238
rect 355542 711002 390986 711238
rect 391222 711002 391306 711238
rect 391542 711002 426986 711238
rect 427222 711002 427306 711238
rect 427542 711002 462986 711238
rect 463222 711002 463306 711238
rect 463542 711002 498986 711238
rect 499222 711002 499306 711238
rect 499542 711002 534986 711238
rect 535222 711002 535306 711238
rect 535542 711002 570986 711238
rect 571222 711002 571306 711238
rect 571542 711002 592062 711238
rect 592298 711002 592382 711238
rect 592618 711002 592650 711238
rect -8726 710970 592650 711002
rect -7766 710598 591690 710630
rect -7766 710362 -7734 710598
rect -7498 710362 -7414 710598
rect -7178 710362 12986 710598
rect 13222 710362 13306 710598
rect 13542 710362 48986 710598
rect 49222 710362 49306 710598
rect 49542 710362 84986 710598
rect 85222 710362 85306 710598
rect 85542 710362 120986 710598
rect 121222 710362 121306 710598
rect 121542 710362 156986 710598
rect 157222 710362 157306 710598
rect 157542 710362 192986 710598
rect 193222 710362 193306 710598
rect 193542 710362 228986 710598
rect 229222 710362 229306 710598
rect 229542 710362 264986 710598
rect 265222 710362 265306 710598
rect 265542 710362 300986 710598
rect 301222 710362 301306 710598
rect 301542 710362 336986 710598
rect 337222 710362 337306 710598
rect 337542 710362 372986 710598
rect 373222 710362 373306 710598
rect 373542 710362 408986 710598
rect 409222 710362 409306 710598
rect 409542 710362 444986 710598
rect 445222 710362 445306 710598
rect 445542 710362 480986 710598
rect 481222 710362 481306 710598
rect 481542 710362 516986 710598
rect 517222 710362 517306 710598
rect 517542 710362 552986 710598
rect 553222 710362 553306 710598
rect 553542 710362 591102 710598
rect 591338 710362 591422 710598
rect 591658 710362 591690 710598
rect -7766 710278 591690 710362
rect -7766 710042 -7734 710278
rect -7498 710042 -7414 710278
rect -7178 710042 12986 710278
rect 13222 710042 13306 710278
rect 13542 710042 48986 710278
rect 49222 710042 49306 710278
rect 49542 710042 84986 710278
rect 85222 710042 85306 710278
rect 85542 710042 120986 710278
rect 121222 710042 121306 710278
rect 121542 710042 156986 710278
rect 157222 710042 157306 710278
rect 157542 710042 192986 710278
rect 193222 710042 193306 710278
rect 193542 710042 228986 710278
rect 229222 710042 229306 710278
rect 229542 710042 264986 710278
rect 265222 710042 265306 710278
rect 265542 710042 300986 710278
rect 301222 710042 301306 710278
rect 301542 710042 336986 710278
rect 337222 710042 337306 710278
rect 337542 710042 372986 710278
rect 373222 710042 373306 710278
rect 373542 710042 408986 710278
rect 409222 710042 409306 710278
rect 409542 710042 444986 710278
rect 445222 710042 445306 710278
rect 445542 710042 480986 710278
rect 481222 710042 481306 710278
rect 481542 710042 516986 710278
rect 517222 710042 517306 710278
rect 517542 710042 552986 710278
rect 553222 710042 553306 710278
rect 553542 710042 591102 710278
rect 591338 710042 591422 710278
rect 591658 710042 591690 710278
rect -7766 710010 591690 710042
rect -6806 709638 590730 709670
rect -6806 709402 -6774 709638
rect -6538 709402 -6454 709638
rect -6218 709402 27266 709638
rect 27502 709402 27586 709638
rect 27822 709402 63266 709638
rect 63502 709402 63586 709638
rect 63822 709402 99266 709638
rect 99502 709402 99586 709638
rect 99822 709402 135266 709638
rect 135502 709402 135586 709638
rect 135822 709402 171266 709638
rect 171502 709402 171586 709638
rect 171822 709402 207266 709638
rect 207502 709402 207586 709638
rect 207822 709402 243266 709638
rect 243502 709402 243586 709638
rect 243822 709402 279266 709638
rect 279502 709402 279586 709638
rect 279822 709402 315266 709638
rect 315502 709402 315586 709638
rect 315822 709402 351266 709638
rect 351502 709402 351586 709638
rect 351822 709402 387266 709638
rect 387502 709402 387586 709638
rect 387822 709402 423266 709638
rect 423502 709402 423586 709638
rect 423822 709402 459266 709638
rect 459502 709402 459586 709638
rect 459822 709402 495266 709638
rect 495502 709402 495586 709638
rect 495822 709402 531266 709638
rect 531502 709402 531586 709638
rect 531822 709402 567266 709638
rect 567502 709402 567586 709638
rect 567822 709402 590142 709638
rect 590378 709402 590462 709638
rect 590698 709402 590730 709638
rect -6806 709318 590730 709402
rect -6806 709082 -6774 709318
rect -6538 709082 -6454 709318
rect -6218 709082 27266 709318
rect 27502 709082 27586 709318
rect 27822 709082 63266 709318
rect 63502 709082 63586 709318
rect 63822 709082 99266 709318
rect 99502 709082 99586 709318
rect 99822 709082 135266 709318
rect 135502 709082 135586 709318
rect 135822 709082 171266 709318
rect 171502 709082 171586 709318
rect 171822 709082 207266 709318
rect 207502 709082 207586 709318
rect 207822 709082 243266 709318
rect 243502 709082 243586 709318
rect 243822 709082 279266 709318
rect 279502 709082 279586 709318
rect 279822 709082 315266 709318
rect 315502 709082 315586 709318
rect 315822 709082 351266 709318
rect 351502 709082 351586 709318
rect 351822 709082 387266 709318
rect 387502 709082 387586 709318
rect 387822 709082 423266 709318
rect 423502 709082 423586 709318
rect 423822 709082 459266 709318
rect 459502 709082 459586 709318
rect 459822 709082 495266 709318
rect 495502 709082 495586 709318
rect 495822 709082 531266 709318
rect 531502 709082 531586 709318
rect 531822 709082 567266 709318
rect 567502 709082 567586 709318
rect 567822 709082 590142 709318
rect 590378 709082 590462 709318
rect 590698 709082 590730 709318
rect -6806 709050 590730 709082
rect -5846 708678 589770 708710
rect -5846 708442 -5814 708678
rect -5578 708442 -5494 708678
rect -5258 708442 9266 708678
rect 9502 708442 9586 708678
rect 9822 708442 45266 708678
rect 45502 708442 45586 708678
rect 45822 708442 81266 708678
rect 81502 708442 81586 708678
rect 81822 708442 117266 708678
rect 117502 708442 117586 708678
rect 117822 708442 153266 708678
rect 153502 708442 153586 708678
rect 153822 708442 189266 708678
rect 189502 708442 189586 708678
rect 189822 708442 225266 708678
rect 225502 708442 225586 708678
rect 225822 708442 261266 708678
rect 261502 708442 261586 708678
rect 261822 708442 297266 708678
rect 297502 708442 297586 708678
rect 297822 708442 333266 708678
rect 333502 708442 333586 708678
rect 333822 708442 369266 708678
rect 369502 708442 369586 708678
rect 369822 708442 405266 708678
rect 405502 708442 405586 708678
rect 405822 708442 441266 708678
rect 441502 708442 441586 708678
rect 441822 708442 477266 708678
rect 477502 708442 477586 708678
rect 477822 708442 513266 708678
rect 513502 708442 513586 708678
rect 513822 708442 549266 708678
rect 549502 708442 549586 708678
rect 549822 708442 589182 708678
rect 589418 708442 589502 708678
rect 589738 708442 589770 708678
rect -5846 708358 589770 708442
rect -5846 708122 -5814 708358
rect -5578 708122 -5494 708358
rect -5258 708122 9266 708358
rect 9502 708122 9586 708358
rect 9822 708122 45266 708358
rect 45502 708122 45586 708358
rect 45822 708122 81266 708358
rect 81502 708122 81586 708358
rect 81822 708122 117266 708358
rect 117502 708122 117586 708358
rect 117822 708122 153266 708358
rect 153502 708122 153586 708358
rect 153822 708122 189266 708358
rect 189502 708122 189586 708358
rect 189822 708122 225266 708358
rect 225502 708122 225586 708358
rect 225822 708122 261266 708358
rect 261502 708122 261586 708358
rect 261822 708122 297266 708358
rect 297502 708122 297586 708358
rect 297822 708122 333266 708358
rect 333502 708122 333586 708358
rect 333822 708122 369266 708358
rect 369502 708122 369586 708358
rect 369822 708122 405266 708358
rect 405502 708122 405586 708358
rect 405822 708122 441266 708358
rect 441502 708122 441586 708358
rect 441822 708122 477266 708358
rect 477502 708122 477586 708358
rect 477822 708122 513266 708358
rect 513502 708122 513586 708358
rect 513822 708122 549266 708358
rect 549502 708122 549586 708358
rect 549822 708122 589182 708358
rect 589418 708122 589502 708358
rect 589738 708122 589770 708358
rect -5846 708090 589770 708122
rect -4886 707718 588810 707750
rect -4886 707482 -4854 707718
rect -4618 707482 -4534 707718
rect -4298 707482 23546 707718
rect 23782 707482 23866 707718
rect 24102 707482 59546 707718
rect 59782 707482 59866 707718
rect 60102 707482 95546 707718
rect 95782 707482 95866 707718
rect 96102 707482 131546 707718
rect 131782 707482 131866 707718
rect 132102 707482 167546 707718
rect 167782 707482 167866 707718
rect 168102 707482 203546 707718
rect 203782 707482 203866 707718
rect 204102 707482 239546 707718
rect 239782 707482 239866 707718
rect 240102 707482 275546 707718
rect 275782 707482 275866 707718
rect 276102 707482 311546 707718
rect 311782 707482 311866 707718
rect 312102 707482 347546 707718
rect 347782 707482 347866 707718
rect 348102 707482 383546 707718
rect 383782 707482 383866 707718
rect 384102 707482 419546 707718
rect 419782 707482 419866 707718
rect 420102 707482 455546 707718
rect 455782 707482 455866 707718
rect 456102 707482 491546 707718
rect 491782 707482 491866 707718
rect 492102 707482 527546 707718
rect 527782 707482 527866 707718
rect 528102 707482 563546 707718
rect 563782 707482 563866 707718
rect 564102 707482 588222 707718
rect 588458 707482 588542 707718
rect 588778 707482 588810 707718
rect -4886 707398 588810 707482
rect -4886 707162 -4854 707398
rect -4618 707162 -4534 707398
rect -4298 707162 23546 707398
rect 23782 707162 23866 707398
rect 24102 707162 59546 707398
rect 59782 707162 59866 707398
rect 60102 707162 95546 707398
rect 95782 707162 95866 707398
rect 96102 707162 131546 707398
rect 131782 707162 131866 707398
rect 132102 707162 167546 707398
rect 167782 707162 167866 707398
rect 168102 707162 203546 707398
rect 203782 707162 203866 707398
rect 204102 707162 239546 707398
rect 239782 707162 239866 707398
rect 240102 707162 275546 707398
rect 275782 707162 275866 707398
rect 276102 707162 311546 707398
rect 311782 707162 311866 707398
rect 312102 707162 347546 707398
rect 347782 707162 347866 707398
rect 348102 707162 383546 707398
rect 383782 707162 383866 707398
rect 384102 707162 419546 707398
rect 419782 707162 419866 707398
rect 420102 707162 455546 707398
rect 455782 707162 455866 707398
rect 456102 707162 491546 707398
rect 491782 707162 491866 707398
rect 492102 707162 527546 707398
rect 527782 707162 527866 707398
rect 528102 707162 563546 707398
rect 563782 707162 563866 707398
rect 564102 707162 588222 707398
rect 588458 707162 588542 707398
rect 588778 707162 588810 707398
rect -4886 707130 588810 707162
rect -3926 706758 587850 706790
rect -3926 706522 -3894 706758
rect -3658 706522 -3574 706758
rect -3338 706522 5546 706758
rect 5782 706522 5866 706758
rect 6102 706522 41546 706758
rect 41782 706522 41866 706758
rect 42102 706522 77546 706758
rect 77782 706522 77866 706758
rect 78102 706522 113546 706758
rect 113782 706522 113866 706758
rect 114102 706522 149546 706758
rect 149782 706522 149866 706758
rect 150102 706522 185546 706758
rect 185782 706522 185866 706758
rect 186102 706522 221546 706758
rect 221782 706522 221866 706758
rect 222102 706522 257546 706758
rect 257782 706522 257866 706758
rect 258102 706522 293546 706758
rect 293782 706522 293866 706758
rect 294102 706522 329546 706758
rect 329782 706522 329866 706758
rect 330102 706522 365546 706758
rect 365782 706522 365866 706758
rect 366102 706522 401546 706758
rect 401782 706522 401866 706758
rect 402102 706522 437546 706758
rect 437782 706522 437866 706758
rect 438102 706522 473546 706758
rect 473782 706522 473866 706758
rect 474102 706522 509546 706758
rect 509782 706522 509866 706758
rect 510102 706522 545546 706758
rect 545782 706522 545866 706758
rect 546102 706522 581546 706758
rect 581782 706522 581866 706758
rect 582102 706522 587262 706758
rect 587498 706522 587582 706758
rect 587818 706522 587850 706758
rect -3926 706438 587850 706522
rect -3926 706202 -3894 706438
rect -3658 706202 -3574 706438
rect -3338 706202 5546 706438
rect 5782 706202 5866 706438
rect 6102 706202 41546 706438
rect 41782 706202 41866 706438
rect 42102 706202 77546 706438
rect 77782 706202 77866 706438
rect 78102 706202 113546 706438
rect 113782 706202 113866 706438
rect 114102 706202 149546 706438
rect 149782 706202 149866 706438
rect 150102 706202 185546 706438
rect 185782 706202 185866 706438
rect 186102 706202 221546 706438
rect 221782 706202 221866 706438
rect 222102 706202 257546 706438
rect 257782 706202 257866 706438
rect 258102 706202 293546 706438
rect 293782 706202 293866 706438
rect 294102 706202 329546 706438
rect 329782 706202 329866 706438
rect 330102 706202 365546 706438
rect 365782 706202 365866 706438
rect 366102 706202 401546 706438
rect 401782 706202 401866 706438
rect 402102 706202 437546 706438
rect 437782 706202 437866 706438
rect 438102 706202 473546 706438
rect 473782 706202 473866 706438
rect 474102 706202 509546 706438
rect 509782 706202 509866 706438
rect 510102 706202 545546 706438
rect 545782 706202 545866 706438
rect 546102 706202 581546 706438
rect 581782 706202 581866 706438
rect 582102 706202 587262 706438
rect 587498 706202 587582 706438
rect 587818 706202 587850 706438
rect -3926 706170 587850 706202
rect -2966 705798 586890 705830
rect -2966 705562 -2934 705798
rect -2698 705562 -2614 705798
rect -2378 705562 19826 705798
rect 20062 705562 20146 705798
rect 20382 705562 55826 705798
rect 56062 705562 56146 705798
rect 56382 705562 91826 705798
rect 92062 705562 92146 705798
rect 92382 705562 127826 705798
rect 128062 705562 128146 705798
rect 128382 705562 163826 705798
rect 164062 705562 164146 705798
rect 164382 705562 199826 705798
rect 200062 705562 200146 705798
rect 200382 705562 235826 705798
rect 236062 705562 236146 705798
rect 236382 705562 271826 705798
rect 272062 705562 272146 705798
rect 272382 705562 307826 705798
rect 308062 705562 308146 705798
rect 308382 705562 343826 705798
rect 344062 705562 344146 705798
rect 344382 705562 379826 705798
rect 380062 705562 380146 705798
rect 380382 705562 415826 705798
rect 416062 705562 416146 705798
rect 416382 705562 451826 705798
rect 452062 705562 452146 705798
rect 452382 705562 487826 705798
rect 488062 705562 488146 705798
rect 488382 705562 523826 705798
rect 524062 705562 524146 705798
rect 524382 705562 559826 705798
rect 560062 705562 560146 705798
rect 560382 705562 586302 705798
rect 586538 705562 586622 705798
rect 586858 705562 586890 705798
rect -2966 705478 586890 705562
rect -2966 705242 -2934 705478
rect -2698 705242 -2614 705478
rect -2378 705242 19826 705478
rect 20062 705242 20146 705478
rect 20382 705242 55826 705478
rect 56062 705242 56146 705478
rect 56382 705242 91826 705478
rect 92062 705242 92146 705478
rect 92382 705242 127826 705478
rect 128062 705242 128146 705478
rect 128382 705242 163826 705478
rect 164062 705242 164146 705478
rect 164382 705242 199826 705478
rect 200062 705242 200146 705478
rect 200382 705242 235826 705478
rect 236062 705242 236146 705478
rect 236382 705242 271826 705478
rect 272062 705242 272146 705478
rect 272382 705242 307826 705478
rect 308062 705242 308146 705478
rect 308382 705242 343826 705478
rect 344062 705242 344146 705478
rect 344382 705242 379826 705478
rect 380062 705242 380146 705478
rect 380382 705242 415826 705478
rect 416062 705242 416146 705478
rect 416382 705242 451826 705478
rect 452062 705242 452146 705478
rect 452382 705242 487826 705478
rect 488062 705242 488146 705478
rect 488382 705242 523826 705478
rect 524062 705242 524146 705478
rect 524382 705242 559826 705478
rect 560062 705242 560146 705478
rect 560382 705242 586302 705478
rect 586538 705242 586622 705478
rect 586858 705242 586890 705478
rect -2966 705210 586890 705242
rect -2006 704838 585930 704870
rect -2006 704602 -1974 704838
rect -1738 704602 -1654 704838
rect -1418 704602 1826 704838
rect 2062 704602 2146 704838
rect 2382 704602 37826 704838
rect 38062 704602 38146 704838
rect 38382 704602 73826 704838
rect 74062 704602 74146 704838
rect 74382 704602 109826 704838
rect 110062 704602 110146 704838
rect 110382 704602 145826 704838
rect 146062 704602 146146 704838
rect 146382 704602 181826 704838
rect 182062 704602 182146 704838
rect 182382 704602 217826 704838
rect 218062 704602 218146 704838
rect 218382 704602 253826 704838
rect 254062 704602 254146 704838
rect 254382 704602 289826 704838
rect 290062 704602 290146 704838
rect 290382 704602 325826 704838
rect 326062 704602 326146 704838
rect 326382 704602 361826 704838
rect 362062 704602 362146 704838
rect 362382 704602 397826 704838
rect 398062 704602 398146 704838
rect 398382 704602 433826 704838
rect 434062 704602 434146 704838
rect 434382 704602 469826 704838
rect 470062 704602 470146 704838
rect 470382 704602 505826 704838
rect 506062 704602 506146 704838
rect 506382 704602 541826 704838
rect 542062 704602 542146 704838
rect 542382 704602 577826 704838
rect 578062 704602 578146 704838
rect 578382 704602 585342 704838
rect 585578 704602 585662 704838
rect 585898 704602 585930 704838
rect -2006 704518 585930 704602
rect -2006 704282 -1974 704518
rect -1738 704282 -1654 704518
rect -1418 704282 1826 704518
rect 2062 704282 2146 704518
rect 2382 704282 37826 704518
rect 38062 704282 38146 704518
rect 38382 704282 73826 704518
rect 74062 704282 74146 704518
rect 74382 704282 109826 704518
rect 110062 704282 110146 704518
rect 110382 704282 145826 704518
rect 146062 704282 146146 704518
rect 146382 704282 181826 704518
rect 182062 704282 182146 704518
rect 182382 704282 217826 704518
rect 218062 704282 218146 704518
rect 218382 704282 253826 704518
rect 254062 704282 254146 704518
rect 254382 704282 289826 704518
rect 290062 704282 290146 704518
rect 290382 704282 325826 704518
rect 326062 704282 326146 704518
rect 326382 704282 361826 704518
rect 362062 704282 362146 704518
rect 362382 704282 397826 704518
rect 398062 704282 398146 704518
rect 398382 704282 433826 704518
rect 434062 704282 434146 704518
rect 434382 704282 469826 704518
rect 470062 704282 470146 704518
rect 470382 704282 505826 704518
rect 506062 704282 506146 704518
rect 506382 704282 541826 704518
rect 542062 704282 542146 704518
rect 542382 704282 577826 704518
rect 578062 704282 578146 704518
rect 578382 704282 585342 704518
rect 585578 704282 585662 704518
rect 585898 704282 585930 704518
rect -2006 704250 585930 704282
rect -8726 698614 592650 698646
rect -8726 698378 -7734 698614
rect -7498 698378 -7414 698614
rect -7178 698378 591102 698614
rect 591338 698378 591422 698614
rect 591658 698378 592650 698614
rect -8726 698294 592650 698378
rect -8726 698058 -7734 698294
rect -7498 698058 -7414 698294
rect -7178 698058 591102 698294
rect 591338 698058 591422 698294
rect 591658 698058 592650 698294
rect -8726 698026 592650 698058
rect -6806 694894 590730 694926
rect -6806 694658 -5814 694894
rect -5578 694658 -5494 694894
rect -5258 694658 589182 694894
rect 589418 694658 589502 694894
rect 589738 694658 590730 694894
rect -6806 694574 590730 694658
rect -6806 694338 -5814 694574
rect -5578 694338 -5494 694574
rect -5258 694338 589182 694574
rect 589418 694338 589502 694574
rect 589738 694338 590730 694574
rect -6806 694306 590730 694338
rect -4886 691174 588810 691206
rect -4886 690938 -3894 691174
rect -3658 690938 -3574 691174
rect -3338 690938 581546 691174
rect 581782 690938 581866 691174
rect 582102 690938 587262 691174
rect 587498 690938 587582 691174
rect 587818 690938 588810 691174
rect -4886 690854 588810 690938
rect -4886 690618 -3894 690854
rect -3658 690618 -3574 690854
rect -3338 690618 581546 690854
rect 581782 690618 581866 690854
rect 582102 690618 587262 690854
rect 587498 690618 587582 690854
rect 587818 690618 588810 690854
rect -4886 690586 588810 690618
rect -2966 687454 586890 687486
rect -2966 687218 -1974 687454
rect -1738 687218 -1654 687454
rect -1418 687218 8250 687454
rect 8486 687218 38970 687454
rect 39206 687218 69690 687454
rect 69926 687218 100410 687454
rect 100646 687218 131130 687454
rect 131366 687218 161850 687454
rect 162086 687218 192570 687454
rect 192806 687218 223290 687454
rect 223526 687218 254010 687454
rect 254246 687218 284730 687454
rect 284966 687218 315450 687454
rect 315686 687218 346170 687454
rect 346406 687218 376890 687454
rect 377126 687218 407610 687454
rect 407846 687218 438330 687454
rect 438566 687218 469050 687454
rect 469286 687218 499770 687454
rect 500006 687218 530490 687454
rect 530726 687218 561210 687454
rect 561446 687218 577826 687454
rect 578062 687218 578146 687454
rect 578382 687218 585342 687454
rect 585578 687218 585662 687454
rect 585898 687218 586890 687454
rect -2966 687134 586890 687218
rect -2966 686898 -1974 687134
rect -1738 686898 -1654 687134
rect -1418 686898 8250 687134
rect 8486 686898 38970 687134
rect 39206 686898 69690 687134
rect 69926 686898 100410 687134
rect 100646 686898 131130 687134
rect 131366 686898 161850 687134
rect 162086 686898 192570 687134
rect 192806 686898 223290 687134
rect 223526 686898 254010 687134
rect 254246 686898 284730 687134
rect 284966 686898 315450 687134
rect 315686 686898 346170 687134
rect 346406 686898 376890 687134
rect 377126 686898 407610 687134
rect 407846 686898 438330 687134
rect 438566 686898 469050 687134
rect 469286 686898 499770 687134
rect 500006 686898 530490 687134
rect 530726 686898 561210 687134
rect 561446 686898 577826 687134
rect 578062 686898 578146 687134
rect 578382 686898 585342 687134
rect 585578 686898 585662 687134
rect 585898 686898 586890 687134
rect -2966 686866 586890 686898
rect -8726 680614 592650 680646
rect -8726 680378 -8694 680614
rect -8458 680378 -8374 680614
rect -8138 680378 570986 680614
rect 571222 680378 571306 680614
rect 571542 680378 592062 680614
rect 592298 680378 592382 680614
rect 592618 680378 592650 680614
rect -8726 680294 592650 680378
rect -8726 680058 -8694 680294
rect -8458 680058 -8374 680294
rect -8138 680058 570986 680294
rect 571222 680058 571306 680294
rect 571542 680058 592062 680294
rect 592298 680058 592382 680294
rect 592618 680058 592650 680294
rect -8726 680026 592650 680058
rect -6806 676894 590730 676926
rect -6806 676658 -6774 676894
rect -6538 676658 -6454 676894
rect -6218 676658 567266 676894
rect 567502 676658 567586 676894
rect 567822 676658 590142 676894
rect 590378 676658 590462 676894
rect 590698 676658 590730 676894
rect -6806 676574 590730 676658
rect -6806 676338 -6774 676574
rect -6538 676338 -6454 676574
rect -6218 676338 567266 676574
rect 567502 676338 567586 676574
rect 567822 676338 590142 676574
rect 590378 676338 590462 676574
rect 590698 676338 590730 676574
rect -6806 676306 590730 676338
rect -4886 673174 588810 673206
rect -4886 672938 -4854 673174
rect -4618 672938 -4534 673174
rect -4298 672938 588222 673174
rect 588458 672938 588542 673174
rect 588778 672938 588810 673174
rect -4886 672854 588810 672938
rect -4886 672618 -4854 672854
rect -4618 672618 -4534 672854
rect -4298 672618 588222 672854
rect 588458 672618 588542 672854
rect 588778 672618 588810 672854
rect -4886 672586 588810 672618
rect -2966 669454 586890 669486
rect -2966 669218 -2934 669454
rect -2698 669218 -2614 669454
rect -2378 669218 23610 669454
rect 23846 669218 54330 669454
rect 54566 669218 85050 669454
rect 85286 669218 115770 669454
rect 116006 669218 146490 669454
rect 146726 669218 177210 669454
rect 177446 669218 207930 669454
rect 208166 669218 238650 669454
rect 238886 669218 269370 669454
rect 269606 669218 300090 669454
rect 300326 669218 330810 669454
rect 331046 669218 361530 669454
rect 361766 669218 392250 669454
rect 392486 669218 422970 669454
rect 423206 669218 453690 669454
rect 453926 669218 484410 669454
rect 484646 669218 515130 669454
rect 515366 669218 545850 669454
rect 546086 669218 586302 669454
rect 586538 669218 586622 669454
rect 586858 669218 586890 669454
rect -2966 669134 586890 669218
rect -2966 668898 -2934 669134
rect -2698 668898 -2614 669134
rect -2378 668898 23610 669134
rect 23846 668898 54330 669134
rect 54566 668898 85050 669134
rect 85286 668898 115770 669134
rect 116006 668898 146490 669134
rect 146726 668898 177210 669134
rect 177446 668898 207930 669134
rect 208166 668898 238650 669134
rect 238886 668898 269370 669134
rect 269606 668898 300090 669134
rect 300326 668898 330810 669134
rect 331046 668898 361530 669134
rect 361766 668898 392250 669134
rect 392486 668898 422970 669134
rect 423206 668898 453690 669134
rect 453926 668898 484410 669134
rect 484646 668898 515130 669134
rect 515366 668898 545850 669134
rect 546086 668898 586302 669134
rect 586538 668898 586622 669134
rect 586858 668898 586890 669134
rect -2966 668866 586890 668898
rect -8726 662614 592650 662646
rect -8726 662378 -7734 662614
rect -7498 662378 -7414 662614
rect -7178 662378 591102 662614
rect 591338 662378 591422 662614
rect 591658 662378 592650 662614
rect -8726 662294 592650 662378
rect -8726 662058 -7734 662294
rect -7498 662058 -7414 662294
rect -7178 662058 591102 662294
rect 591338 662058 591422 662294
rect 591658 662058 592650 662294
rect -8726 662026 592650 662058
rect -6806 658894 590730 658926
rect -6806 658658 -5814 658894
rect -5578 658658 -5494 658894
rect -5258 658658 589182 658894
rect 589418 658658 589502 658894
rect 589738 658658 590730 658894
rect -6806 658574 590730 658658
rect -6806 658338 -5814 658574
rect -5578 658338 -5494 658574
rect -5258 658338 589182 658574
rect 589418 658338 589502 658574
rect 589738 658338 590730 658574
rect -6806 658306 590730 658338
rect -4886 655174 588810 655206
rect -4886 654938 -3894 655174
rect -3658 654938 -3574 655174
rect -3338 654938 581546 655174
rect 581782 654938 581866 655174
rect 582102 654938 587262 655174
rect 587498 654938 587582 655174
rect 587818 654938 588810 655174
rect -4886 654854 588810 654938
rect -4886 654618 -3894 654854
rect -3658 654618 -3574 654854
rect -3338 654618 581546 654854
rect 581782 654618 581866 654854
rect 582102 654618 587262 654854
rect 587498 654618 587582 654854
rect 587818 654618 588810 654854
rect -4886 654586 588810 654618
rect -2966 651454 586890 651486
rect -2966 651218 -1974 651454
rect -1738 651218 -1654 651454
rect -1418 651218 8250 651454
rect 8486 651218 38970 651454
rect 39206 651218 69690 651454
rect 69926 651218 100410 651454
rect 100646 651218 131130 651454
rect 131366 651218 161850 651454
rect 162086 651218 192570 651454
rect 192806 651218 223290 651454
rect 223526 651218 254010 651454
rect 254246 651218 284730 651454
rect 284966 651218 315450 651454
rect 315686 651218 346170 651454
rect 346406 651218 376890 651454
rect 377126 651218 407610 651454
rect 407846 651218 438330 651454
rect 438566 651218 469050 651454
rect 469286 651218 499770 651454
rect 500006 651218 530490 651454
rect 530726 651218 561210 651454
rect 561446 651218 577826 651454
rect 578062 651218 578146 651454
rect 578382 651218 585342 651454
rect 585578 651218 585662 651454
rect 585898 651218 586890 651454
rect -2966 651134 586890 651218
rect -2966 650898 -1974 651134
rect -1738 650898 -1654 651134
rect -1418 650898 8250 651134
rect 8486 650898 38970 651134
rect 39206 650898 69690 651134
rect 69926 650898 100410 651134
rect 100646 650898 131130 651134
rect 131366 650898 161850 651134
rect 162086 650898 192570 651134
rect 192806 650898 223290 651134
rect 223526 650898 254010 651134
rect 254246 650898 284730 651134
rect 284966 650898 315450 651134
rect 315686 650898 346170 651134
rect 346406 650898 376890 651134
rect 377126 650898 407610 651134
rect 407846 650898 438330 651134
rect 438566 650898 469050 651134
rect 469286 650898 499770 651134
rect 500006 650898 530490 651134
rect 530726 650898 561210 651134
rect 561446 650898 577826 651134
rect 578062 650898 578146 651134
rect 578382 650898 585342 651134
rect 585578 650898 585662 651134
rect 585898 650898 586890 651134
rect -2966 650866 586890 650898
rect -8726 644614 592650 644646
rect -8726 644378 -8694 644614
rect -8458 644378 -8374 644614
rect -8138 644378 570986 644614
rect 571222 644378 571306 644614
rect 571542 644378 592062 644614
rect 592298 644378 592382 644614
rect 592618 644378 592650 644614
rect -8726 644294 592650 644378
rect -8726 644058 -8694 644294
rect -8458 644058 -8374 644294
rect -8138 644058 570986 644294
rect 571222 644058 571306 644294
rect 571542 644058 592062 644294
rect 592298 644058 592382 644294
rect 592618 644058 592650 644294
rect -8726 644026 592650 644058
rect -6806 640894 590730 640926
rect -6806 640658 -6774 640894
rect -6538 640658 -6454 640894
rect -6218 640658 567266 640894
rect 567502 640658 567586 640894
rect 567822 640658 590142 640894
rect 590378 640658 590462 640894
rect 590698 640658 590730 640894
rect -6806 640574 590730 640658
rect -6806 640338 -6774 640574
rect -6538 640338 -6454 640574
rect -6218 640338 567266 640574
rect 567502 640338 567586 640574
rect 567822 640338 590142 640574
rect 590378 640338 590462 640574
rect 590698 640338 590730 640574
rect -6806 640306 590730 640338
rect -4886 637174 588810 637206
rect -4886 636938 -4854 637174
rect -4618 636938 -4534 637174
rect -4298 636938 588222 637174
rect 588458 636938 588542 637174
rect 588778 636938 588810 637174
rect -4886 636854 588810 636938
rect -4886 636618 -4854 636854
rect -4618 636618 -4534 636854
rect -4298 636618 588222 636854
rect 588458 636618 588542 636854
rect 588778 636618 588810 636854
rect -4886 636586 588810 636618
rect -2966 633454 586890 633486
rect -2966 633218 -2934 633454
rect -2698 633218 -2614 633454
rect -2378 633218 23610 633454
rect 23846 633218 54330 633454
rect 54566 633218 85050 633454
rect 85286 633218 115770 633454
rect 116006 633218 146490 633454
rect 146726 633218 177210 633454
rect 177446 633218 207930 633454
rect 208166 633218 238650 633454
rect 238886 633218 269370 633454
rect 269606 633218 300090 633454
rect 300326 633218 330810 633454
rect 331046 633218 361530 633454
rect 361766 633218 392250 633454
rect 392486 633218 422970 633454
rect 423206 633218 453690 633454
rect 453926 633218 484410 633454
rect 484646 633218 515130 633454
rect 515366 633218 545850 633454
rect 546086 633218 586302 633454
rect 586538 633218 586622 633454
rect 586858 633218 586890 633454
rect -2966 633134 586890 633218
rect -2966 632898 -2934 633134
rect -2698 632898 -2614 633134
rect -2378 632898 23610 633134
rect 23846 632898 54330 633134
rect 54566 632898 85050 633134
rect 85286 632898 115770 633134
rect 116006 632898 146490 633134
rect 146726 632898 177210 633134
rect 177446 632898 207930 633134
rect 208166 632898 238650 633134
rect 238886 632898 269370 633134
rect 269606 632898 300090 633134
rect 300326 632898 330810 633134
rect 331046 632898 361530 633134
rect 361766 632898 392250 633134
rect 392486 632898 422970 633134
rect 423206 632898 453690 633134
rect 453926 632898 484410 633134
rect 484646 632898 515130 633134
rect 515366 632898 545850 633134
rect 546086 632898 586302 633134
rect 586538 632898 586622 633134
rect 586858 632898 586890 633134
rect -2966 632866 586890 632898
rect -8726 626614 592650 626646
rect -8726 626378 -7734 626614
rect -7498 626378 -7414 626614
rect -7178 626378 591102 626614
rect 591338 626378 591422 626614
rect 591658 626378 592650 626614
rect -8726 626294 592650 626378
rect -8726 626058 -7734 626294
rect -7498 626058 -7414 626294
rect -7178 626058 591102 626294
rect 591338 626058 591422 626294
rect 591658 626058 592650 626294
rect -8726 626026 592650 626058
rect -6806 622894 590730 622926
rect -6806 622658 -5814 622894
rect -5578 622658 -5494 622894
rect -5258 622658 589182 622894
rect 589418 622658 589502 622894
rect 589738 622658 590730 622894
rect -6806 622574 590730 622658
rect -6806 622338 -5814 622574
rect -5578 622338 -5494 622574
rect -5258 622338 589182 622574
rect 589418 622338 589502 622574
rect 589738 622338 590730 622574
rect -6806 622306 590730 622338
rect -4886 619174 588810 619206
rect -4886 618938 -3894 619174
rect -3658 618938 -3574 619174
rect -3338 618938 581546 619174
rect 581782 618938 581866 619174
rect 582102 618938 587262 619174
rect 587498 618938 587582 619174
rect 587818 618938 588810 619174
rect -4886 618854 588810 618938
rect -4886 618618 -3894 618854
rect -3658 618618 -3574 618854
rect -3338 618618 581546 618854
rect 581782 618618 581866 618854
rect 582102 618618 587262 618854
rect 587498 618618 587582 618854
rect 587818 618618 588810 618854
rect -4886 618586 588810 618618
rect -2966 615454 586890 615486
rect -2966 615218 -1974 615454
rect -1738 615218 -1654 615454
rect -1418 615218 8250 615454
rect 8486 615218 38970 615454
rect 39206 615218 69690 615454
rect 69926 615218 100410 615454
rect 100646 615218 131130 615454
rect 131366 615218 161850 615454
rect 162086 615218 192570 615454
rect 192806 615218 223290 615454
rect 223526 615218 254010 615454
rect 254246 615218 284730 615454
rect 284966 615218 315450 615454
rect 315686 615218 346170 615454
rect 346406 615218 376890 615454
rect 377126 615218 407610 615454
rect 407846 615218 438330 615454
rect 438566 615218 469050 615454
rect 469286 615218 499770 615454
rect 500006 615218 530490 615454
rect 530726 615218 561210 615454
rect 561446 615218 577826 615454
rect 578062 615218 578146 615454
rect 578382 615218 585342 615454
rect 585578 615218 585662 615454
rect 585898 615218 586890 615454
rect -2966 615134 586890 615218
rect -2966 614898 -1974 615134
rect -1738 614898 -1654 615134
rect -1418 614898 8250 615134
rect 8486 614898 38970 615134
rect 39206 614898 69690 615134
rect 69926 614898 100410 615134
rect 100646 614898 131130 615134
rect 131366 614898 161850 615134
rect 162086 614898 192570 615134
rect 192806 614898 223290 615134
rect 223526 614898 254010 615134
rect 254246 614898 284730 615134
rect 284966 614898 315450 615134
rect 315686 614898 346170 615134
rect 346406 614898 376890 615134
rect 377126 614898 407610 615134
rect 407846 614898 438330 615134
rect 438566 614898 469050 615134
rect 469286 614898 499770 615134
rect 500006 614898 530490 615134
rect 530726 614898 561210 615134
rect 561446 614898 577826 615134
rect 578062 614898 578146 615134
rect 578382 614898 585342 615134
rect 585578 614898 585662 615134
rect 585898 614898 586890 615134
rect -2966 614866 586890 614898
rect -8726 608614 592650 608646
rect -8726 608378 -8694 608614
rect -8458 608378 -8374 608614
rect -8138 608378 570986 608614
rect 571222 608378 571306 608614
rect 571542 608378 592062 608614
rect 592298 608378 592382 608614
rect 592618 608378 592650 608614
rect -8726 608294 592650 608378
rect -8726 608058 -8694 608294
rect -8458 608058 -8374 608294
rect -8138 608058 570986 608294
rect 571222 608058 571306 608294
rect 571542 608058 592062 608294
rect 592298 608058 592382 608294
rect 592618 608058 592650 608294
rect -8726 608026 592650 608058
rect -6806 604894 590730 604926
rect -6806 604658 -6774 604894
rect -6538 604658 -6454 604894
rect -6218 604658 567266 604894
rect 567502 604658 567586 604894
rect 567822 604658 590142 604894
rect 590378 604658 590462 604894
rect 590698 604658 590730 604894
rect -6806 604574 590730 604658
rect -6806 604338 -6774 604574
rect -6538 604338 -6454 604574
rect -6218 604338 567266 604574
rect 567502 604338 567586 604574
rect 567822 604338 590142 604574
rect 590378 604338 590462 604574
rect 590698 604338 590730 604574
rect -6806 604306 590730 604338
rect -4886 601174 588810 601206
rect -4886 600938 -4854 601174
rect -4618 600938 -4534 601174
rect -4298 600938 588222 601174
rect 588458 600938 588542 601174
rect 588778 600938 588810 601174
rect -4886 600854 588810 600938
rect -4886 600618 -4854 600854
rect -4618 600618 -4534 600854
rect -4298 600618 588222 600854
rect 588458 600618 588542 600854
rect 588778 600618 588810 600854
rect -4886 600586 588810 600618
rect -2966 597454 586890 597486
rect -2966 597218 -2934 597454
rect -2698 597218 -2614 597454
rect -2378 597218 23610 597454
rect 23846 597218 54330 597454
rect 54566 597218 85050 597454
rect 85286 597218 115770 597454
rect 116006 597218 146490 597454
rect 146726 597218 177210 597454
rect 177446 597218 207930 597454
rect 208166 597218 238650 597454
rect 238886 597218 269370 597454
rect 269606 597218 300090 597454
rect 300326 597218 330810 597454
rect 331046 597218 361530 597454
rect 361766 597218 392250 597454
rect 392486 597218 422970 597454
rect 423206 597218 453690 597454
rect 453926 597218 484410 597454
rect 484646 597218 515130 597454
rect 515366 597218 545850 597454
rect 546086 597218 586302 597454
rect 586538 597218 586622 597454
rect 586858 597218 586890 597454
rect -2966 597134 586890 597218
rect -2966 596898 -2934 597134
rect -2698 596898 -2614 597134
rect -2378 596898 23610 597134
rect 23846 596898 54330 597134
rect 54566 596898 85050 597134
rect 85286 596898 115770 597134
rect 116006 596898 146490 597134
rect 146726 596898 177210 597134
rect 177446 596898 207930 597134
rect 208166 596898 238650 597134
rect 238886 596898 269370 597134
rect 269606 596898 300090 597134
rect 300326 596898 330810 597134
rect 331046 596898 361530 597134
rect 361766 596898 392250 597134
rect 392486 596898 422970 597134
rect 423206 596898 453690 597134
rect 453926 596898 484410 597134
rect 484646 596898 515130 597134
rect 515366 596898 545850 597134
rect 546086 596898 586302 597134
rect 586538 596898 586622 597134
rect 586858 596898 586890 597134
rect -2966 596866 586890 596898
rect -8726 590614 592650 590646
rect -8726 590378 -7734 590614
rect -7498 590378 -7414 590614
rect -7178 590378 591102 590614
rect 591338 590378 591422 590614
rect 591658 590378 592650 590614
rect -8726 590294 592650 590378
rect -8726 590058 -7734 590294
rect -7498 590058 -7414 590294
rect -7178 590058 591102 590294
rect 591338 590058 591422 590294
rect 591658 590058 592650 590294
rect -8726 590026 592650 590058
rect -6806 586894 590730 586926
rect -6806 586658 -5814 586894
rect -5578 586658 -5494 586894
rect -5258 586658 589182 586894
rect 589418 586658 589502 586894
rect 589738 586658 590730 586894
rect -6806 586574 590730 586658
rect -6806 586338 -5814 586574
rect -5578 586338 -5494 586574
rect -5258 586338 589182 586574
rect 589418 586338 589502 586574
rect 589738 586338 590730 586574
rect -6806 586306 590730 586338
rect -4886 583174 588810 583206
rect -4886 582938 -3894 583174
rect -3658 582938 -3574 583174
rect -3338 582938 581546 583174
rect 581782 582938 581866 583174
rect 582102 582938 587262 583174
rect 587498 582938 587582 583174
rect 587818 582938 588810 583174
rect -4886 582854 588810 582938
rect -4886 582618 -3894 582854
rect -3658 582618 -3574 582854
rect -3338 582618 581546 582854
rect 581782 582618 581866 582854
rect 582102 582618 587262 582854
rect 587498 582618 587582 582854
rect 587818 582618 588810 582854
rect -4886 582586 588810 582618
rect -2966 579454 586890 579486
rect -2966 579218 -1974 579454
rect -1738 579218 -1654 579454
rect -1418 579218 8250 579454
rect 8486 579218 38970 579454
rect 39206 579218 69690 579454
rect 69926 579218 100410 579454
rect 100646 579218 131130 579454
rect 131366 579218 161850 579454
rect 162086 579218 192570 579454
rect 192806 579218 223290 579454
rect 223526 579218 254010 579454
rect 254246 579218 284730 579454
rect 284966 579218 315450 579454
rect 315686 579218 346170 579454
rect 346406 579218 376890 579454
rect 377126 579218 407610 579454
rect 407846 579218 438330 579454
rect 438566 579218 469050 579454
rect 469286 579218 499770 579454
rect 500006 579218 530490 579454
rect 530726 579218 561210 579454
rect 561446 579218 577826 579454
rect 578062 579218 578146 579454
rect 578382 579218 585342 579454
rect 585578 579218 585662 579454
rect 585898 579218 586890 579454
rect -2966 579134 586890 579218
rect -2966 578898 -1974 579134
rect -1738 578898 -1654 579134
rect -1418 578898 8250 579134
rect 8486 578898 38970 579134
rect 39206 578898 69690 579134
rect 69926 578898 100410 579134
rect 100646 578898 131130 579134
rect 131366 578898 161850 579134
rect 162086 578898 192570 579134
rect 192806 578898 223290 579134
rect 223526 578898 254010 579134
rect 254246 578898 284730 579134
rect 284966 578898 315450 579134
rect 315686 578898 346170 579134
rect 346406 578898 376890 579134
rect 377126 578898 407610 579134
rect 407846 578898 438330 579134
rect 438566 578898 469050 579134
rect 469286 578898 499770 579134
rect 500006 578898 530490 579134
rect 530726 578898 561210 579134
rect 561446 578898 577826 579134
rect 578062 578898 578146 579134
rect 578382 578898 585342 579134
rect 585578 578898 585662 579134
rect 585898 578898 586890 579134
rect -2966 578866 586890 578898
rect -8726 572614 592650 572646
rect -8726 572378 -8694 572614
rect -8458 572378 -8374 572614
rect -8138 572378 570986 572614
rect 571222 572378 571306 572614
rect 571542 572378 592062 572614
rect 592298 572378 592382 572614
rect 592618 572378 592650 572614
rect -8726 572294 592650 572378
rect -8726 572058 -8694 572294
rect -8458 572058 -8374 572294
rect -8138 572058 570986 572294
rect 571222 572058 571306 572294
rect 571542 572058 592062 572294
rect 592298 572058 592382 572294
rect 592618 572058 592650 572294
rect -8726 572026 592650 572058
rect -6806 568894 590730 568926
rect -6806 568658 -6774 568894
rect -6538 568658 -6454 568894
rect -6218 568658 567266 568894
rect 567502 568658 567586 568894
rect 567822 568658 590142 568894
rect 590378 568658 590462 568894
rect 590698 568658 590730 568894
rect -6806 568574 590730 568658
rect -6806 568338 -6774 568574
rect -6538 568338 -6454 568574
rect -6218 568338 567266 568574
rect 567502 568338 567586 568574
rect 567822 568338 590142 568574
rect 590378 568338 590462 568574
rect 590698 568338 590730 568574
rect -6806 568306 590730 568338
rect -4886 565174 588810 565206
rect -4886 564938 -4854 565174
rect -4618 564938 -4534 565174
rect -4298 564938 588222 565174
rect 588458 564938 588542 565174
rect 588778 564938 588810 565174
rect -4886 564854 588810 564938
rect -4886 564618 -4854 564854
rect -4618 564618 -4534 564854
rect -4298 564618 588222 564854
rect 588458 564618 588542 564854
rect 588778 564618 588810 564854
rect -4886 564586 588810 564618
rect -2966 561454 586890 561486
rect -2966 561218 -2934 561454
rect -2698 561218 -2614 561454
rect -2378 561218 23610 561454
rect 23846 561218 54330 561454
rect 54566 561218 85050 561454
rect 85286 561218 115770 561454
rect 116006 561218 146490 561454
rect 146726 561218 177210 561454
rect 177446 561218 207930 561454
rect 208166 561218 238650 561454
rect 238886 561218 269370 561454
rect 269606 561218 300090 561454
rect 300326 561218 330810 561454
rect 331046 561218 361530 561454
rect 361766 561218 392250 561454
rect 392486 561218 422970 561454
rect 423206 561218 453690 561454
rect 453926 561218 484410 561454
rect 484646 561218 515130 561454
rect 515366 561218 545850 561454
rect 546086 561218 586302 561454
rect 586538 561218 586622 561454
rect 586858 561218 586890 561454
rect -2966 561134 586890 561218
rect -2966 560898 -2934 561134
rect -2698 560898 -2614 561134
rect -2378 560898 23610 561134
rect 23846 560898 54330 561134
rect 54566 560898 85050 561134
rect 85286 560898 115770 561134
rect 116006 560898 146490 561134
rect 146726 560898 177210 561134
rect 177446 560898 207930 561134
rect 208166 560898 238650 561134
rect 238886 560898 269370 561134
rect 269606 560898 300090 561134
rect 300326 560898 330810 561134
rect 331046 560898 361530 561134
rect 361766 560898 392250 561134
rect 392486 560898 422970 561134
rect 423206 560898 453690 561134
rect 453926 560898 484410 561134
rect 484646 560898 515130 561134
rect 515366 560898 545850 561134
rect 546086 560898 586302 561134
rect 586538 560898 586622 561134
rect 586858 560898 586890 561134
rect -2966 560866 586890 560898
rect -8726 554614 592650 554646
rect -8726 554378 -7734 554614
rect -7498 554378 -7414 554614
rect -7178 554378 591102 554614
rect 591338 554378 591422 554614
rect 591658 554378 592650 554614
rect -8726 554294 592650 554378
rect -8726 554058 -7734 554294
rect -7498 554058 -7414 554294
rect -7178 554058 591102 554294
rect 591338 554058 591422 554294
rect 591658 554058 592650 554294
rect -8726 554026 592650 554058
rect -6806 550894 590730 550926
rect -6806 550658 -5814 550894
rect -5578 550658 -5494 550894
rect -5258 550658 589182 550894
rect 589418 550658 589502 550894
rect 589738 550658 590730 550894
rect -6806 550574 590730 550658
rect -6806 550338 -5814 550574
rect -5578 550338 -5494 550574
rect -5258 550338 589182 550574
rect 589418 550338 589502 550574
rect 589738 550338 590730 550574
rect -6806 550306 590730 550338
rect -4886 547174 588810 547206
rect -4886 546938 -3894 547174
rect -3658 546938 -3574 547174
rect -3338 546938 581546 547174
rect 581782 546938 581866 547174
rect 582102 546938 587262 547174
rect 587498 546938 587582 547174
rect 587818 546938 588810 547174
rect -4886 546854 588810 546938
rect -4886 546618 -3894 546854
rect -3658 546618 -3574 546854
rect -3338 546618 581546 546854
rect 581782 546618 581866 546854
rect 582102 546618 587262 546854
rect 587498 546618 587582 546854
rect 587818 546618 588810 546854
rect -4886 546586 588810 546618
rect -2966 543454 586890 543486
rect -2966 543218 -1974 543454
rect -1738 543218 -1654 543454
rect -1418 543218 8250 543454
rect 8486 543218 38970 543454
rect 39206 543218 69690 543454
rect 69926 543218 100410 543454
rect 100646 543218 131130 543454
rect 131366 543218 161850 543454
rect 162086 543218 192570 543454
rect 192806 543218 223290 543454
rect 223526 543218 254010 543454
rect 254246 543218 284730 543454
rect 284966 543218 315450 543454
rect 315686 543218 346170 543454
rect 346406 543218 376890 543454
rect 377126 543218 407610 543454
rect 407846 543218 438330 543454
rect 438566 543218 469050 543454
rect 469286 543218 499770 543454
rect 500006 543218 530490 543454
rect 530726 543218 561210 543454
rect 561446 543218 577826 543454
rect 578062 543218 578146 543454
rect 578382 543218 585342 543454
rect 585578 543218 585662 543454
rect 585898 543218 586890 543454
rect -2966 543134 586890 543218
rect -2966 542898 -1974 543134
rect -1738 542898 -1654 543134
rect -1418 542898 8250 543134
rect 8486 542898 38970 543134
rect 39206 542898 69690 543134
rect 69926 542898 100410 543134
rect 100646 542898 131130 543134
rect 131366 542898 161850 543134
rect 162086 542898 192570 543134
rect 192806 542898 223290 543134
rect 223526 542898 254010 543134
rect 254246 542898 284730 543134
rect 284966 542898 315450 543134
rect 315686 542898 346170 543134
rect 346406 542898 376890 543134
rect 377126 542898 407610 543134
rect 407846 542898 438330 543134
rect 438566 542898 469050 543134
rect 469286 542898 499770 543134
rect 500006 542898 530490 543134
rect 530726 542898 561210 543134
rect 561446 542898 577826 543134
rect 578062 542898 578146 543134
rect 578382 542898 585342 543134
rect 585578 542898 585662 543134
rect 585898 542898 586890 543134
rect -2966 542866 586890 542898
rect -8726 536614 592650 536646
rect -8726 536378 -8694 536614
rect -8458 536378 -8374 536614
rect -8138 536378 570986 536614
rect 571222 536378 571306 536614
rect 571542 536378 592062 536614
rect 592298 536378 592382 536614
rect 592618 536378 592650 536614
rect -8726 536294 592650 536378
rect -8726 536058 -8694 536294
rect -8458 536058 -8374 536294
rect -8138 536058 570986 536294
rect 571222 536058 571306 536294
rect 571542 536058 592062 536294
rect 592298 536058 592382 536294
rect 592618 536058 592650 536294
rect -8726 536026 592650 536058
rect -6806 532894 590730 532926
rect -6806 532658 -6774 532894
rect -6538 532658 -6454 532894
rect -6218 532658 567266 532894
rect 567502 532658 567586 532894
rect 567822 532658 590142 532894
rect 590378 532658 590462 532894
rect 590698 532658 590730 532894
rect -6806 532574 590730 532658
rect -6806 532338 -6774 532574
rect -6538 532338 -6454 532574
rect -6218 532338 567266 532574
rect 567502 532338 567586 532574
rect 567822 532338 590142 532574
rect 590378 532338 590462 532574
rect 590698 532338 590730 532574
rect -6806 532306 590730 532338
rect -4886 529174 588810 529206
rect -4886 528938 -4854 529174
rect -4618 528938 -4534 529174
rect -4298 528938 588222 529174
rect 588458 528938 588542 529174
rect 588778 528938 588810 529174
rect -4886 528854 588810 528938
rect -4886 528618 -4854 528854
rect -4618 528618 -4534 528854
rect -4298 528618 588222 528854
rect 588458 528618 588542 528854
rect 588778 528618 588810 528854
rect -4886 528586 588810 528618
rect -2966 525454 586890 525486
rect -2966 525218 -2934 525454
rect -2698 525218 -2614 525454
rect -2378 525218 23610 525454
rect 23846 525218 54330 525454
rect 54566 525218 85050 525454
rect 85286 525218 115770 525454
rect 116006 525218 146490 525454
rect 146726 525218 177210 525454
rect 177446 525218 207930 525454
rect 208166 525218 238650 525454
rect 238886 525218 269370 525454
rect 269606 525218 300090 525454
rect 300326 525218 330810 525454
rect 331046 525218 361530 525454
rect 361766 525218 392250 525454
rect 392486 525218 422970 525454
rect 423206 525218 453690 525454
rect 453926 525218 484410 525454
rect 484646 525218 515130 525454
rect 515366 525218 545850 525454
rect 546086 525218 586302 525454
rect 586538 525218 586622 525454
rect 586858 525218 586890 525454
rect -2966 525134 586890 525218
rect -2966 524898 -2934 525134
rect -2698 524898 -2614 525134
rect -2378 524898 23610 525134
rect 23846 524898 54330 525134
rect 54566 524898 85050 525134
rect 85286 524898 115770 525134
rect 116006 524898 146490 525134
rect 146726 524898 177210 525134
rect 177446 524898 207930 525134
rect 208166 524898 238650 525134
rect 238886 524898 269370 525134
rect 269606 524898 300090 525134
rect 300326 524898 330810 525134
rect 331046 524898 361530 525134
rect 361766 524898 392250 525134
rect 392486 524898 422970 525134
rect 423206 524898 453690 525134
rect 453926 524898 484410 525134
rect 484646 524898 515130 525134
rect 515366 524898 545850 525134
rect 546086 524898 586302 525134
rect 586538 524898 586622 525134
rect 586858 524898 586890 525134
rect -2966 524866 586890 524898
rect -8726 518614 592650 518646
rect -8726 518378 -7734 518614
rect -7498 518378 -7414 518614
rect -7178 518378 591102 518614
rect 591338 518378 591422 518614
rect 591658 518378 592650 518614
rect -8726 518294 592650 518378
rect -8726 518058 -7734 518294
rect -7498 518058 -7414 518294
rect -7178 518058 591102 518294
rect 591338 518058 591422 518294
rect 591658 518058 592650 518294
rect -8726 518026 592650 518058
rect -6806 514894 590730 514926
rect -6806 514658 -5814 514894
rect -5578 514658 -5494 514894
rect -5258 514658 589182 514894
rect 589418 514658 589502 514894
rect 589738 514658 590730 514894
rect -6806 514574 590730 514658
rect -6806 514338 -5814 514574
rect -5578 514338 -5494 514574
rect -5258 514338 589182 514574
rect 589418 514338 589502 514574
rect 589738 514338 590730 514574
rect -6806 514306 590730 514338
rect -4886 511174 588810 511206
rect -4886 510938 -3894 511174
rect -3658 510938 -3574 511174
rect -3338 510938 581546 511174
rect 581782 510938 581866 511174
rect 582102 510938 587262 511174
rect 587498 510938 587582 511174
rect 587818 510938 588810 511174
rect -4886 510854 588810 510938
rect -4886 510618 -3894 510854
rect -3658 510618 -3574 510854
rect -3338 510618 581546 510854
rect 581782 510618 581866 510854
rect 582102 510618 587262 510854
rect 587498 510618 587582 510854
rect 587818 510618 588810 510854
rect -4886 510586 588810 510618
rect -2966 507454 586890 507486
rect -2966 507218 -1974 507454
rect -1738 507218 -1654 507454
rect -1418 507218 8250 507454
rect 8486 507218 38970 507454
rect 39206 507218 69690 507454
rect 69926 507218 100410 507454
rect 100646 507218 131130 507454
rect 131366 507218 161850 507454
rect 162086 507218 192570 507454
rect 192806 507218 223290 507454
rect 223526 507218 254010 507454
rect 254246 507218 284730 507454
rect 284966 507218 315450 507454
rect 315686 507218 346170 507454
rect 346406 507218 376890 507454
rect 377126 507218 407610 507454
rect 407846 507218 438330 507454
rect 438566 507218 469050 507454
rect 469286 507218 499770 507454
rect 500006 507218 530490 507454
rect 530726 507218 561210 507454
rect 561446 507218 577826 507454
rect 578062 507218 578146 507454
rect 578382 507218 585342 507454
rect 585578 507218 585662 507454
rect 585898 507218 586890 507454
rect -2966 507134 586890 507218
rect -2966 506898 -1974 507134
rect -1738 506898 -1654 507134
rect -1418 506898 8250 507134
rect 8486 506898 38970 507134
rect 39206 506898 69690 507134
rect 69926 506898 100410 507134
rect 100646 506898 131130 507134
rect 131366 506898 161850 507134
rect 162086 506898 192570 507134
rect 192806 506898 223290 507134
rect 223526 506898 254010 507134
rect 254246 506898 284730 507134
rect 284966 506898 315450 507134
rect 315686 506898 346170 507134
rect 346406 506898 376890 507134
rect 377126 506898 407610 507134
rect 407846 506898 438330 507134
rect 438566 506898 469050 507134
rect 469286 506898 499770 507134
rect 500006 506898 530490 507134
rect 530726 506898 561210 507134
rect 561446 506898 577826 507134
rect 578062 506898 578146 507134
rect 578382 506898 585342 507134
rect 585578 506898 585662 507134
rect 585898 506898 586890 507134
rect -2966 506866 586890 506898
rect -8726 500614 592650 500646
rect -8726 500378 -8694 500614
rect -8458 500378 -8374 500614
rect -8138 500378 570986 500614
rect 571222 500378 571306 500614
rect 571542 500378 592062 500614
rect 592298 500378 592382 500614
rect 592618 500378 592650 500614
rect -8726 500294 592650 500378
rect -8726 500058 -8694 500294
rect -8458 500058 -8374 500294
rect -8138 500058 570986 500294
rect 571222 500058 571306 500294
rect 571542 500058 592062 500294
rect 592298 500058 592382 500294
rect 592618 500058 592650 500294
rect -8726 500026 592650 500058
rect -6806 496894 590730 496926
rect -6806 496658 -6774 496894
rect -6538 496658 -6454 496894
rect -6218 496658 567266 496894
rect 567502 496658 567586 496894
rect 567822 496658 590142 496894
rect 590378 496658 590462 496894
rect 590698 496658 590730 496894
rect -6806 496574 590730 496658
rect -6806 496338 -6774 496574
rect -6538 496338 -6454 496574
rect -6218 496338 567266 496574
rect 567502 496338 567586 496574
rect 567822 496338 590142 496574
rect 590378 496338 590462 496574
rect 590698 496338 590730 496574
rect -6806 496306 590730 496338
rect -4886 493174 588810 493206
rect -4886 492938 -4854 493174
rect -4618 492938 -4534 493174
rect -4298 492938 588222 493174
rect 588458 492938 588542 493174
rect 588778 492938 588810 493174
rect -4886 492854 588810 492938
rect -4886 492618 -4854 492854
rect -4618 492618 -4534 492854
rect -4298 492618 588222 492854
rect 588458 492618 588542 492854
rect 588778 492618 588810 492854
rect -4886 492586 588810 492618
rect -2966 489454 586890 489486
rect -2966 489218 -2934 489454
rect -2698 489218 -2614 489454
rect -2378 489218 23610 489454
rect 23846 489218 54330 489454
rect 54566 489218 85050 489454
rect 85286 489218 115770 489454
rect 116006 489218 146490 489454
rect 146726 489218 177210 489454
rect 177446 489218 207930 489454
rect 208166 489218 238650 489454
rect 238886 489218 269370 489454
rect 269606 489218 300090 489454
rect 300326 489218 330810 489454
rect 331046 489218 361530 489454
rect 361766 489218 392250 489454
rect 392486 489218 422970 489454
rect 423206 489218 453690 489454
rect 453926 489218 484410 489454
rect 484646 489218 515130 489454
rect 515366 489218 545850 489454
rect 546086 489218 586302 489454
rect 586538 489218 586622 489454
rect 586858 489218 586890 489454
rect -2966 489134 586890 489218
rect -2966 488898 -2934 489134
rect -2698 488898 -2614 489134
rect -2378 488898 23610 489134
rect 23846 488898 54330 489134
rect 54566 488898 85050 489134
rect 85286 488898 115770 489134
rect 116006 488898 146490 489134
rect 146726 488898 177210 489134
rect 177446 488898 207930 489134
rect 208166 488898 238650 489134
rect 238886 488898 269370 489134
rect 269606 488898 300090 489134
rect 300326 488898 330810 489134
rect 331046 488898 361530 489134
rect 361766 488898 392250 489134
rect 392486 488898 422970 489134
rect 423206 488898 453690 489134
rect 453926 488898 484410 489134
rect 484646 488898 515130 489134
rect 515366 488898 545850 489134
rect 546086 488898 586302 489134
rect 586538 488898 586622 489134
rect 586858 488898 586890 489134
rect -2966 488866 586890 488898
rect -8726 482614 592650 482646
rect -8726 482378 -7734 482614
rect -7498 482378 -7414 482614
rect -7178 482378 591102 482614
rect 591338 482378 591422 482614
rect 591658 482378 592650 482614
rect -8726 482294 592650 482378
rect -8726 482058 -7734 482294
rect -7498 482058 -7414 482294
rect -7178 482058 591102 482294
rect 591338 482058 591422 482294
rect 591658 482058 592650 482294
rect -8726 482026 592650 482058
rect -6806 478894 590730 478926
rect -6806 478658 -5814 478894
rect -5578 478658 -5494 478894
rect -5258 478658 589182 478894
rect 589418 478658 589502 478894
rect 589738 478658 590730 478894
rect -6806 478574 590730 478658
rect -6806 478338 -5814 478574
rect -5578 478338 -5494 478574
rect -5258 478338 589182 478574
rect 589418 478338 589502 478574
rect 589738 478338 590730 478574
rect -6806 478306 590730 478338
rect -4886 475174 588810 475206
rect -4886 474938 -3894 475174
rect -3658 474938 -3574 475174
rect -3338 474938 581546 475174
rect 581782 474938 581866 475174
rect 582102 474938 587262 475174
rect 587498 474938 587582 475174
rect 587818 474938 588810 475174
rect -4886 474854 588810 474938
rect -4886 474618 -3894 474854
rect -3658 474618 -3574 474854
rect -3338 474618 581546 474854
rect 581782 474618 581866 474854
rect 582102 474618 587262 474854
rect 587498 474618 587582 474854
rect 587818 474618 588810 474854
rect -4886 474586 588810 474618
rect -2966 471454 586890 471486
rect -2966 471218 -1974 471454
rect -1738 471218 -1654 471454
rect -1418 471218 8250 471454
rect 8486 471218 38970 471454
rect 39206 471218 69690 471454
rect 69926 471218 100410 471454
rect 100646 471218 131130 471454
rect 131366 471218 161850 471454
rect 162086 471218 192570 471454
rect 192806 471218 223290 471454
rect 223526 471218 254010 471454
rect 254246 471218 284730 471454
rect 284966 471218 315450 471454
rect 315686 471218 346170 471454
rect 346406 471218 376890 471454
rect 377126 471218 407610 471454
rect 407846 471218 438330 471454
rect 438566 471218 469050 471454
rect 469286 471218 499770 471454
rect 500006 471218 530490 471454
rect 530726 471218 561210 471454
rect 561446 471218 577826 471454
rect 578062 471218 578146 471454
rect 578382 471218 585342 471454
rect 585578 471218 585662 471454
rect 585898 471218 586890 471454
rect -2966 471134 586890 471218
rect -2966 470898 -1974 471134
rect -1738 470898 -1654 471134
rect -1418 470898 8250 471134
rect 8486 470898 38970 471134
rect 39206 470898 69690 471134
rect 69926 470898 100410 471134
rect 100646 470898 131130 471134
rect 131366 470898 161850 471134
rect 162086 470898 192570 471134
rect 192806 470898 223290 471134
rect 223526 470898 254010 471134
rect 254246 470898 284730 471134
rect 284966 470898 315450 471134
rect 315686 470898 346170 471134
rect 346406 470898 376890 471134
rect 377126 470898 407610 471134
rect 407846 470898 438330 471134
rect 438566 470898 469050 471134
rect 469286 470898 499770 471134
rect 500006 470898 530490 471134
rect 530726 470898 561210 471134
rect 561446 470898 577826 471134
rect 578062 470898 578146 471134
rect 578382 470898 585342 471134
rect 585578 470898 585662 471134
rect 585898 470898 586890 471134
rect -2966 470866 586890 470898
rect -8726 464614 592650 464646
rect -8726 464378 -8694 464614
rect -8458 464378 -8374 464614
rect -8138 464378 570986 464614
rect 571222 464378 571306 464614
rect 571542 464378 592062 464614
rect 592298 464378 592382 464614
rect 592618 464378 592650 464614
rect -8726 464294 592650 464378
rect -8726 464058 -8694 464294
rect -8458 464058 -8374 464294
rect -8138 464058 570986 464294
rect 571222 464058 571306 464294
rect 571542 464058 592062 464294
rect 592298 464058 592382 464294
rect 592618 464058 592650 464294
rect -8726 464026 592650 464058
rect -6806 460894 590730 460926
rect -6806 460658 -6774 460894
rect -6538 460658 -6454 460894
rect -6218 460658 567266 460894
rect 567502 460658 567586 460894
rect 567822 460658 590142 460894
rect 590378 460658 590462 460894
rect 590698 460658 590730 460894
rect -6806 460574 590730 460658
rect -6806 460338 -6774 460574
rect -6538 460338 -6454 460574
rect -6218 460338 567266 460574
rect 567502 460338 567586 460574
rect 567822 460338 590142 460574
rect 590378 460338 590462 460574
rect 590698 460338 590730 460574
rect -6806 460306 590730 460338
rect -4886 457174 588810 457206
rect -4886 456938 -4854 457174
rect -4618 456938 -4534 457174
rect -4298 456938 588222 457174
rect 588458 456938 588542 457174
rect 588778 456938 588810 457174
rect -4886 456854 588810 456938
rect -4886 456618 -4854 456854
rect -4618 456618 -4534 456854
rect -4298 456618 588222 456854
rect 588458 456618 588542 456854
rect 588778 456618 588810 456854
rect -4886 456586 588810 456618
rect -2966 453454 586890 453486
rect -2966 453218 -2934 453454
rect -2698 453218 -2614 453454
rect -2378 453218 23610 453454
rect 23846 453218 54330 453454
rect 54566 453218 85050 453454
rect 85286 453218 115770 453454
rect 116006 453218 146490 453454
rect 146726 453218 177210 453454
rect 177446 453218 207930 453454
rect 208166 453218 238650 453454
rect 238886 453218 269370 453454
rect 269606 453218 300090 453454
rect 300326 453218 330810 453454
rect 331046 453218 361530 453454
rect 361766 453218 392250 453454
rect 392486 453218 422970 453454
rect 423206 453218 453690 453454
rect 453926 453218 484410 453454
rect 484646 453218 515130 453454
rect 515366 453218 545850 453454
rect 546086 453218 586302 453454
rect 586538 453218 586622 453454
rect 586858 453218 586890 453454
rect -2966 453134 586890 453218
rect -2966 452898 -2934 453134
rect -2698 452898 -2614 453134
rect -2378 452898 23610 453134
rect 23846 452898 54330 453134
rect 54566 452898 85050 453134
rect 85286 452898 115770 453134
rect 116006 452898 146490 453134
rect 146726 452898 177210 453134
rect 177446 452898 207930 453134
rect 208166 452898 238650 453134
rect 238886 452898 269370 453134
rect 269606 452898 300090 453134
rect 300326 452898 330810 453134
rect 331046 452898 361530 453134
rect 361766 452898 392250 453134
rect 392486 452898 422970 453134
rect 423206 452898 453690 453134
rect 453926 452898 484410 453134
rect 484646 452898 515130 453134
rect 515366 452898 545850 453134
rect 546086 452898 586302 453134
rect 586538 452898 586622 453134
rect 586858 452898 586890 453134
rect -2966 452866 586890 452898
rect -8726 446614 592650 446646
rect -8726 446378 -7734 446614
rect -7498 446378 -7414 446614
rect -7178 446378 591102 446614
rect 591338 446378 591422 446614
rect 591658 446378 592650 446614
rect -8726 446294 592650 446378
rect -8726 446058 -7734 446294
rect -7498 446058 -7414 446294
rect -7178 446058 591102 446294
rect 591338 446058 591422 446294
rect 591658 446058 592650 446294
rect -8726 446026 592650 446058
rect -6806 442894 590730 442926
rect -6806 442658 -5814 442894
rect -5578 442658 -5494 442894
rect -5258 442658 589182 442894
rect 589418 442658 589502 442894
rect 589738 442658 590730 442894
rect -6806 442574 590730 442658
rect -6806 442338 -5814 442574
rect -5578 442338 -5494 442574
rect -5258 442338 589182 442574
rect 589418 442338 589502 442574
rect 589738 442338 590730 442574
rect -6806 442306 590730 442338
rect -4886 439174 588810 439206
rect -4886 438938 -3894 439174
rect -3658 438938 -3574 439174
rect -3338 438938 581546 439174
rect 581782 438938 581866 439174
rect 582102 438938 587262 439174
rect 587498 438938 587582 439174
rect 587818 438938 588810 439174
rect -4886 438854 588810 438938
rect -4886 438618 -3894 438854
rect -3658 438618 -3574 438854
rect -3338 438618 581546 438854
rect 581782 438618 581866 438854
rect 582102 438618 587262 438854
rect 587498 438618 587582 438854
rect 587818 438618 588810 438854
rect -4886 438586 588810 438618
rect -2966 435454 586890 435486
rect -2966 435218 -1974 435454
rect -1738 435218 -1654 435454
rect -1418 435218 8250 435454
rect 8486 435218 38970 435454
rect 39206 435218 69690 435454
rect 69926 435218 100410 435454
rect 100646 435218 131130 435454
rect 131366 435218 161850 435454
rect 162086 435218 192570 435454
rect 192806 435218 223290 435454
rect 223526 435218 254010 435454
rect 254246 435218 284730 435454
rect 284966 435218 315450 435454
rect 315686 435218 346170 435454
rect 346406 435218 376890 435454
rect 377126 435218 407610 435454
rect 407846 435218 438330 435454
rect 438566 435218 469050 435454
rect 469286 435218 499770 435454
rect 500006 435218 530490 435454
rect 530726 435218 561210 435454
rect 561446 435218 577826 435454
rect 578062 435218 578146 435454
rect 578382 435218 585342 435454
rect 585578 435218 585662 435454
rect 585898 435218 586890 435454
rect -2966 435134 586890 435218
rect -2966 434898 -1974 435134
rect -1738 434898 -1654 435134
rect -1418 434898 8250 435134
rect 8486 434898 38970 435134
rect 39206 434898 69690 435134
rect 69926 434898 100410 435134
rect 100646 434898 131130 435134
rect 131366 434898 161850 435134
rect 162086 434898 192570 435134
rect 192806 434898 223290 435134
rect 223526 434898 254010 435134
rect 254246 434898 284730 435134
rect 284966 434898 315450 435134
rect 315686 434898 346170 435134
rect 346406 434898 376890 435134
rect 377126 434898 407610 435134
rect 407846 434898 438330 435134
rect 438566 434898 469050 435134
rect 469286 434898 499770 435134
rect 500006 434898 530490 435134
rect 530726 434898 561210 435134
rect 561446 434898 577826 435134
rect 578062 434898 578146 435134
rect 578382 434898 585342 435134
rect 585578 434898 585662 435134
rect 585898 434898 586890 435134
rect -2966 434866 586890 434898
rect -8726 428614 592650 428646
rect -8726 428378 -8694 428614
rect -8458 428378 -8374 428614
rect -8138 428378 570986 428614
rect 571222 428378 571306 428614
rect 571542 428378 592062 428614
rect 592298 428378 592382 428614
rect 592618 428378 592650 428614
rect -8726 428294 592650 428378
rect -8726 428058 -8694 428294
rect -8458 428058 -8374 428294
rect -8138 428058 570986 428294
rect 571222 428058 571306 428294
rect 571542 428058 592062 428294
rect 592298 428058 592382 428294
rect 592618 428058 592650 428294
rect -8726 428026 592650 428058
rect -6806 424894 590730 424926
rect -6806 424658 -6774 424894
rect -6538 424658 -6454 424894
rect -6218 424658 567266 424894
rect 567502 424658 567586 424894
rect 567822 424658 590142 424894
rect 590378 424658 590462 424894
rect 590698 424658 590730 424894
rect -6806 424574 590730 424658
rect -6806 424338 -6774 424574
rect -6538 424338 -6454 424574
rect -6218 424338 567266 424574
rect 567502 424338 567586 424574
rect 567822 424338 590142 424574
rect 590378 424338 590462 424574
rect 590698 424338 590730 424574
rect -6806 424306 590730 424338
rect -4886 421174 588810 421206
rect -4886 420938 -4854 421174
rect -4618 420938 -4534 421174
rect -4298 420938 588222 421174
rect 588458 420938 588542 421174
rect 588778 420938 588810 421174
rect -4886 420854 588810 420938
rect -4886 420618 -4854 420854
rect -4618 420618 -4534 420854
rect -4298 420618 588222 420854
rect 588458 420618 588542 420854
rect 588778 420618 588810 420854
rect -4886 420586 588810 420618
rect -2966 417454 586890 417486
rect -2966 417218 -2934 417454
rect -2698 417218 -2614 417454
rect -2378 417218 23610 417454
rect 23846 417218 54330 417454
rect 54566 417218 85050 417454
rect 85286 417218 115770 417454
rect 116006 417218 146490 417454
rect 146726 417218 177210 417454
rect 177446 417218 207930 417454
rect 208166 417218 238650 417454
rect 238886 417218 269370 417454
rect 269606 417218 300090 417454
rect 300326 417218 330810 417454
rect 331046 417218 361530 417454
rect 361766 417218 392250 417454
rect 392486 417218 422970 417454
rect 423206 417218 453690 417454
rect 453926 417218 484410 417454
rect 484646 417218 515130 417454
rect 515366 417218 545850 417454
rect 546086 417218 586302 417454
rect 586538 417218 586622 417454
rect 586858 417218 586890 417454
rect -2966 417134 586890 417218
rect -2966 416898 -2934 417134
rect -2698 416898 -2614 417134
rect -2378 416898 23610 417134
rect 23846 416898 54330 417134
rect 54566 416898 85050 417134
rect 85286 416898 115770 417134
rect 116006 416898 146490 417134
rect 146726 416898 177210 417134
rect 177446 416898 207930 417134
rect 208166 416898 238650 417134
rect 238886 416898 269370 417134
rect 269606 416898 300090 417134
rect 300326 416898 330810 417134
rect 331046 416898 361530 417134
rect 361766 416898 392250 417134
rect 392486 416898 422970 417134
rect 423206 416898 453690 417134
rect 453926 416898 484410 417134
rect 484646 416898 515130 417134
rect 515366 416898 545850 417134
rect 546086 416898 586302 417134
rect 586538 416898 586622 417134
rect 586858 416898 586890 417134
rect -2966 416866 586890 416898
rect -8726 410614 592650 410646
rect -8726 410378 -7734 410614
rect -7498 410378 -7414 410614
rect -7178 410378 591102 410614
rect 591338 410378 591422 410614
rect 591658 410378 592650 410614
rect -8726 410294 592650 410378
rect -8726 410058 -7734 410294
rect -7498 410058 -7414 410294
rect -7178 410058 591102 410294
rect 591338 410058 591422 410294
rect 591658 410058 592650 410294
rect -8726 410026 592650 410058
rect -6806 406894 590730 406926
rect -6806 406658 -5814 406894
rect -5578 406658 -5494 406894
rect -5258 406658 589182 406894
rect 589418 406658 589502 406894
rect 589738 406658 590730 406894
rect -6806 406574 590730 406658
rect -6806 406338 -5814 406574
rect -5578 406338 -5494 406574
rect -5258 406338 589182 406574
rect 589418 406338 589502 406574
rect 589738 406338 590730 406574
rect -6806 406306 590730 406338
rect -4886 403174 588810 403206
rect -4886 402938 -3894 403174
rect -3658 402938 -3574 403174
rect -3338 402938 581546 403174
rect 581782 402938 581866 403174
rect 582102 402938 587262 403174
rect 587498 402938 587582 403174
rect 587818 402938 588810 403174
rect -4886 402854 588810 402938
rect -4886 402618 -3894 402854
rect -3658 402618 -3574 402854
rect -3338 402618 581546 402854
rect 581782 402618 581866 402854
rect 582102 402618 587262 402854
rect 587498 402618 587582 402854
rect 587818 402618 588810 402854
rect -4886 402586 588810 402618
rect -2966 399454 586890 399486
rect -2966 399218 -1974 399454
rect -1738 399218 -1654 399454
rect -1418 399218 8250 399454
rect 8486 399218 38970 399454
rect 39206 399218 69690 399454
rect 69926 399218 100410 399454
rect 100646 399218 131130 399454
rect 131366 399218 161850 399454
rect 162086 399218 192570 399454
rect 192806 399218 223290 399454
rect 223526 399218 254010 399454
rect 254246 399218 284730 399454
rect 284966 399218 315450 399454
rect 315686 399218 346170 399454
rect 346406 399218 376890 399454
rect 377126 399218 407610 399454
rect 407846 399218 438330 399454
rect 438566 399218 469050 399454
rect 469286 399218 499770 399454
rect 500006 399218 530490 399454
rect 530726 399218 561210 399454
rect 561446 399218 577826 399454
rect 578062 399218 578146 399454
rect 578382 399218 585342 399454
rect 585578 399218 585662 399454
rect 585898 399218 586890 399454
rect -2966 399134 586890 399218
rect -2966 398898 -1974 399134
rect -1738 398898 -1654 399134
rect -1418 398898 8250 399134
rect 8486 398898 38970 399134
rect 39206 398898 69690 399134
rect 69926 398898 100410 399134
rect 100646 398898 131130 399134
rect 131366 398898 161850 399134
rect 162086 398898 192570 399134
rect 192806 398898 223290 399134
rect 223526 398898 254010 399134
rect 254246 398898 284730 399134
rect 284966 398898 315450 399134
rect 315686 398898 346170 399134
rect 346406 398898 376890 399134
rect 377126 398898 407610 399134
rect 407846 398898 438330 399134
rect 438566 398898 469050 399134
rect 469286 398898 499770 399134
rect 500006 398898 530490 399134
rect 530726 398898 561210 399134
rect 561446 398898 577826 399134
rect 578062 398898 578146 399134
rect 578382 398898 585342 399134
rect 585578 398898 585662 399134
rect 585898 398898 586890 399134
rect -2966 398866 586890 398898
rect -8726 392614 592650 392646
rect -8726 392378 -8694 392614
rect -8458 392378 -8374 392614
rect -8138 392378 570986 392614
rect 571222 392378 571306 392614
rect 571542 392378 592062 392614
rect 592298 392378 592382 392614
rect 592618 392378 592650 392614
rect -8726 392294 592650 392378
rect -8726 392058 -8694 392294
rect -8458 392058 -8374 392294
rect -8138 392058 570986 392294
rect 571222 392058 571306 392294
rect 571542 392058 592062 392294
rect 592298 392058 592382 392294
rect 592618 392058 592650 392294
rect -8726 392026 592650 392058
rect -6806 388894 590730 388926
rect -6806 388658 -6774 388894
rect -6538 388658 -6454 388894
rect -6218 388658 567266 388894
rect 567502 388658 567586 388894
rect 567822 388658 590142 388894
rect 590378 388658 590462 388894
rect 590698 388658 590730 388894
rect -6806 388574 590730 388658
rect -6806 388338 -6774 388574
rect -6538 388338 -6454 388574
rect -6218 388338 567266 388574
rect 567502 388338 567586 388574
rect 567822 388338 590142 388574
rect 590378 388338 590462 388574
rect 590698 388338 590730 388574
rect -6806 388306 590730 388338
rect -4886 385174 588810 385206
rect -4886 384938 -4854 385174
rect -4618 384938 -4534 385174
rect -4298 384938 588222 385174
rect 588458 384938 588542 385174
rect 588778 384938 588810 385174
rect -4886 384854 588810 384938
rect -4886 384618 -4854 384854
rect -4618 384618 -4534 384854
rect -4298 384618 588222 384854
rect 588458 384618 588542 384854
rect 588778 384618 588810 384854
rect -4886 384586 588810 384618
rect -2966 381454 586890 381486
rect -2966 381218 -2934 381454
rect -2698 381218 -2614 381454
rect -2378 381218 23610 381454
rect 23846 381218 54330 381454
rect 54566 381218 85050 381454
rect 85286 381218 115770 381454
rect 116006 381218 146490 381454
rect 146726 381218 177210 381454
rect 177446 381218 207930 381454
rect 208166 381218 238650 381454
rect 238886 381218 269370 381454
rect 269606 381218 300090 381454
rect 300326 381218 330810 381454
rect 331046 381218 361530 381454
rect 361766 381218 392250 381454
rect 392486 381218 422970 381454
rect 423206 381218 453690 381454
rect 453926 381218 484410 381454
rect 484646 381218 515130 381454
rect 515366 381218 545850 381454
rect 546086 381218 586302 381454
rect 586538 381218 586622 381454
rect 586858 381218 586890 381454
rect -2966 381134 586890 381218
rect -2966 380898 -2934 381134
rect -2698 380898 -2614 381134
rect -2378 380898 23610 381134
rect 23846 380898 54330 381134
rect 54566 380898 85050 381134
rect 85286 380898 115770 381134
rect 116006 380898 146490 381134
rect 146726 380898 177210 381134
rect 177446 380898 207930 381134
rect 208166 380898 238650 381134
rect 238886 380898 269370 381134
rect 269606 380898 300090 381134
rect 300326 380898 330810 381134
rect 331046 380898 361530 381134
rect 361766 380898 392250 381134
rect 392486 380898 422970 381134
rect 423206 380898 453690 381134
rect 453926 380898 484410 381134
rect 484646 380898 515130 381134
rect 515366 380898 545850 381134
rect 546086 380898 586302 381134
rect 586538 380898 586622 381134
rect 586858 380898 586890 381134
rect -2966 380866 586890 380898
rect -8726 374614 592650 374646
rect -8726 374378 -7734 374614
rect -7498 374378 -7414 374614
rect -7178 374378 591102 374614
rect 591338 374378 591422 374614
rect 591658 374378 592650 374614
rect -8726 374294 592650 374378
rect -8726 374058 -7734 374294
rect -7498 374058 -7414 374294
rect -7178 374058 591102 374294
rect 591338 374058 591422 374294
rect 591658 374058 592650 374294
rect -8726 374026 592650 374058
rect -6806 370894 590730 370926
rect -6806 370658 -5814 370894
rect -5578 370658 -5494 370894
rect -5258 370658 589182 370894
rect 589418 370658 589502 370894
rect 589738 370658 590730 370894
rect -6806 370574 590730 370658
rect -6806 370338 -5814 370574
rect -5578 370338 -5494 370574
rect -5258 370338 589182 370574
rect 589418 370338 589502 370574
rect 589738 370338 590730 370574
rect -6806 370306 590730 370338
rect -4886 367174 588810 367206
rect -4886 366938 -3894 367174
rect -3658 366938 -3574 367174
rect -3338 366938 581546 367174
rect 581782 366938 581866 367174
rect 582102 366938 587262 367174
rect 587498 366938 587582 367174
rect 587818 366938 588810 367174
rect -4886 366854 588810 366938
rect -4886 366618 -3894 366854
rect -3658 366618 -3574 366854
rect -3338 366618 581546 366854
rect 581782 366618 581866 366854
rect 582102 366618 587262 366854
rect 587498 366618 587582 366854
rect 587818 366618 588810 366854
rect -4886 366586 588810 366618
rect -2966 363454 586890 363486
rect -2966 363218 -1974 363454
rect -1738 363218 -1654 363454
rect -1418 363218 8250 363454
rect 8486 363218 38970 363454
rect 39206 363218 69690 363454
rect 69926 363218 100410 363454
rect 100646 363218 131130 363454
rect 131366 363218 161850 363454
rect 162086 363218 192570 363454
rect 192806 363218 223290 363454
rect 223526 363218 254010 363454
rect 254246 363218 284730 363454
rect 284966 363218 315450 363454
rect 315686 363218 346170 363454
rect 346406 363218 376890 363454
rect 377126 363218 407610 363454
rect 407846 363218 438330 363454
rect 438566 363218 469050 363454
rect 469286 363218 499770 363454
rect 500006 363218 530490 363454
rect 530726 363218 561210 363454
rect 561446 363218 577826 363454
rect 578062 363218 578146 363454
rect 578382 363218 585342 363454
rect 585578 363218 585662 363454
rect 585898 363218 586890 363454
rect -2966 363134 586890 363218
rect -2966 362898 -1974 363134
rect -1738 362898 -1654 363134
rect -1418 362898 8250 363134
rect 8486 362898 38970 363134
rect 39206 362898 69690 363134
rect 69926 362898 100410 363134
rect 100646 362898 131130 363134
rect 131366 362898 161850 363134
rect 162086 362898 192570 363134
rect 192806 362898 223290 363134
rect 223526 362898 254010 363134
rect 254246 362898 284730 363134
rect 284966 362898 315450 363134
rect 315686 362898 346170 363134
rect 346406 362898 376890 363134
rect 377126 362898 407610 363134
rect 407846 362898 438330 363134
rect 438566 362898 469050 363134
rect 469286 362898 499770 363134
rect 500006 362898 530490 363134
rect 530726 362898 561210 363134
rect 561446 362898 577826 363134
rect 578062 362898 578146 363134
rect 578382 362898 585342 363134
rect 585578 362898 585662 363134
rect 585898 362898 586890 363134
rect -2966 362866 586890 362898
rect -8726 356614 592650 356646
rect -8726 356378 -8694 356614
rect -8458 356378 -8374 356614
rect -8138 356378 570986 356614
rect 571222 356378 571306 356614
rect 571542 356378 592062 356614
rect 592298 356378 592382 356614
rect 592618 356378 592650 356614
rect -8726 356294 592650 356378
rect -8726 356058 -8694 356294
rect -8458 356058 -8374 356294
rect -8138 356058 570986 356294
rect 571222 356058 571306 356294
rect 571542 356058 592062 356294
rect 592298 356058 592382 356294
rect 592618 356058 592650 356294
rect -8726 356026 592650 356058
rect -6806 352894 590730 352926
rect -6806 352658 -6774 352894
rect -6538 352658 -6454 352894
rect -6218 352658 567266 352894
rect 567502 352658 567586 352894
rect 567822 352658 590142 352894
rect 590378 352658 590462 352894
rect 590698 352658 590730 352894
rect -6806 352574 590730 352658
rect -6806 352338 -6774 352574
rect -6538 352338 -6454 352574
rect -6218 352338 567266 352574
rect 567502 352338 567586 352574
rect 567822 352338 590142 352574
rect 590378 352338 590462 352574
rect 590698 352338 590730 352574
rect -6806 352306 590730 352338
rect -4886 349174 588810 349206
rect -4886 348938 -4854 349174
rect -4618 348938 -4534 349174
rect -4298 348938 588222 349174
rect 588458 348938 588542 349174
rect 588778 348938 588810 349174
rect -4886 348854 588810 348938
rect -4886 348618 -4854 348854
rect -4618 348618 -4534 348854
rect -4298 348618 588222 348854
rect 588458 348618 588542 348854
rect 588778 348618 588810 348854
rect -4886 348586 588810 348618
rect -2966 345454 586890 345486
rect -2966 345218 -2934 345454
rect -2698 345218 -2614 345454
rect -2378 345218 23610 345454
rect 23846 345218 54330 345454
rect 54566 345218 85050 345454
rect 85286 345218 115770 345454
rect 116006 345218 146490 345454
rect 146726 345218 177210 345454
rect 177446 345218 207930 345454
rect 208166 345218 238650 345454
rect 238886 345218 269370 345454
rect 269606 345218 300090 345454
rect 300326 345218 330810 345454
rect 331046 345218 361530 345454
rect 361766 345218 392250 345454
rect 392486 345218 422970 345454
rect 423206 345218 453690 345454
rect 453926 345218 484410 345454
rect 484646 345218 515130 345454
rect 515366 345218 545850 345454
rect 546086 345218 586302 345454
rect 586538 345218 586622 345454
rect 586858 345218 586890 345454
rect -2966 345134 586890 345218
rect -2966 344898 -2934 345134
rect -2698 344898 -2614 345134
rect -2378 344898 23610 345134
rect 23846 344898 54330 345134
rect 54566 344898 85050 345134
rect 85286 344898 115770 345134
rect 116006 344898 146490 345134
rect 146726 344898 177210 345134
rect 177446 344898 207930 345134
rect 208166 344898 238650 345134
rect 238886 344898 269370 345134
rect 269606 344898 300090 345134
rect 300326 344898 330810 345134
rect 331046 344898 361530 345134
rect 361766 344898 392250 345134
rect 392486 344898 422970 345134
rect 423206 344898 453690 345134
rect 453926 344898 484410 345134
rect 484646 344898 515130 345134
rect 515366 344898 545850 345134
rect 546086 344898 586302 345134
rect 586538 344898 586622 345134
rect 586858 344898 586890 345134
rect -2966 344866 586890 344898
rect -8726 338614 592650 338646
rect -8726 338378 -7734 338614
rect -7498 338378 -7414 338614
rect -7178 338378 591102 338614
rect 591338 338378 591422 338614
rect 591658 338378 592650 338614
rect -8726 338294 592650 338378
rect -8726 338058 -7734 338294
rect -7498 338058 -7414 338294
rect -7178 338058 591102 338294
rect 591338 338058 591422 338294
rect 591658 338058 592650 338294
rect -8726 338026 592650 338058
rect -6806 334894 590730 334926
rect -6806 334658 -5814 334894
rect -5578 334658 -5494 334894
rect -5258 334658 589182 334894
rect 589418 334658 589502 334894
rect 589738 334658 590730 334894
rect -6806 334574 590730 334658
rect -6806 334338 -5814 334574
rect -5578 334338 -5494 334574
rect -5258 334338 589182 334574
rect 589418 334338 589502 334574
rect 589738 334338 590730 334574
rect -6806 334306 590730 334338
rect -4886 331174 588810 331206
rect -4886 330938 -3894 331174
rect -3658 330938 -3574 331174
rect -3338 330938 581546 331174
rect 581782 330938 581866 331174
rect 582102 330938 587262 331174
rect 587498 330938 587582 331174
rect 587818 330938 588810 331174
rect -4886 330854 588810 330938
rect -4886 330618 -3894 330854
rect -3658 330618 -3574 330854
rect -3338 330618 581546 330854
rect 581782 330618 581866 330854
rect 582102 330618 587262 330854
rect 587498 330618 587582 330854
rect 587818 330618 588810 330854
rect -4886 330586 588810 330618
rect -2966 327454 586890 327486
rect -2966 327218 -1974 327454
rect -1738 327218 -1654 327454
rect -1418 327218 8250 327454
rect 8486 327218 38970 327454
rect 39206 327218 69690 327454
rect 69926 327218 100410 327454
rect 100646 327218 131130 327454
rect 131366 327218 161850 327454
rect 162086 327218 192570 327454
rect 192806 327218 223290 327454
rect 223526 327218 254010 327454
rect 254246 327218 284730 327454
rect 284966 327218 315450 327454
rect 315686 327218 346170 327454
rect 346406 327218 376890 327454
rect 377126 327218 407610 327454
rect 407846 327218 438330 327454
rect 438566 327218 469050 327454
rect 469286 327218 499770 327454
rect 500006 327218 530490 327454
rect 530726 327218 561210 327454
rect 561446 327218 577826 327454
rect 578062 327218 578146 327454
rect 578382 327218 585342 327454
rect 585578 327218 585662 327454
rect 585898 327218 586890 327454
rect -2966 327134 586890 327218
rect -2966 326898 -1974 327134
rect -1738 326898 -1654 327134
rect -1418 326898 8250 327134
rect 8486 326898 38970 327134
rect 39206 326898 69690 327134
rect 69926 326898 100410 327134
rect 100646 326898 131130 327134
rect 131366 326898 161850 327134
rect 162086 326898 192570 327134
rect 192806 326898 223290 327134
rect 223526 326898 254010 327134
rect 254246 326898 284730 327134
rect 284966 326898 315450 327134
rect 315686 326898 346170 327134
rect 346406 326898 376890 327134
rect 377126 326898 407610 327134
rect 407846 326898 438330 327134
rect 438566 326898 469050 327134
rect 469286 326898 499770 327134
rect 500006 326898 530490 327134
rect 530726 326898 561210 327134
rect 561446 326898 577826 327134
rect 578062 326898 578146 327134
rect 578382 326898 585342 327134
rect 585578 326898 585662 327134
rect 585898 326898 586890 327134
rect -2966 326866 586890 326898
rect -8726 320614 592650 320646
rect -8726 320378 -8694 320614
rect -8458 320378 -8374 320614
rect -8138 320378 570986 320614
rect 571222 320378 571306 320614
rect 571542 320378 592062 320614
rect 592298 320378 592382 320614
rect 592618 320378 592650 320614
rect -8726 320294 592650 320378
rect -8726 320058 -8694 320294
rect -8458 320058 -8374 320294
rect -8138 320058 570986 320294
rect 571222 320058 571306 320294
rect 571542 320058 592062 320294
rect 592298 320058 592382 320294
rect 592618 320058 592650 320294
rect -8726 320026 592650 320058
rect -6806 316894 590730 316926
rect -6806 316658 -6774 316894
rect -6538 316658 -6454 316894
rect -6218 316658 567266 316894
rect 567502 316658 567586 316894
rect 567822 316658 590142 316894
rect 590378 316658 590462 316894
rect 590698 316658 590730 316894
rect -6806 316574 590730 316658
rect -6806 316338 -6774 316574
rect -6538 316338 -6454 316574
rect -6218 316338 567266 316574
rect 567502 316338 567586 316574
rect 567822 316338 590142 316574
rect 590378 316338 590462 316574
rect 590698 316338 590730 316574
rect -6806 316306 590730 316338
rect -4886 313174 588810 313206
rect -4886 312938 -4854 313174
rect -4618 312938 -4534 313174
rect -4298 312938 588222 313174
rect 588458 312938 588542 313174
rect 588778 312938 588810 313174
rect -4886 312854 588810 312938
rect -4886 312618 -4854 312854
rect -4618 312618 -4534 312854
rect -4298 312618 588222 312854
rect 588458 312618 588542 312854
rect 588778 312618 588810 312854
rect -4886 312586 588810 312618
rect -2966 309454 586890 309486
rect -2966 309218 -2934 309454
rect -2698 309218 -2614 309454
rect -2378 309218 23610 309454
rect 23846 309218 54330 309454
rect 54566 309218 85050 309454
rect 85286 309218 115770 309454
rect 116006 309218 146490 309454
rect 146726 309218 177210 309454
rect 177446 309218 207930 309454
rect 208166 309218 238650 309454
rect 238886 309218 269370 309454
rect 269606 309218 300090 309454
rect 300326 309218 330810 309454
rect 331046 309218 361530 309454
rect 361766 309218 392250 309454
rect 392486 309218 422970 309454
rect 423206 309218 453690 309454
rect 453926 309218 484410 309454
rect 484646 309218 515130 309454
rect 515366 309218 545850 309454
rect 546086 309218 586302 309454
rect 586538 309218 586622 309454
rect 586858 309218 586890 309454
rect -2966 309134 586890 309218
rect -2966 308898 -2934 309134
rect -2698 308898 -2614 309134
rect -2378 308898 23610 309134
rect 23846 308898 54330 309134
rect 54566 308898 85050 309134
rect 85286 308898 115770 309134
rect 116006 308898 146490 309134
rect 146726 308898 177210 309134
rect 177446 308898 207930 309134
rect 208166 308898 238650 309134
rect 238886 308898 269370 309134
rect 269606 308898 300090 309134
rect 300326 308898 330810 309134
rect 331046 308898 361530 309134
rect 361766 308898 392250 309134
rect 392486 308898 422970 309134
rect 423206 308898 453690 309134
rect 453926 308898 484410 309134
rect 484646 308898 515130 309134
rect 515366 308898 545850 309134
rect 546086 308898 586302 309134
rect 586538 308898 586622 309134
rect 586858 308898 586890 309134
rect -2966 308866 586890 308898
rect -8726 302614 592650 302646
rect -8726 302378 -7734 302614
rect -7498 302378 -7414 302614
rect -7178 302378 591102 302614
rect 591338 302378 591422 302614
rect 591658 302378 592650 302614
rect -8726 302294 592650 302378
rect -8726 302058 -7734 302294
rect -7498 302058 -7414 302294
rect -7178 302058 591102 302294
rect 591338 302058 591422 302294
rect 591658 302058 592650 302294
rect -8726 302026 592650 302058
rect -6806 298894 590730 298926
rect -6806 298658 -5814 298894
rect -5578 298658 -5494 298894
rect -5258 298658 589182 298894
rect 589418 298658 589502 298894
rect 589738 298658 590730 298894
rect -6806 298574 590730 298658
rect -6806 298338 -5814 298574
rect -5578 298338 -5494 298574
rect -5258 298338 589182 298574
rect 589418 298338 589502 298574
rect 589738 298338 590730 298574
rect -6806 298306 590730 298338
rect -4886 295174 588810 295206
rect -4886 294938 -3894 295174
rect -3658 294938 -3574 295174
rect -3338 294938 581546 295174
rect 581782 294938 581866 295174
rect 582102 294938 587262 295174
rect 587498 294938 587582 295174
rect 587818 294938 588810 295174
rect -4886 294854 588810 294938
rect -4886 294618 -3894 294854
rect -3658 294618 -3574 294854
rect -3338 294618 581546 294854
rect 581782 294618 581866 294854
rect 582102 294618 587262 294854
rect 587498 294618 587582 294854
rect 587818 294618 588810 294854
rect -4886 294586 588810 294618
rect -2966 291454 586890 291486
rect -2966 291218 -1974 291454
rect -1738 291218 -1654 291454
rect -1418 291218 8250 291454
rect 8486 291218 38970 291454
rect 39206 291218 69690 291454
rect 69926 291218 100410 291454
rect 100646 291218 131130 291454
rect 131366 291218 161850 291454
rect 162086 291218 192570 291454
rect 192806 291218 223290 291454
rect 223526 291218 254010 291454
rect 254246 291218 284730 291454
rect 284966 291218 315450 291454
rect 315686 291218 346170 291454
rect 346406 291218 376890 291454
rect 377126 291218 407610 291454
rect 407846 291218 438330 291454
rect 438566 291218 469050 291454
rect 469286 291218 499770 291454
rect 500006 291218 530490 291454
rect 530726 291218 561210 291454
rect 561446 291218 577826 291454
rect 578062 291218 578146 291454
rect 578382 291218 585342 291454
rect 585578 291218 585662 291454
rect 585898 291218 586890 291454
rect -2966 291134 586890 291218
rect -2966 290898 -1974 291134
rect -1738 290898 -1654 291134
rect -1418 290898 8250 291134
rect 8486 290898 38970 291134
rect 39206 290898 69690 291134
rect 69926 290898 100410 291134
rect 100646 290898 131130 291134
rect 131366 290898 161850 291134
rect 162086 290898 192570 291134
rect 192806 290898 223290 291134
rect 223526 290898 254010 291134
rect 254246 290898 284730 291134
rect 284966 290898 315450 291134
rect 315686 290898 346170 291134
rect 346406 290898 376890 291134
rect 377126 290898 407610 291134
rect 407846 290898 438330 291134
rect 438566 290898 469050 291134
rect 469286 290898 499770 291134
rect 500006 290898 530490 291134
rect 530726 290898 561210 291134
rect 561446 290898 577826 291134
rect 578062 290898 578146 291134
rect 578382 290898 585342 291134
rect 585578 290898 585662 291134
rect 585898 290898 586890 291134
rect -2966 290866 586890 290898
rect -8726 284614 592650 284646
rect -8726 284378 -8694 284614
rect -8458 284378 -8374 284614
rect -8138 284378 570986 284614
rect 571222 284378 571306 284614
rect 571542 284378 592062 284614
rect 592298 284378 592382 284614
rect 592618 284378 592650 284614
rect -8726 284294 592650 284378
rect -8726 284058 -8694 284294
rect -8458 284058 -8374 284294
rect -8138 284058 570986 284294
rect 571222 284058 571306 284294
rect 571542 284058 592062 284294
rect 592298 284058 592382 284294
rect 592618 284058 592650 284294
rect -8726 284026 592650 284058
rect -6806 280894 590730 280926
rect -6806 280658 -6774 280894
rect -6538 280658 -6454 280894
rect -6218 280658 567266 280894
rect 567502 280658 567586 280894
rect 567822 280658 590142 280894
rect 590378 280658 590462 280894
rect 590698 280658 590730 280894
rect -6806 280574 590730 280658
rect -6806 280338 -6774 280574
rect -6538 280338 -6454 280574
rect -6218 280338 567266 280574
rect 567502 280338 567586 280574
rect 567822 280338 590142 280574
rect 590378 280338 590462 280574
rect 590698 280338 590730 280574
rect -6806 280306 590730 280338
rect -4886 277174 588810 277206
rect -4886 276938 -4854 277174
rect -4618 276938 -4534 277174
rect -4298 276938 588222 277174
rect 588458 276938 588542 277174
rect 588778 276938 588810 277174
rect -4886 276854 588810 276938
rect -4886 276618 -4854 276854
rect -4618 276618 -4534 276854
rect -4298 276618 588222 276854
rect 588458 276618 588542 276854
rect 588778 276618 588810 276854
rect -4886 276586 588810 276618
rect -2966 273454 586890 273486
rect -2966 273218 -2934 273454
rect -2698 273218 -2614 273454
rect -2378 273218 23610 273454
rect 23846 273218 54330 273454
rect 54566 273218 85050 273454
rect 85286 273218 115770 273454
rect 116006 273218 146490 273454
rect 146726 273218 177210 273454
rect 177446 273218 207930 273454
rect 208166 273218 238650 273454
rect 238886 273218 269370 273454
rect 269606 273218 300090 273454
rect 300326 273218 330810 273454
rect 331046 273218 361530 273454
rect 361766 273218 392250 273454
rect 392486 273218 422970 273454
rect 423206 273218 453690 273454
rect 453926 273218 484410 273454
rect 484646 273218 515130 273454
rect 515366 273218 545850 273454
rect 546086 273218 586302 273454
rect 586538 273218 586622 273454
rect 586858 273218 586890 273454
rect -2966 273134 586890 273218
rect -2966 272898 -2934 273134
rect -2698 272898 -2614 273134
rect -2378 272898 23610 273134
rect 23846 272898 54330 273134
rect 54566 272898 85050 273134
rect 85286 272898 115770 273134
rect 116006 272898 146490 273134
rect 146726 272898 177210 273134
rect 177446 272898 207930 273134
rect 208166 272898 238650 273134
rect 238886 272898 269370 273134
rect 269606 272898 300090 273134
rect 300326 272898 330810 273134
rect 331046 272898 361530 273134
rect 361766 272898 392250 273134
rect 392486 272898 422970 273134
rect 423206 272898 453690 273134
rect 453926 272898 484410 273134
rect 484646 272898 515130 273134
rect 515366 272898 545850 273134
rect 546086 272898 586302 273134
rect 586538 272898 586622 273134
rect 586858 272898 586890 273134
rect -2966 272866 586890 272898
rect -8726 266614 592650 266646
rect -8726 266378 -7734 266614
rect -7498 266378 -7414 266614
rect -7178 266378 591102 266614
rect 591338 266378 591422 266614
rect 591658 266378 592650 266614
rect -8726 266294 592650 266378
rect -8726 266058 -7734 266294
rect -7498 266058 -7414 266294
rect -7178 266058 591102 266294
rect 591338 266058 591422 266294
rect 591658 266058 592650 266294
rect -8726 266026 592650 266058
rect -6806 262894 590730 262926
rect -6806 262658 -5814 262894
rect -5578 262658 -5494 262894
rect -5258 262658 589182 262894
rect 589418 262658 589502 262894
rect 589738 262658 590730 262894
rect -6806 262574 590730 262658
rect -6806 262338 -5814 262574
rect -5578 262338 -5494 262574
rect -5258 262338 589182 262574
rect 589418 262338 589502 262574
rect 589738 262338 590730 262574
rect -6806 262306 590730 262338
rect -4886 259174 588810 259206
rect -4886 258938 -3894 259174
rect -3658 258938 -3574 259174
rect -3338 258938 581546 259174
rect 581782 258938 581866 259174
rect 582102 258938 587262 259174
rect 587498 258938 587582 259174
rect 587818 258938 588810 259174
rect -4886 258854 588810 258938
rect -4886 258618 -3894 258854
rect -3658 258618 -3574 258854
rect -3338 258618 581546 258854
rect 581782 258618 581866 258854
rect 582102 258618 587262 258854
rect 587498 258618 587582 258854
rect 587818 258618 588810 258854
rect -4886 258586 588810 258618
rect -2966 255454 586890 255486
rect -2966 255218 -1974 255454
rect -1738 255218 -1654 255454
rect -1418 255218 8250 255454
rect 8486 255218 38970 255454
rect 39206 255218 69690 255454
rect 69926 255218 100410 255454
rect 100646 255218 131130 255454
rect 131366 255218 161850 255454
rect 162086 255218 192570 255454
rect 192806 255218 223290 255454
rect 223526 255218 254010 255454
rect 254246 255218 284730 255454
rect 284966 255218 315450 255454
rect 315686 255218 346170 255454
rect 346406 255218 376890 255454
rect 377126 255218 407610 255454
rect 407846 255218 438330 255454
rect 438566 255218 469050 255454
rect 469286 255218 499770 255454
rect 500006 255218 530490 255454
rect 530726 255218 561210 255454
rect 561446 255218 577826 255454
rect 578062 255218 578146 255454
rect 578382 255218 585342 255454
rect 585578 255218 585662 255454
rect 585898 255218 586890 255454
rect -2966 255134 586890 255218
rect -2966 254898 -1974 255134
rect -1738 254898 -1654 255134
rect -1418 254898 8250 255134
rect 8486 254898 38970 255134
rect 39206 254898 69690 255134
rect 69926 254898 100410 255134
rect 100646 254898 131130 255134
rect 131366 254898 161850 255134
rect 162086 254898 192570 255134
rect 192806 254898 223290 255134
rect 223526 254898 254010 255134
rect 254246 254898 284730 255134
rect 284966 254898 315450 255134
rect 315686 254898 346170 255134
rect 346406 254898 376890 255134
rect 377126 254898 407610 255134
rect 407846 254898 438330 255134
rect 438566 254898 469050 255134
rect 469286 254898 499770 255134
rect 500006 254898 530490 255134
rect 530726 254898 561210 255134
rect 561446 254898 577826 255134
rect 578062 254898 578146 255134
rect 578382 254898 585342 255134
rect 585578 254898 585662 255134
rect 585898 254898 586890 255134
rect -2966 254866 586890 254898
rect -8726 248614 592650 248646
rect -8726 248378 -8694 248614
rect -8458 248378 -8374 248614
rect -8138 248378 570986 248614
rect 571222 248378 571306 248614
rect 571542 248378 592062 248614
rect 592298 248378 592382 248614
rect 592618 248378 592650 248614
rect -8726 248294 592650 248378
rect -8726 248058 -8694 248294
rect -8458 248058 -8374 248294
rect -8138 248058 570986 248294
rect 571222 248058 571306 248294
rect 571542 248058 592062 248294
rect 592298 248058 592382 248294
rect 592618 248058 592650 248294
rect -8726 248026 592650 248058
rect -6806 244894 590730 244926
rect -6806 244658 -6774 244894
rect -6538 244658 -6454 244894
rect -6218 244658 567266 244894
rect 567502 244658 567586 244894
rect 567822 244658 590142 244894
rect 590378 244658 590462 244894
rect 590698 244658 590730 244894
rect -6806 244574 590730 244658
rect -6806 244338 -6774 244574
rect -6538 244338 -6454 244574
rect -6218 244338 567266 244574
rect 567502 244338 567586 244574
rect 567822 244338 590142 244574
rect 590378 244338 590462 244574
rect 590698 244338 590730 244574
rect -6806 244306 590730 244338
rect -4886 241174 588810 241206
rect -4886 240938 -4854 241174
rect -4618 240938 -4534 241174
rect -4298 240938 588222 241174
rect 588458 240938 588542 241174
rect 588778 240938 588810 241174
rect -4886 240854 588810 240938
rect -4886 240618 -4854 240854
rect -4618 240618 -4534 240854
rect -4298 240618 588222 240854
rect 588458 240618 588542 240854
rect 588778 240618 588810 240854
rect -4886 240586 588810 240618
rect -2966 237454 586890 237486
rect -2966 237218 -2934 237454
rect -2698 237218 -2614 237454
rect -2378 237218 23610 237454
rect 23846 237218 54330 237454
rect 54566 237218 85050 237454
rect 85286 237218 115770 237454
rect 116006 237218 146490 237454
rect 146726 237218 177210 237454
rect 177446 237218 207930 237454
rect 208166 237218 238650 237454
rect 238886 237218 269370 237454
rect 269606 237218 300090 237454
rect 300326 237218 330810 237454
rect 331046 237218 361530 237454
rect 361766 237218 392250 237454
rect 392486 237218 422970 237454
rect 423206 237218 453690 237454
rect 453926 237218 484410 237454
rect 484646 237218 515130 237454
rect 515366 237218 545850 237454
rect 546086 237218 586302 237454
rect 586538 237218 586622 237454
rect 586858 237218 586890 237454
rect -2966 237134 586890 237218
rect -2966 236898 -2934 237134
rect -2698 236898 -2614 237134
rect -2378 236898 23610 237134
rect 23846 236898 54330 237134
rect 54566 236898 85050 237134
rect 85286 236898 115770 237134
rect 116006 236898 146490 237134
rect 146726 236898 177210 237134
rect 177446 236898 207930 237134
rect 208166 236898 238650 237134
rect 238886 236898 269370 237134
rect 269606 236898 300090 237134
rect 300326 236898 330810 237134
rect 331046 236898 361530 237134
rect 361766 236898 392250 237134
rect 392486 236898 422970 237134
rect 423206 236898 453690 237134
rect 453926 236898 484410 237134
rect 484646 236898 515130 237134
rect 515366 236898 545850 237134
rect 546086 236898 586302 237134
rect 586538 236898 586622 237134
rect 586858 236898 586890 237134
rect -2966 236866 586890 236898
rect -8726 230614 592650 230646
rect -8726 230378 -7734 230614
rect -7498 230378 -7414 230614
rect -7178 230378 591102 230614
rect 591338 230378 591422 230614
rect 591658 230378 592650 230614
rect -8726 230294 592650 230378
rect -8726 230058 -7734 230294
rect -7498 230058 -7414 230294
rect -7178 230058 591102 230294
rect 591338 230058 591422 230294
rect 591658 230058 592650 230294
rect -8726 230026 592650 230058
rect -6806 226894 590730 226926
rect -6806 226658 -5814 226894
rect -5578 226658 -5494 226894
rect -5258 226658 589182 226894
rect 589418 226658 589502 226894
rect 589738 226658 590730 226894
rect -6806 226574 590730 226658
rect -6806 226338 -5814 226574
rect -5578 226338 -5494 226574
rect -5258 226338 589182 226574
rect 589418 226338 589502 226574
rect 589738 226338 590730 226574
rect -6806 226306 590730 226338
rect -4886 223174 588810 223206
rect -4886 222938 -3894 223174
rect -3658 222938 -3574 223174
rect -3338 222938 581546 223174
rect 581782 222938 581866 223174
rect 582102 222938 587262 223174
rect 587498 222938 587582 223174
rect 587818 222938 588810 223174
rect -4886 222854 588810 222938
rect -4886 222618 -3894 222854
rect -3658 222618 -3574 222854
rect -3338 222618 581546 222854
rect 581782 222618 581866 222854
rect 582102 222618 587262 222854
rect 587498 222618 587582 222854
rect 587818 222618 588810 222854
rect -4886 222586 588810 222618
rect -2966 219454 586890 219486
rect -2966 219218 -1974 219454
rect -1738 219218 -1654 219454
rect -1418 219218 8250 219454
rect 8486 219218 38970 219454
rect 39206 219218 69690 219454
rect 69926 219218 100410 219454
rect 100646 219218 131130 219454
rect 131366 219218 161850 219454
rect 162086 219218 192570 219454
rect 192806 219218 223290 219454
rect 223526 219218 254010 219454
rect 254246 219218 284730 219454
rect 284966 219218 315450 219454
rect 315686 219218 346170 219454
rect 346406 219218 376890 219454
rect 377126 219218 407610 219454
rect 407846 219218 438330 219454
rect 438566 219218 469050 219454
rect 469286 219218 499770 219454
rect 500006 219218 530490 219454
rect 530726 219218 561210 219454
rect 561446 219218 577826 219454
rect 578062 219218 578146 219454
rect 578382 219218 585342 219454
rect 585578 219218 585662 219454
rect 585898 219218 586890 219454
rect -2966 219134 586890 219218
rect -2966 218898 -1974 219134
rect -1738 218898 -1654 219134
rect -1418 218898 8250 219134
rect 8486 218898 38970 219134
rect 39206 218898 69690 219134
rect 69926 218898 100410 219134
rect 100646 218898 131130 219134
rect 131366 218898 161850 219134
rect 162086 218898 192570 219134
rect 192806 218898 223290 219134
rect 223526 218898 254010 219134
rect 254246 218898 284730 219134
rect 284966 218898 315450 219134
rect 315686 218898 346170 219134
rect 346406 218898 376890 219134
rect 377126 218898 407610 219134
rect 407846 218898 438330 219134
rect 438566 218898 469050 219134
rect 469286 218898 499770 219134
rect 500006 218898 530490 219134
rect 530726 218898 561210 219134
rect 561446 218898 577826 219134
rect 578062 218898 578146 219134
rect 578382 218898 585342 219134
rect 585578 218898 585662 219134
rect 585898 218898 586890 219134
rect -2966 218866 586890 218898
rect -8726 212614 592650 212646
rect -8726 212378 -8694 212614
rect -8458 212378 -8374 212614
rect -8138 212378 570986 212614
rect 571222 212378 571306 212614
rect 571542 212378 592062 212614
rect 592298 212378 592382 212614
rect 592618 212378 592650 212614
rect -8726 212294 592650 212378
rect -8726 212058 -8694 212294
rect -8458 212058 -8374 212294
rect -8138 212058 570986 212294
rect 571222 212058 571306 212294
rect 571542 212058 592062 212294
rect 592298 212058 592382 212294
rect 592618 212058 592650 212294
rect -8726 212026 592650 212058
rect -6806 208894 590730 208926
rect -6806 208658 -6774 208894
rect -6538 208658 -6454 208894
rect -6218 208658 567266 208894
rect 567502 208658 567586 208894
rect 567822 208658 590142 208894
rect 590378 208658 590462 208894
rect 590698 208658 590730 208894
rect -6806 208574 590730 208658
rect -6806 208338 -6774 208574
rect -6538 208338 -6454 208574
rect -6218 208338 567266 208574
rect 567502 208338 567586 208574
rect 567822 208338 590142 208574
rect 590378 208338 590462 208574
rect 590698 208338 590730 208574
rect -6806 208306 590730 208338
rect -4886 205174 588810 205206
rect -4886 204938 -4854 205174
rect -4618 204938 -4534 205174
rect -4298 204938 588222 205174
rect 588458 204938 588542 205174
rect 588778 204938 588810 205174
rect -4886 204854 588810 204938
rect -4886 204618 -4854 204854
rect -4618 204618 -4534 204854
rect -4298 204618 588222 204854
rect 588458 204618 588542 204854
rect 588778 204618 588810 204854
rect -4886 204586 588810 204618
rect -2966 201454 586890 201486
rect -2966 201218 -2934 201454
rect -2698 201218 -2614 201454
rect -2378 201218 23610 201454
rect 23846 201218 54330 201454
rect 54566 201218 85050 201454
rect 85286 201218 115770 201454
rect 116006 201218 146490 201454
rect 146726 201218 177210 201454
rect 177446 201218 207930 201454
rect 208166 201218 238650 201454
rect 238886 201218 269370 201454
rect 269606 201218 300090 201454
rect 300326 201218 330810 201454
rect 331046 201218 361530 201454
rect 361766 201218 392250 201454
rect 392486 201218 422970 201454
rect 423206 201218 453690 201454
rect 453926 201218 484410 201454
rect 484646 201218 515130 201454
rect 515366 201218 545850 201454
rect 546086 201218 586302 201454
rect 586538 201218 586622 201454
rect 586858 201218 586890 201454
rect -2966 201134 586890 201218
rect -2966 200898 -2934 201134
rect -2698 200898 -2614 201134
rect -2378 200898 23610 201134
rect 23846 200898 54330 201134
rect 54566 200898 85050 201134
rect 85286 200898 115770 201134
rect 116006 200898 146490 201134
rect 146726 200898 177210 201134
rect 177446 200898 207930 201134
rect 208166 200898 238650 201134
rect 238886 200898 269370 201134
rect 269606 200898 300090 201134
rect 300326 200898 330810 201134
rect 331046 200898 361530 201134
rect 361766 200898 392250 201134
rect 392486 200898 422970 201134
rect 423206 200898 453690 201134
rect 453926 200898 484410 201134
rect 484646 200898 515130 201134
rect 515366 200898 545850 201134
rect 546086 200898 586302 201134
rect 586538 200898 586622 201134
rect 586858 200898 586890 201134
rect -2966 200866 586890 200898
rect -8726 194614 592650 194646
rect -8726 194378 -7734 194614
rect -7498 194378 -7414 194614
rect -7178 194378 591102 194614
rect 591338 194378 591422 194614
rect 591658 194378 592650 194614
rect -8726 194294 592650 194378
rect -8726 194058 -7734 194294
rect -7498 194058 -7414 194294
rect -7178 194058 591102 194294
rect 591338 194058 591422 194294
rect 591658 194058 592650 194294
rect -8726 194026 592650 194058
rect -6806 190894 590730 190926
rect -6806 190658 -5814 190894
rect -5578 190658 -5494 190894
rect -5258 190658 589182 190894
rect 589418 190658 589502 190894
rect 589738 190658 590730 190894
rect -6806 190574 590730 190658
rect -6806 190338 -5814 190574
rect -5578 190338 -5494 190574
rect -5258 190338 589182 190574
rect 589418 190338 589502 190574
rect 589738 190338 590730 190574
rect -6806 190306 590730 190338
rect -4886 187174 588810 187206
rect -4886 186938 -3894 187174
rect -3658 186938 -3574 187174
rect -3338 186938 581546 187174
rect 581782 186938 581866 187174
rect 582102 186938 587262 187174
rect 587498 186938 587582 187174
rect 587818 186938 588810 187174
rect -4886 186854 588810 186938
rect -4886 186618 -3894 186854
rect -3658 186618 -3574 186854
rect -3338 186618 581546 186854
rect 581782 186618 581866 186854
rect 582102 186618 587262 186854
rect 587498 186618 587582 186854
rect 587818 186618 588810 186854
rect -4886 186586 588810 186618
rect -2966 183454 586890 183486
rect -2966 183218 -1974 183454
rect -1738 183218 -1654 183454
rect -1418 183218 8250 183454
rect 8486 183218 38970 183454
rect 39206 183218 69690 183454
rect 69926 183218 100410 183454
rect 100646 183218 131130 183454
rect 131366 183218 161850 183454
rect 162086 183218 192570 183454
rect 192806 183218 223290 183454
rect 223526 183218 254010 183454
rect 254246 183218 284730 183454
rect 284966 183218 315450 183454
rect 315686 183218 346170 183454
rect 346406 183218 376890 183454
rect 377126 183218 407610 183454
rect 407846 183218 438330 183454
rect 438566 183218 469050 183454
rect 469286 183218 499770 183454
rect 500006 183218 530490 183454
rect 530726 183218 561210 183454
rect 561446 183218 577826 183454
rect 578062 183218 578146 183454
rect 578382 183218 585342 183454
rect 585578 183218 585662 183454
rect 585898 183218 586890 183454
rect -2966 183134 586890 183218
rect -2966 182898 -1974 183134
rect -1738 182898 -1654 183134
rect -1418 182898 8250 183134
rect 8486 182898 38970 183134
rect 39206 182898 69690 183134
rect 69926 182898 100410 183134
rect 100646 182898 131130 183134
rect 131366 182898 161850 183134
rect 162086 182898 192570 183134
rect 192806 182898 223290 183134
rect 223526 182898 254010 183134
rect 254246 182898 284730 183134
rect 284966 182898 315450 183134
rect 315686 182898 346170 183134
rect 346406 182898 376890 183134
rect 377126 182898 407610 183134
rect 407846 182898 438330 183134
rect 438566 182898 469050 183134
rect 469286 182898 499770 183134
rect 500006 182898 530490 183134
rect 530726 182898 561210 183134
rect 561446 182898 577826 183134
rect 578062 182898 578146 183134
rect 578382 182898 585342 183134
rect 585578 182898 585662 183134
rect 585898 182898 586890 183134
rect -2966 182866 586890 182898
rect -8726 176614 592650 176646
rect -8726 176378 -8694 176614
rect -8458 176378 -8374 176614
rect -8138 176378 570986 176614
rect 571222 176378 571306 176614
rect 571542 176378 592062 176614
rect 592298 176378 592382 176614
rect 592618 176378 592650 176614
rect -8726 176294 592650 176378
rect -8726 176058 -8694 176294
rect -8458 176058 -8374 176294
rect -8138 176058 570986 176294
rect 571222 176058 571306 176294
rect 571542 176058 592062 176294
rect 592298 176058 592382 176294
rect 592618 176058 592650 176294
rect -8726 176026 592650 176058
rect -6806 172894 590730 172926
rect -6806 172658 -6774 172894
rect -6538 172658 -6454 172894
rect -6218 172658 567266 172894
rect 567502 172658 567586 172894
rect 567822 172658 590142 172894
rect 590378 172658 590462 172894
rect 590698 172658 590730 172894
rect -6806 172574 590730 172658
rect -6806 172338 -6774 172574
rect -6538 172338 -6454 172574
rect -6218 172338 567266 172574
rect 567502 172338 567586 172574
rect 567822 172338 590142 172574
rect 590378 172338 590462 172574
rect 590698 172338 590730 172574
rect -6806 172306 590730 172338
rect -4886 169174 588810 169206
rect -4886 168938 -4854 169174
rect -4618 168938 -4534 169174
rect -4298 168938 588222 169174
rect 588458 168938 588542 169174
rect 588778 168938 588810 169174
rect -4886 168854 588810 168938
rect -4886 168618 -4854 168854
rect -4618 168618 -4534 168854
rect -4298 168618 588222 168854
rect 588458 168618 588542 168854
rect 588778 168618 588810 168854
rect -4886 168586 588810 168618
rect -2966 165454 586890 165486
rect -2966 165218 -2934 165454
rect -2698 165218 -2614 165454
rect -2378 165218 23610 165454
rect 23846 165218 54330 165454
rect 54566 165218 85050 165454
rect 85286 165218 115770 165454
rect 116006 165218 146490 165454
rect 146726 165218 177210 165454
rect 177446 165218 207930 165454
rect 208166 165218 238650 165454
rect 238886 165218 269370 165454
rect 269606 165218 300090 165454
rect 300326 165218 330810 165454
rect 331046 165218 361530 165454
rect 361766 165218 392250 165454
rect 392486 165218 422970 165454
rect 423206 165218 453690 165454
rect 453926 165218 484410 165454
rect 484646 165218 515130 165454
rect 515366 165218 545850 165454
rect 546086 165218 586302 165454
rect 586538 165218 586622 165454
rect 586858 165218 586890 165454
rect -2966 165134 586890 165218
rect -2966 164898 -2934 165134
rect -2698 164898 -2614 165134
rect -2378 164898 23610 165134
rect 23846 164898 54330 165134
rect 54566 164898 85050 165134
rect 85286 164898 115770 165134
rect 116006 164898 146490 165134
rect 146726 164898 177210 165134
rect 177446 164898 207930 165134
rect 208166 164898 238650 165134
rect 238886 164898 269370 165134
rect 269606 164898 300090 165134
rect 300326 164898 330810 165134
rect 331046 164898 361530 165134
rect 361766 164898 392250 165134
rect 392486 164898 422970 165134
rect 423206 164898 453690 165134
rect 453926 164898 484410 165134
rect 484646 164898 515130 165134
rect 515366 164898 545850 165134
rect 546086 164898 586302 165134
rect 586538 164898 586622 165134
rect 586858 164898 586890 165134
rect -2966 164866 586890 164898
rect -8726 158614 592650 158646
rect -8726 158378 -7734 158614
rect -7498 158378 -7414 158614
rect -7178 158378 591102 158614
rect 591338 158378 591422 158614
rect 591658 158378 592650 158614
rect -8726 158294 592650 158378
rect -8726 158058 -7734 158294
rect -7498 158058 -7414 158294
rect -7178 158058 591102 158294
rect 591338 158058 591422 158294
rect 591658 158058 592650 158294
rect -8726 158026 592650 158058
rect -6806 154894 590730 154926
rect -6806 154658 -5814 154894
rect -5578 154658 -5494 154894
rect -5258 154658 589182 154894
rect 589418 154658 589502 154894
rect 589738 154658 590730 154894
rect -6806 154574 590730 154658
rect -6806 154338 -5814 154574
rect -5578 154338 -5494 154574
rect -5258 154338 589182 154574
rect 589418 154338 589502 154574
rect 589738 154338 590730 154574
rect -6806 154306 590730 154338
rect -4886 151174 588810 151206
rect -4886 150938 -3894 151174
rect -3658 150938 -3574 151174
rect -3338 150938 581546 151174
rect 581782 150938 581866 151174
rect 582102 150938 587262 151174
rect 587498 150938 587582 151174
rect 587818 150938 588810 151174
rect -4886 150854 588810 150938
rect -4886 150618 -3894 150854
rect -3658 150618 -3574 150854
rect -3338 150618 581546 150854
rect 581782 150618 581866 150854
rect 582102 150618 587262 150854
rect 587498 150618 587582 150854
rect 587818 150618 588810 150854
rect -4886 150586 588810 150618
rect -2966 147454 586890 147486
rect -2966 147218 -1974 147454
rect -1738 147218 -1654 147454
rect -1418 147218 8250 147454
rect 8486 147218 38970 147454
rect 39206 147218 69690 147454
rect 69926 147218 100410 147454
rect 100646 147218 131130 147454
rect 131366 147218 161850 147454
rect 162086 147218 192570 147454
rect 192806 147218 223290 147454
rect 223526 147218 254010 147454
rect 254246 147218 284730 147454
rect 284966 147218 315450 147454
rect 315686 147218 346170 147454
rect 346406 147218 376890 147454
rect 377126 147218 407610 147454
rect 407846 147218 438330 147454
rect 438566 147218 469050 147454
rect 469286 147218 499770 147454
rect 500006 147218 530490 147454
rect 530726 147218 561210 147454
rect 561446 147218 577826 147454
rect 578062 147218 578146 147454
rect 578382 147218 585342 147454
rect 585578 147218 585662 147454
rect 585898 147218 586890 147454
rect -2966 147134 586890 147218
rect -2966 146898 -1974 147134
rect -1738 146898 -1654 147134
rect -1418 146898 8250 147134
rect 8486 146898 38970 147134
rect 39206 146898 69690 147134
rect 69926 146898 100410 147134
rect 100646 146898 131130 147134
rect 131366 146898 161850 147134
rect 162086 146898 192570 147134
rect 192806 146898 223290 147134
rect 223526 146898 254010 147134
rect 254246 146898 284730 147134
rect 284966 146898 315450 147134
rect 315686 146898 346170 147134
rect 346406 146898 376890 147134
rect 377126 146898 407610 147134
rect 407846 146898 438330 147134
rect 438566 146898 469050 147134
rect 469286 146898 499770 147134
rect 500006 146898 530490 147134
rect 530726 146898 561210 147134
rect 561446 146898 577826 147134
rect 578062 146898 578146 147134
rect 578382 146898 585342 147134
rect 585578 146898 585662 147134
rect 585898 146898 586890 147134
rect -2966 146866 586890 146898
rect -8726 140614 592650 140646
rect -8726 140378 -8694 140614
rect -8458 140378 -8374 140614
rect -8138 140378 570986 140614
rect 571222 140378 571306 140614
rect 571542 140378 592062 140614
rect 592298 140378 592382 140614
rect 592618 140378 592650 140614
rect -8726 140294 592650 140378
rect -8726 140058 -8694 140294
rect -8458 140058 -8374 140294
rect -8138 140058 570986 140294
rect 571222 140058 571306 140294
rect 571542 140058 592062 140294
rect 592298 140058 592382 140294
rect 592618 140058 592650 140294
rect -8726 140026 592650 140058
rect -6806 136894 590730 136926
rect -6806 136658 -6774 136894
rect -6538 136658 -6454 136894
rect -6218 136658 567266 136894
rect 567502 136658 567586 136894
rect 567822 136658 590142 136894
rect 590378 136658 590462 136894
rect 590698 136658 590730 136894
rect -6806 136574 590730 136658
rect -6806 136338 -6774 136574
rect -6538 136338 -6454 136574
rect -6218 136338 567266 136574
rect 567502 136338 567586 136574
rect 567822 136338 590142 136574
rect 590378 136338 590462 136574
rect 590698 136338 590730 136574
rect -6806 136306 590730 136338
rect -4886 133174 588810 133206
rect -4886 132938 -4854 133174
rect -4618 132938 -4534 133174
rect -4298 132938 588222 133174
rect 588458 132938 588542 133174
rect 588778 132938 588810 133174
rect -4886 132854 588810 132938
rect -4886 132618 -4854 132854
rect -4618 132618 -4534 132854
rect -4298 132618 588222 132854
rect 588458 132618 588542 132854
rect 588778 132618 588810 132854
rect -4886 132586 588810 132618
rect -2966 129454 586890 129486
rect -2966 129218 -2934 129454
rect -2698 129218 -2614 129454
rect -2378 129218 23610 129454
rect 23846 129218 54330 129454
rect 54566 129218 85050 129454
rect 85286 129218 115770 129454
rect 116006 129218 146490 129454
rect 146726 129218 177210 129454
rect 177446 129218 207930 129454
rect 208166 129218 238650 129454
rect 238886 129218 269370 129454
rect 269606 129218 300090 129454
rect 300326 129218 330810 129454
rect 331046 129218 361530 129454
rect 361766 129218 392250 129454
rect 392486 129218 422970 129454
rect 423206 129218 453690 129454
rect 453926 129218 484410 129454
rect 484646 129218 515130 129454
rect 515366 129218 545850 129454
rect 546086 129218 586302 129454
rect 586538 129218 586622 129454
rect 586858 129218 586890 129454
rect -2966 129134 586890 129218
rect -2966 128898 -2934 129134
rect -2698 128898 -2614 129134
rect -2378 128898 23610 129134
rect 23846 128898 54330 129134
rect 54566 128898 85050 129134
rect 85286 128898 115770 129134
rect 116006 128898 146490 129134
rect 146726 128898 177210 129134
rect 177446 128898 207930 129134
rect 208166 128898 238650 129134
rect 238886 128898 269370 129134
rect 269606 128898 300090 129134
rect 300326 128898 330810 129134
rect 331046 128898 361530 129134
rect 361766 128898 392250 129134
rect 392486 128898 422970 129134
rect 423206 128898 453690 129134
rect 453926 128898 484410 129134
rect 484646 128898 515130 129134
rect 515366 128898 545850 129134
rect 546086 128898 586302 129134
rect 586538 128898 586622 129134
rect 586858 128898 586890 129134
rect -2966 128866 586890 128898
rect -8726 122614 592650 122646
rect -8726 122378 -7734 122614
rect -7498 122378 -7414 122614
rect -7178 122378 591102 122614
rect 591338 122378 591422 122614
rect 591658 122378 592650 122614
rect -8726 122294 592650 122378
rect -8726 122058 -7734 122294
rect -7498 122058 -7414 122294
rect -7178 122058 591102 122294
rect 591338 122058 591422 122294
rect 591658 122058 592650 122294
rect -8726 122026 592650 122058
rect -6806 118894 590730 118926
rect -6806 118658 -5814 118894
rect -5578 118658 -5494 118894
rect -5258 118658 589182 118894
rect 589418 118658 589502 118894
rect 589738 118658 590730 118894
rect -6806 118574 590730 118658
rect -6806 118338 -5814 118574
rect -5578 118338 -5494 118574
rect -5258 118338 589182 118574
rect 589418 118338 589502 118574
rect 589738 118338 590730 118574
rect -6806 118306 590730 118338
rect -4886 115174 588810 115206
rect -4886 114938 -3894 115174
rect -3658 114938 -3574 115174
rect -3338 114938 581546 115174
rect 581782 114938 581866 115174
rect 582102 114938 587262 115174
rect 587498 114938 587582 115174
rect 587818 114938 588810 115174
rect -4886 114854 588810 114938
rect -4886 114618 -3894 114854
rect -3658 114618 -3574 114854
rect -3338 114618 581546 114854
rect 581782 114618 581866 114854
rect 582102 114618 587262 114854
rect 587498 114618 587582 114854
rect 587818 114618 588810 114854
rect -4886 114586 588810 114618
rect -2966 111454 586890 111486
rect -2966 111218 -1974 111454
rect -1738 111218 -1654 111454
rect -1418 111218 8250 111454
rect 8486 111218 38970 111454
rect 39206 111218 69690 111454
rect 69926 111218 100410 111454
rect 100646 111218 131130 111454
rect 131366 111218 161850 111454
rect 162086 111218 192570 111454
rect 192806 111218 223290 111454
rect 223526 111218 254010 111454
rect 254246 111218 284730 111454
rect 284966 111218 315450 111454
rect 315686 111218 346170 111454
rect 346406 111218 376890 111454
rect 377126 111218 407610 111454
rect 407846 111218 438330 111454
rect 438566 111218 469050 111454
rect 469286 111218 499770 111454
rect 500006 111218 530490 111454
rect 530726 111218 561210 111454
rect 561446 111218 577826 111454
rect 578062 111218 578146 111454
rect 578382 111218 585342 111454
rect 585578 111218 585662 111454
rect 585898 111218 586890 111454
rect -2966 111134 586890 111218
rect -2966 110898 -1974 111134
rect -1738 110898 -1654 111134
rect -1418 110898 8250 111134
rect 8486 110898 38970 111134
rect 39206 110898 69690 111134
rect 69926 110898 100410 111134
rect 100646 110898 131130 111134
rect 131366 110898 161850 111134
rect 162086 110898 192570 111134
rect 192806 110898 223290 111134
rect 223526 110898 254010 111134
rect 254246 110898 284730 111134
rect 284966 110898 315450 111134
rect 315686 110898 346170 111134
rect 346406 110898 376890 111134
rect 377126 110898 407610 111134
rect 407846 110898 438330 111134
rect 438566 110898 469050 111134
rect 469286 110898 499770 111134
rect 500006 110898 530490 111134
rect 530726 110898 561210 111134
rect 561446 110898 577826 111134
rect 578062 110898 578146 111134
rect 578382 110898 585342 111134
rect 585578 110898 585662 111134
rect 585898 110898 586890 111134
rect -2966 110866 586890 110898
rect -8726 104614 592650 104646
rect -8726 104378 -8694 104614
rect -8458 104378 -8374 104614
rect -8138 104378 570986 104614
rect 571222 104378 571306 104614
rect 571542 104378 592062 104614
rect 592298 104378 592382 104614
rect 592618 104378 592650 104614
rect -8726 104294 592650 104378
rect -8726 104058 -8694 104294
rect -8458 104058 -8374 104294
rect -8138 104058 570986 104294
rect 571222 104058 571306 104294
rect 571542 104058 592062 104294
rect 592298 104058 592382 104294
rect 592618 104058 592650 104294
rect -8726 104026 592650 104058
rect -6806 100894 590730 100926
rect -6806 100658 -6774 100894
rect -6538 100658 -6454 100894
rect -6218 100658 567266 100894
rect 567502 100658 567586 100894
rect 567822 100658 590142 100894
rect 590378 100658 590462 100894
rect 590698 100658 590730 100894
rect -6806 100574 590730 100658
rect -6806 100338 -6774 100574
rect -6538 100338 -6454 100574
rect -6218 100338 567266 100574
rect 567502 100338 567586 100574
rect 567822 100338 590142 100574
rect 590378 100338 590462 100574
rect 590698 100338 590730 100574
rect -6806 100306 590730 100338
rect -4886 97174 588810 97206
rect -4886 96938 -4854 97174
rect -4618 96938 -4534 97174
rect -4298 96938 588222 97174
rect 588458 96938 588542 97174
rect 588778 96938 588810 97174
rect -4886 96854 588810 96938
rect -4886 96618 -4854 96854
rect -4618 96618 -4534 96854
rect -4298 96618 588222 96854
rect 588458 96618 588542 96854
rect 588778 96618 588810 96854
rect -4886 96586 588810 96618
rect -2966 93454 586890 93486
rect -2966 93218 -2934 93454
rect -2698 93218 -2614 93454
rect -2378 93218 23610 93454
rect 23846 93218 54330 93454
rect 54566 93218 85050 93454
rect 85286 93218 115770 93454
rect 116006 93218 146490 93454
rect 146726 93218 177210 93454
rect 177446 93218 207930 93454
rect 208166 93218 238650 93454
rect 238886 93218 269370 93454
rect 269606 93218 300090 93454
rect 300326 93218 330810 93454
rect 331046 93218 361530 93454
rect 361766 93218 392250 93454
rect 392486 93218 422970 93454
rect 423206 93218 453690 93454
rect 453926 93218 484410 93454
rect 484646 93218 515130 93454
rect 515366 93218 545850 93454
rect 546086 93218 586302 93454
rect 586538 93218 586622 93454
rect 586858 93218 586890 93454
rect -2966 93134 586890 93218
rect -2966 92898 -2934 93134
rect -2698 92898 -2614 93134
rect -2378 92898 23610 93134
rect 23846 92898 54330 93134
rect 54566 92898 85050 93134
rect 85286 92898 115770 93134
rect 116006 92898 146490 93134
rect 146726 92898 177210 93134
rect 177446 92898 207930 93134
rect 208166 92898 238650 93134
rect 238886 92898 269370 93134
rect 269606 92898 300090 93134
rect 300326 92898 330810 93134
rect 331046 92898 361530 93134
rect 361766 92898 392250 93134
rect 392486 92898 422970 93134
rect 423206 92898 453690 93134
rect 453926 92898 484410 93134
rect 484646 92898 515130 93134
rect 515366 92898 545850 93134
rect 546086 92898 586302 93134
rect 586538 92898 586622 93134
rect 586858 92898 586890 93134
rect -2966 92866 586890 92898
rect -8726 86614 592650 86646
rect -8726 86378 -7734 86614
rect -7498 86378 -7414 86614
rect -7178 86378 591102 86614
rect 591338 86378 591422 86614
rect 591658 86378 592650 86614
rect -8726 86294 592650 86378
rect -8726 86058 -7734 86294
rect -7498 86058 -7414 86294
rect -7178 86058 591102 86294
rect 591338 86058 591422 86294
rect 591658 86058 592650 86294
rect -8726 86026 592650 86058
rect -6806 82894 590730 82926
rect -6806 82658 -5814 82894
rect -5578 82658 -5494 82894
rect -5258 82658 589182 82894
rect 589418 82658 589502 82894
rect 589738 82658 590730 82894
rect -6806 82574 590730 82658
rect -6806 82338 -5814 82574
rect -5578 82338 -5494 82574
rect -5258 82338 589182 82574
rect 589418 82338 589502 82574
rect 589738 82338 590730 82574
rect -6806 82306 590730 82338
rect -4886 79174 588810 79206
rect -4886 78938 -3894 79174
rect -3658 78938 -3574 79174
rect -3338 78938 581546 79174
rect 581782 78938 581866 79174
rect 582102 78938 587262 79174
rect 587498 78938 587582 79174
rect 587818 78938 588810 79174
rect -4886 78854 588810 78938
rect -4886 78618 -3894 78854
rect -3658 78618 -3574 78854
rect -3338 78618 581546 78854
rect 581782 78618 581866 78854
rect 582102 78618 587262 78854
rect 587498 78618 587582 78854
rect 587818 78618 588810 78854
rect -4886 78586 588810 78618
rect -2966 75454 586890 75486
rect -2966 75218 -1974 75454
rect -1738 75218 -1654 75454
rect -1418 75218 8250 75454
rect 8486 75218 38970 75454
rect 39206 75218 69690 75454
rect 69926 75218 100410 75454
rect 100646 75218 131130 75454
rect 131366 75218 161850 75454
rect 162086 75218 192570 75454
rect 192806 75218 223290 75454
rect 223526 75218 254010 75454
rect 254246 75218 284730 75454
rect 284966 75218 315450 75454
rect 315686 75218 346170 75454
rect 346406 75218 376890 75454
rect 377126 75218 407610 75454
rect 407846 75218 438330 75454
rect 438566 75218 469050 75454
rect 469286 75218 499770 75454
rect 500006 75218 530490 75454
rect 530726 75218 561210 75454
rect 561446 75218 577826 75454
rect 578062 75218 578146 75454
rect 578382 75218 585342 75454
rect 585578 75218 585662 75454
rect 585898 75218 586890 75454
rect -2966 75134 586890 75218
rect -2966 74898 -1974 75134
rect -1738 74898 -1654 75134
rect -1418 74898 8250 75134
rect 8486 74898 38970 75134
rect 39206 74898 69690 75134
rect 69926 74898 100410 75134
rect 100646 74898 131130 75134
rect 131366 74898 161850 75134
rect 162086 74898 192570 75134
rect 192806 74898 223290 75134
rect 223526 74898 254010 75134
rect 254246 74898 284730 75134
rect 284966 74898 315450 75134
rect 315686 74898 346170 75134
rect 346406 74898 376890 75134
rect 377126 74898 407610 75134
rect 407846 74898 438330 75134
rect 438566 74898 469050 75134
rect 469286 74898 499770 75134
rect 500006 74898 530490 75134
rect 530726 74898 561210 75134
rect 561446 74898 577826 75134
rect 578062 74898 578146 75134
rect 578382 74898 585342 75134
rect 585578 74898 585662 75134
rect 585898 74898 586890 75134
rect -2966 74866 586890 74898
rect -8726 68614 592650 68646
rect -8726 68378 -8694 68614
rect -8458 68378 -8374 68614
rect -8138 68378 570986 68614
rect 571222 68378 571306 68614
rect 571542 68378 592062 68614
rect 592298 68378 592382 68614
rect 592618 68378 592650 68614
rect -8726 68294 592650 68378
rect -8726 68058 -8694 68294
rect -8458 68058 -8374 68294
rect -8138 68058 570986 68294
rect 571222 68058 571306 68294
rect 571542 68058 592062 68294
rect 592298 68058 592382 68294
rect 592618 68058 592650 68294
rect -8726 68026 592650 68058
rect -6806 64894 590730 64926
rect -6806 64658 -6774 64894
rect -6538 64658 -6454 64894
rect -6218 64658 567266 64894
rect 567502 64658 567586 64894
rect 567822 64658 590142 64894
rect 590378 64658 590462 64894
rect 590698 64658 590730 64894
rect -6806 64574 590730 64658
rect -6806 64338 -6774 64574
rect -6538 64338 -6454 64574
rect -6218 64338 567266 64574
rect 567502 64338 567586 64574
rect 567822 64338 590142 64574
rect 590378 64338 590462 64574
rect 590698 64338 590730 64574
rect -6806 64306 590730 64338
rect -4886 61174 588810 61206
rect -4886 60938 -4854 61174
rect -4618 60938 -4534 61174
rect -4298 60938 588222 61174
rect 588458 60938 588542 61174
rect 588778 60938 588810 61174
rect -4886 60854 588810 60938
rect -4886 60618 -4854 60854
rect -4618 60618 -4534 60854
rect -4298 60618 588222 60854
rect 588458 60618 588542 60854
rect 588778 60618 588810 60854
rect -4886 60586 588810 60618
rect -2966 57454 586890 57486
rect -2966 57218 -2934 57454
rect -2698 57218 -2614 57454
rect -2378 57218 23610 57454
rect 23846 57218 54330 57454
rect 54566 57218 85050 57454
rect 85286 57218 115770 57454
rect 116006 57218 146490 57454
rect 146726 57218 177210 57454
rect 177446 57218 207930 57454
rect 208166 57218 238650 57454
rect 238886 57218 269370 57454
rect 269606 57218 300090 57454
rect 300326 57218 330810 57454
rect 331046 57218 361530 57454
rect 361766 57218 392250 57454
rect 392486 57218 422970 57454
rect 423206 57218 453690 57454
rect 453926 57218 484410 57454
rect 484646 57218 515130 57454
rect 515366 57218 545850 57454
rect 546086 57218 586302 57454
rect 586538 57218 586622 57454
rect 586858 57218 586890 57454
rect -2966 57134 586890 57218
rect -2966 56898 -2934 57134
rect -2698 56898 -2614 57134
rect -2378 56898 23610 57134
rect 23846 56898 54330 57134
rect 54566 56898 85050 57134
rect 85286 56898 115770 57134
rect 116006 56898 146490 57134
rect 146726 56898 177210 57134
rect 177446 56898 207930 57134
rect 208166 56898 238650 57134
rect 238886 56898 269370 57134
rect 269606 56898 300090 57134
rect 300326 56898 330810 57134
rect 331046 56898 361530 57134
rect 361766 56898 392250 57134
rect 392486 56898 422970 57134
rect 423206 56898 453690 57134
rect 453926 56898 484410 57134
rect 484646 56898 515130 57134
rect 515366 56898 545850 57134
rect 546086 56898 586302 57134
rect 586538 56898 586622 57134
rect 586858 56898 586890 57134
rect -2966 56866 586890 56898
rect -8726 50614 592650 50646
rect -8726 50378 -7734 50614
rect -7498 50378 -7414 50614
rect -7178 50378 591102 50614
rect 591338 50378 591422 50614
rect 591658 50378 592650 50614
rect -8726 50294 592650 50378
rect -8726 50058 -7734 50294
rect -7498 50058 -7414 50294
rect -7178 50058 591102 50294
rect 591338 50058 591422 50294
rect 591658 50058 592650 50294
rect -8726 50026 592650 50058
rect -6806 46894 590730 46926
rect -6806 46658 -5814 46894
rect -5578 46658 -5494 46894
rect -5258 46658 589182 46894
rect 589418 46658 589502 46894
rect 589738 46658 590730 46894
rect -6806 46574 590730 46658
rect -6806 46338 -5814 46574
rect -5578 46338 -5494 46574
rect -5258 46338 589182 46574
rect 589418 46338 589502 46574
rect 589738 46338 590730 46574
rect -6806 46306 590730 46338
rect -4886 43174 588810 43206
rect -4886 42938 -3894 43174
rect -3658 42938 -3574 43174
rect -3338 42938 581546 43174
rect 581782 42938 581866 43174
rect 582102 42938 587262 43174
rect 587498 42938 587582 43174
rect 587818 42938 588810 43174
rect -4886 42854 588810 42938
rect -4886 42618 -3894 42854
rect -3658 42618 -3574 42854
rect -3338 42618 581546 42854
rect 581782 42618 581866 42854
rect 582102 42618 587262 42854
rect 587498 42618 587582 42854
rect 587818 42618 588810 42854
rect -4886 42586 588810 42618
rect -2966 39454 586890 39486
rect -2966 39218 -1974 39454
rect -1738 39218 -1654 39454
rect -1418 39218 8250 39454
rect 8486 39218 38970 39454
rect 39206 39218 69690 39454
rect 69926 39218 100410 39454
rect 100646 39218 131130 39454
rect 131366 39218 161850 39454
rect 162086 39218 192570 39454
rect 192806 39218 223290 39454
rect 223526 39218 254010 39454
rect 254246 39218 284730 39454
rect 284966 39218 315450 39454
rect 315686 39218 346170 39454
rect 346406 39218 376890 39454
rect 377126 39218 407610 39454
rect 407846 39218 438330 39454
rect 438566 39218 469050 39454
rect 469286 39218 499770 39454
rect 500006 39218 530490 39454
rect 530726 39218 561210 39454
rect 561446 39218 577826 39454
rect 578062 39218 578146 39454
rect 578382 39218 585342 39454
rect 585578 39218 585662 39454
rect 585898 39218 586890 39454
rect -2966 39134 586890 39218
rect -2966 38898 -1974 39134
rect -1738 38898 -1654 39134
rect -1418 38898 8250 39134
rect 8486 38898 38970 39134
rect 39206 38898 69690 39134
rect 69926 38898 100410 39134
rect 100646 38898 131130 39134
rect 131366 38898 161850 39134
rect 162086 38898 192570 39134
rect 192806 38898 223290 39134
rect 223526 38898 254010 39134
rect 254246 38898 284730 39134
rect 284966 38898 315450 39134
rect 315686 38898 346170 39134
rect 346406 38898 376890 39134
rect 377126 38898 407610 39134
rect 407846 38898 438330 39134
rect 438566 38898 469050 39134
rect 469286 38898 499770 39134
rect 500006 38898 530490 39134
rect 530726 38898 561210 39134
rect 561446 38898 577826 39134
rect 578062 38898 578146 39134
rect 578382 38898 585342 39134
rect 585578 38898 585662 39134
rect 585898 38898 586890 39134
rect -2966 38866 586890 38898
rect -8726 32614 592650 32646
rect -8726 32378 -8694 32614
rect -8458 32378 -8374 32614
rect -8138 32378 570986 32614
rect 571222 32378 571306 32614
rect 571542 32378 592062 32614
rect 592298 32378 592382 32614
rect 592618 32378 592650 32614
rect -8726 32294 592650 32378
rect -8726 32058 -8694 32294
rect -8458 32058 -8374 32294
rect -8138 32058 570986 32294
rect 571222 32058 571306 32294
rect 571542 32058 592062 32294
rect 592298 32058 592382 32294
rect 592618 32058 592650 32294
rect -8726 32026 592650 32058
rect -6806 28894 590730 28926
rect -6806 28658 -6774 28894
rect -6538 28658 -6454 28894
rect -6218 28658 567266 28894
rect 567502 28658 567586 28894
rect 567822 28658 590142 28894
rect 590378 28658 590462 28894
rect 590698 28658 590730 28894
rect -6806 28574 590730 28658
rect -6806 28338 -6774 28574
rect -6538 28338 -6454 28574
rect -6218 28338 567266 28574
rect 567502 28338 567586 28574
rect 567822 28338 590142 28574
rect 590378 28338 590462 28574
rect 590698 28338 590730 28574
rect -6806 28306 590730 28338
rect -4886 25174 588810 25206
rect -4886 24938 -4854 25174
rect -4618 24938 -4534 25174
rect -4298 24938 588222 25174
rect 588458 24938 588542 25174
rect 588778 24938 588810 25174
rect -4886 24854 588810 24938
rect -4886 24618 -4854 24854
rect -4618 24618 -4534 24854
rect -4298 24618 588222 24854
rect 588458 24618 588542 24854
rect 588778 24618 588810 24854
rect -4886 24586 588810 24618
rect -2966 21454 586890 21486
rect -2966 21218 -2934 21454
rect -2698 21218 -2614 21454
rect -2378 21218 23610 21454
rect 23846 21218 54330 21454
rect 54566 21218 85050 21454
rect 85286 21218 115770 21454
rect 116006 21218 146490 21454
rect 146726 21218 177210 21454
rect 177446 21218 207930 21454
rect 208166 21218 238650 21454
rect 238886 21218 269370 21454
rect 269606 21218 300090 21454
rect 300326 21218 330810 21454
rect 331046 21218 361530 21454
rect 361766 21218 392250 21454
rect 392486 21218 422970 21454
rect 423206 21218 453690 21454
rect 453926 21218 484410 21454
rect 484646 21218 515130 21454
rect 515366 21218 545850 21454
rect 546086 21218 586302 21454
rect 586538 21218 586622 21454
rect 586858 21218 586890 21454
rect -2966 21134 586890 21218
rect -2966 20898 -2934 21134
rect -2698 20898 -2614 21134
rect -2378 20898 23610 21134
rect 23846 20898 54330 21134
rect 54566 20898 85050 21134
rect 85286 20898 115770 21134
rect 116006 20898 146490 21134
rect 146726 20898 177210 21134
rect 177446 20898 207930 21134
rect 208166 20898 238650 21134
rect 238886 20898 269370 21134
rect 269606 20898 300090 21134
rect 300326 20898 330810 21134
rect 331046 20898 361530 21134
rect 361766 20898 392250 21134
rect 392486 20898 422970 21134
rect 423206 20898 453690 21134
rect 453926 20898 484410 21134
rect 484646 20898 515130 21134
rect 515366 20898 545850 21134
rect 546086 20898 586302 21134
rect 586538 20898 586622 21134
rect 586858 20898 586890 21134
rect -2966 20866 586890 20898
rect -8726 14614 592650 14646
rect -8726 14378 -7734 14614
rect -7498 14378 -7414 14614
rect -7178 14378 591102 14614
rect 591338 14378 591422 14614
rect 591658 14378 592650 14614
rect -8726 14294 592650 14378
rect -8726 14058 -7734 14294
rect -7498 14058 -7414 14294
rect -7178 14058 591102 14294
rect 591338 14058 591422 14294
rect 591658 14058 592650 14294
rect -8726 14026 592650 14058
rect -6806 10894 590730 10926
rect -6806 10658 -5814 10894
rect -5578 10658 -5494 10894
rect -5258 10658 589182 10894
rect 589418 10658 589502 10894
rect 589738 10658 590730 10894
rect -6806 10574 590730 10658
rect -6806 10338 -5814 10574
rect -5578 10338 -5494 10574
rect -5258 10338 589182 10574
rect 589418 10338 589502 10574
rect 589738 10338 590730 10574
rect -6806 10306 590730 10338
rect -4886 7174 588810 7206
rect -4886 6938 -3894 7174
rect -3658 6938 -3574 7174
rect -3338 6938 581546 7174
rect 581782 6938 581866 7174
rect 582102 6938 587262 7174
rect 587498 6938 587582 7174
rect 587818 6938 588810 7174
rect -4886 6854 588810 6938
rect -4886 6618 -3894 6854
rect -3658 6618 -3574 6854
rect -3338 6618 581546 6854
rect 581782 6618 581866 6854
rect 582102 6618 587262 6854
rect 587498 6618 587582 6854
rect 587818 6618 588810 6854
rect -4886 6586 588810 6618
rect -2966 3454 586890 3486
rect -2966 3218 -1974 3454
rect -1738 3218 -1654 3454
rect -1418 3218 8250 3454
rect 8486 3218 38970 3454
rect 39206 3218 69690 3454
rect 69926 3218 100410 3454
rect 100646 3218 131130 3454
rect 131366 3218 161850 3454
rect 162086 3218 192570 3454
rect 192806 3218 223290 3454
rect 223526 3218 254010 3454
rect 254246 3218 284730 3454
rect 284966 3218 315450 3454
rect 315686 3218 346170 3454
rect 346406 3218 376890 3454
rect 377126 3218 407610 3454
rect 407846 3218 438330 3454
rect 438566 3218 469050 3454
rect 469286 3218 499770 3454
rect 500006 3218 530490 3454
rect 530726 3218 561210 3454
rect 561446 3218 577826 3454
rect 578062 3218 578146 3454
rect 578382 3218 585342 3454
rect 585578 3218 585662 3454
rect 585898 3218 586890 3454
rect -2966 3134 586890 3218
rect -2966 2898 -1974 3134
rect -1738 2898 -1654 3134
rect -1418 2898 8250 3134
rect 8486 2898 38970 3134
rect 39206 2898 69690 3134
rect 69926 2898 100410 3134
rect 100646 2898 131130 3134
rect 131366 2898 161850 3134
rect 162086 2898 192570 3134
rect 192806 2898 223290 3134
rect 223526 2898 254010 3134
rect 254246 2898 284730 3134
rect 284966 2898 315450 3134
rect 315686 2898 346170 3134
rect 346406 2898 376890 3134
rect 377126 2898 407610 3134
rect 407846 2898 438330 3134
rect 438566 2898 469050 3134
rect 469286 2898 499770 3134
rect 500006 2898 530490 3134
rect 530726 2898 561210 3134
rect 561446 2898 577826 3134
rect 578062 2898 578146 3134
rect 578382 2898 585342 3134
rect 585578 2898 585662 3134
rect 585898 2898 586890 3134
rect -2966 2866 586890 2898
rect -2006 -346 585930 -314
rect -2006 -582 -1974 -346
rect -1738 -582 -1654 -346
rect -1418 -582 577826 -346
rect 578062 -582 578146 -346
rect 578382 -582 585342 -346
rect 585578 -582 585662 -346
rect 585898 -582 585930 -346
rect -2006 -666 585930 -582
rect -2006 -902 -1974 -666
rect -1738 -902 -1654 -666
rect -1418 -902 577826 -666
rect 578062 -902 578146 -666
rect 578382 -902 585342 -666
rect 585578 -902 585662 -666
rect 585898 -902 585930 -666
rect -2006 -934 585930 -902
rect -2966 -1306 586890 -1274
rect -2966 -1542 -2934 -1306
rect -2698 -1542 -2614 -1306
rect -2378 -1542 586302 -1306
rect 586538 -1542 586622 -1306
rect 586858 -1542 586890 -1306
rect -2966 -1626 586890 -1542
rect -2966 -1862 -2934 -1626
rect -2698 -1862 -2614 -1626
rect -2378 -1862 586302 -1626
rect 586538 -1862 586622 -1626
rect 586858 -1862 586890 -1626
rect -2966 -1894 586890 -1862
rect -3926 -2266 587850 -2234
rect -3926 -2502 -3894 -2266
rect -3658 -2502 -3574 -2266
rect -3338 -2502 5546 -2266
rect 5782 -2502 5866 -2266
rect 6102 -2502 41546 -2266
rect 41782 -2502 41866 -2266
rect 42102 -2502 77546 -2266
rect 77782 -2502 77866 -2266
rect 78102 -2502 113546 -2266
rect 113782 -2502 113866 -2266
rect 114102 -2502 149546 -2266
rect 149782 -2502 149866 -2266
rect 150102 -2502 185546 -2266
rect 185782 -2502 185866 -2266
rect 186102 -2502 221546 -2266
rect 221782 -2502 221866 -2266
rect 222102 -2502 257546 -2266
rect 257782 -2502 257866 -2266
rect 258102 -2502 293546 -2266
rect 293782 -2502 293866 -2266
rect 294102 -2502 329546 -2266
rect 329782 -2502 329866 -2266
rect 330102 -2502 365546 -2266
rect 365782 -2502 365866 -2266
rect 366102 -2502 401546 -2266
rect 401782 -2502 401866 -2266
rect 402102 -2502 437546 -2266
rect 437782 -2502 437866 -2266
rect 438102 -2502 473546 -2266
rect 473782 -2502 473866 -2266
rect 474102 -2502 509546 -2266
rect 509782 -2502 509866 -2266
rect 510102 -2502 545546 -2266
rect 545782 -2502 545866 -2266
rect 546102 -2502 581546 -2266
rect 581782 -2502 581866 -2266
rect 582102 -2502 587262 -2266
rect 587498 -2502 587582 -2266
rect 587818 -2502 587850 -2266
rect -3926 -2586 587850 -2502
rect -3926 -2822 -3894 -2586
rect -3658 -2822 -3574 -2586
rect -3338 -2822 5546 -2586
rect 5782 -2822 5866 -2586
rect 6102 -2822 41546 -2586
rect 41782 -2822 41866 -2586
rect 42102 -2822 77546 -2586
rect 77782 -2822 77866 -2586
rect 78102 -2822 113546 -2586
rect 113782 -2822 113866 -2586
rect 114102 -2822 149546 -2586
rect 149782 -2822 149866 -2586
rect 150102 -2822 185546 -2586
rect 185782 -2822 185866 -2586
rect 186102 -2822 221546 -2586
rect 221782 -2822 221866 -2586
rect 222102 -2822 257546 -2586
rect 257782 -2822 257866 -2586
rect 258102 -2822 293546 -2586
rect 293782 -2822 293866 -2586
rect 294102 -2822 329546 -2586
rect 329782 -2822 329866 -2586
rect 330102 -2822 365546 -2586
rect 365782 -2822 365866 -2586
rect 366102 -2822 401546 -2586
rect 401782 -2822 401866 -2586
rect 402102 -2822 437546 -2586
rect 437782 -2822 437866 -2586
rect 438102 -2822 473546 -2586
rect 473782 -2822 473866 -2586
rect 474102 -2822 509546 -2586
rect 509782 -2822 509866 -2586
rect 510102 -2822 545546 -2586
rect 545782 -2822 545866 -2586
rect 546102 -2822 581546 -2586
rect 581782 -2822 581866 -2586
rect 582102 -2822 587262 -2586
rect 587498 -2822 587582 -2586
rect 587818 -2822 587850 -2586
rect -3926 -2854 587850 -2822
rect -4886 -3226 588810 -3194
rect -4886 -3462 -4854 -3226
rect -4618 -3462 -4534 -3226
rect -4298 -3462 23546 -3226
rect 23782 -3462 23866 -3226
rect 24102 -3462 59546 -3226
rect 59782 -3462 59866 -3226
rect 60102 -3462 95546 -3226
rect 95782 -3462 95866 -3226
rect 96102 -3462 131546 -3226
rect 131782 -3462 131866 -3226
rect 132102 -3462 167546 -3226
rect 167782 -3462 167866 -3226
rect 168102 -3462 203546 -3226
rect 203782 -3462 203866 -3226
rect 204102 -3462 239546 -3226
rect 239782 -3462 239866 -3226
rect 240102 -3462 275546 -3226
rect 275782 -3462 275866 -3226
rect 276102 -3462 311546 -3226
rect 311782 -3462 311866 -3226
rect 312102 -3462 347546 -3226
rect 347782 -3462 347866 -3226
rect 348102 -3462 383546 -3226
rect 383782 -3462 383866 -3226
rect 384102 -3462 419546 -3226
rect 419782 -3462 419866 -3226
rect 420102 -3462 455546 -3226
rect 455782 -3462 455866 -3226
rect 456102 -3462 491546 -3226
rect 491782 -3462 491866 -3226
rect 492102 -3462 527546 -3226
rect 527782 -3462 527866 -3226
rect 528102 -3462 563546 -3226
rect 563782 -3462 563866 -3226
rect 564102 -3462 588222 -3226
rect 588458 -3462 588542 -3226
rect 588778 -3462 588810 -3226
rect -4886 -3546 588810 -3462
rect -4886 -3782 -4854 -3546
rect -4618 -3782 -4534 -3546
rect -4298 -3782 23546 -3546
rect 23782 -3782 23866 -3546
rect 24102 -3782 59546 -3546
rect 59782 -3782 59866 -3546
rect 60102 -3782 95546 -3546
rect 95782 -3782 95866 -3546
rect 96102 -3782 131546 -3546
rect 131782 -3782 131866 -3546
rect 132102 -3782 167546 -3546
rect 167782 -3782 167866 -3546
rect 168102 -3782 203546 -3546
rect 203782 -3782 203866 -3546
rect 204102 -3782 239546 -3546
rect 239782 -3782 239866 -3546
rect 240102 -3782 275546 -3546
rect 275782 -3782 275866 -3546
rect 276102 -3782 311546 -3546
rect 311782 -3782 311866 -3546
rect 312102 -3782 347546 -3546
rect 347782 -3782 347866 -3546
rect 348102 -3782 383546 -3546
rect 383782 -3782 383866 -3546
rect 384102 -3782 419546 -3546
rect 419782 -3782 419866 -3546
rect 420102 -3782 455546 -3546
rect 455782 -3782 455866 -3546
rect 456102 -3782 491546 -3546
rect 491782 -3782 491866 -3546
rect 492102 -3782 527546 -3546
rect 527782 -3782 527866 -3546
rect 528102 -3782 563546 -3546
rect 563782 -3782 563866 -3546
rect 564102 -3782 588222 -3546
rect 588458 -3782 588542 -3546
rect 588778 -3782 588810 -3546
rect -4886 -3814 588810 -3782
rect -5846 -4186 589770 -4154
rect -5846 -4422 -5814 -4186
rect -5578 -4422 -5494 -4186
rect -5258 -4422 9266 -4186
rect 9502 -4422 9586 -4186
rect 9822 -4422 45266 -4186
rect 45502 -4422 45586 -4186
rect 45822 -4422 81266 -4186
rect 81502 -4422 81586 -4186
rect 81822 -4422 117266 -4186
rect 117502 -4422 117586 -4186
rect 117822 -4422 153266 -4186
rect 153502 -4422 153586 -4186
rect 153822 -4422 189266 -4186
rect 189502 -4422 189586 -4186
rect 189822 -4422 225266 -4186
rect 225502 -4422 225586 -4186
rect 225822 -4422 261266 -4186
rect 261502 -4422 261586 -4186
rect 261822 -4422 297266 -4186
rect 297502 -4422 297586 -4186
rect 297822 -4422 333266 -4186
rect 333502 -4422 333586 -4186
rect 333822 -4422 369266 -4186
rect 369502 -4422 369586 -4186
rect 369822 -4422 405266 -4186
rect 405502 -4422 405586 -4186
rect 405822 -4422 441266 -4186
rect 441502 -4422 441586 -4186
rect 441822 -4422 477266 -4186
rect 477502 -4422 477586 -4186
rect 477822 -4422 513266 -4186
rect 513502 -4422 513586 -4186
rect 513822 -4422 549266 -4186
rect 549502 -4422 549586 -4186
rect 549822 -4422 589182 -4186
rect 589418 -4422 589502 -4186
rect 589738 -4422 589770 -4186
rect -5846 -4506 589770 -4422
rect -5846 -4742 -5814 -4506
rect -5578 -4742 -5494 -4506
rect -5258 -4742 9266 -4506
rect 9502 -4742 9586 -4506
rect 9822 -4742 45266 -4506
rect 45502 -4742 45586 -4506
rect 45822 -4742 81266 -4506
rect 81502 -4742 81586 -4506
rect 81822 -4742 117266 -4506
rect 117502 -4742 117586 -4506
rect 117822 -4742 153266 -4506
rect 153502 -4742 153586 -4506
rect 153822 -4742 189266 -4506
rect 189502 -4742 189586 -4506
rect 189822 -4742 225266 -4506
rect 225502 -4742 225586 -4506
rect 225822 -4742 261266 -4506
rect 261502 -4742 261586 -4506
rect 261822 -4742 297266 -4506
rect 297502 -4742 297586 -4506
rect 297822 -4742 333266 -4506
rect 333502 -4742 333586 -4506
rect 333822 -4742 369266 -4506
rect 369502 -4742 369586 -4506
rect 369822 -4742 405266 -4506
rect 405502 -4742 405586 -4506
rect 405822 -4742 441266 -4506
rect 441502 -4742 441586 -4506
rect 441822 -4742 477266 -4506
rect 477502 -4742 477586 -4506
rect 477822 -4742 513266 -4506
rect 513502 -4742 513586 -4506
rect 513822 -4742 549266 -4506
rect 549502 -4742 549586 -4506
rect 549822 -4742 589182 -4506
rect 589418 -4742 589502 -4506
rect 589738 -4742 589770 -4506
rect -5846 -4774 589770 -4742
rect -6806 -5146 590730 -5114
rect -6806 -5382 -6774 -5146
rect -6538 -5382 -6454 -5146
rect -6218 -5382 27266 -5146
rect 27502 -5382 27586 -5146
rect 27822 -5382 63266 -5146
rect 63502 -5382 63586 -5146
rect 63822 -5382 99266 -5146
rect 99502 -5382 99586 -5146
rect 99822 -5382 135266 -5146
rect 135502 -5382 135586 -5146
rect 135822 -5382 171266 -5146
rect 171502 -5382 171586 -5146
rect 171822 -5382 207266 -5146
rect 207502 -5382 207586 -5146
rect 207822 -5382 243266 -5146
rect 243502 -5382 243586 -5146
rect 243822 -5382 279266 -5146
rect 279502 -5382 279586 -5146
rect 279822 -5382 315266 -5146
rect 315502 -5382 315586 -5146
rect 315822 -5382 351266 -5146
rect 351502 -5382 351586 -5146
rect 351822 -5382 387266 -5146
rect 387502 -5382 387586 -5146
rect 387822 -5382 423266 -5146
rect 423502 -5382 423586 -5146
rect 423822 -5382 459266 -5146
rect 459502 -5382 459586 -5146
rect 459822 -5382 495266 -5146
rect 495502 -5382 495586 -5146
rect 495822 -5382 531266 -5146
rect 531502 -5382 531586 -5146
rect 531822 -5382 567266 -5146
rect 567502 -5382 567586 -5146
rect 567822 -5382 590142 -5146
rect 590378 -5382 590462 -5146
rect 590698 -5382 590730 -5146
rect -6806 -5466 590730 -5382
rect -6806 -5702 -6774 -5466
rect -6538 -5702 -6454 -5466
rect -6218 -5702 27266 -5466
rect 27502 -5702 27586 -5466
rect 27822 -5702 63266 -5466
rect 63502 -5702 63586 -5466
rect 63822 -5702 99266 -5466
rect 99502 -5702 99586 -5466
rect 99822 -5702 135266 -5466
rect 135502 -5702 135586 -5466
rect 135822 -5702 171266 -5466
rect 171502 -5702 171586 -5466
rect 171822 -5702 207266 -5466
rect 207502 -5702 207586 -5466
rect 207822 -5702 243266 -5466
rect 243502 -5702 243586 -5466
rect 243822 -5702 279266 -5466
rect 279502 -5702 279586 -5466
rect 279822 -5702 315266 -5466
rect 315502 -5702 315586 -5466
rect 315822 -5702 351266 -5466
rect 351502 -5702 351586 -5466
rect 351822 -5702 387266 -5466
rect 387502 -5702 387586 -5466
rect 387822 -5702 423266 -5466
rect 423502 -5702 423586 -5466
rect 423822 -5702 459266 -5466
rect 459502 -5702 459586 -5466
rect 459822 -5702 495266 -5466
rect 495502 -5702 495586 -5466
rect 495822 -5702 531266 -5466
rect 531502 -5702 531586 -5466
rect 531822 -5702 567266 -5466
rect 567502 -5702 567586 -5466
rect 567822 -5702 590142 -5466
rect 590378 -5702 590462 -5466
rect 590698 -5702 590730 -5466
rect -6806 -5734 590730 -5702
rect -7766 -6106 591690 -6074
rect -7766 -6342 -7734 -6106
rect -7498 -6342 -7414 -6106
rect -7178 -6342 12986 -6106
rect 13222 -6342 13306 -6106
rect 13542 -6342 48986 -6106
rect 49222 -6342 49306 -6106
rect 49542 -6342 84986 -6106
rect 85222 -6342 85306 -6106
rect 85542 -6342 120986 -6106
rect 121222 -6342 121306 -6106
rect 121542 -6342 156986 -6106
rect 157222 -6342 157306 -6106
rect 157542 -6342 192986 -6106
rect 193222 -6342 193306 -6106
rect 193542 -6342 228986 -6106
rect 229222 -6342 229306 -6106
rect 229542 -6342 264986 -6106
rect 265222 -6342 265306 -6106
rect 265542 -6342 300986 -6106
rect 301222 -6342 301306 -6106
rect 301542 -6342 336986 -6106
rect 337222 -6342 337306 -6106
rect 337542 -6342 372986 -6106
rect 373222 -6342 373306 -6106
rect 373542 -6342 408986 -6106
rect 409222 -6342 409306 -6106
rect 409542 -6342 444986 -6106
rect 445222 -6342 445306 -6106
rect 445542 -6342 480986 -6106
rect 481222 -6342 481306 -6106
rect 481542 -6342 516986 -6106
rect 517222 -6342 517306 -6106
rect 517542 -6342 552986 -6106
rect 553222 -6342 553306 -6106
rect 553542 -6342 591102 -6106
rect 591338 -6342 591422 -6106
rect 591658 -6342 591690 -6106
rect -7766 -6426 591690 -6342
rect -7766 -6662 -7734 -6426
rect -7498 -6662 -7414 -6426
rect -7178 -6662 12986 -6426
rect 13222 -6662 13306 -6426
rect 13542 -6662 48986 -6426
rect 49222 -6662 49306 -6426
rect 49542 -6662 84986 -6426
rect 85222 -6662 85306 -6426
rect 85542 -6662 120986 -6426
rect 121222 -6662 121306 -6426
rect 121542 -6662 156986 -6426
rect 157222 -6662 157306 -6426
rect 157542 -6662 192986 -6426
rect 193222 -6662 193306 -6426
rect 193542 -6662 228986 -6426
rect 229222 -6662 229306 -6426
rect 229542 -6662 264986 -6426
rect 265222 -6662 265306 -6426
rect 265542 -6662 300986 -6426
rect 301222 -6662 301306 -6426
rect 301542 -6662 336986 -6426
rect 337222 -6662 337306 -6426
rect 337542 -6662 372986 -6426
rect 373222 -6662 373306 -6426
rect 373542 -6662 408986 -6426
rect 409222 -6662 409306 -6426
rect 409542 -6662 444986 -6426
rect 445222 -6662 445306 -6426
rect 445542 -6662 480986 -6426
rect 481222 -6662 481306 -6426
rect 481542 -6662 516986 -6426
rect 517222 -6662 517306 -6426
rect 517542 -6662 552986 -6426
rect 553222 -6662 553306 -6426
rect 553542 -6662 591102 -6426
rect 591338 -6662 591422 -6426
rect 591658 -6662 591690 -6426
rect -7766 -6694 591690 -6662
rect -8726 -7066 592650 -7034
rect -8726 -7302 -8694 -7066
rect -8458 -7302 -8374 -7066
rect -8138 -7302 30986 -7066
rect 31222 -7302 31306 -7066
rect 31542 -7302 66986 -7066
rect 67222 -7302 67306 -7066
rect 67542 -7302 102986 -7066
rect 103222 -7302 103306 -7066
rect 103542 -7302 138986 -7066
rect 139222 -7302 139306 -7066
rect 139542 -7302 174986 -7066
rect 175222 -7302 175306 -7066
rect 175542 -7302 210986 -7066
rect 211222 -7302 211306 -7066
rect 211542 -7302 246986 -7066
rect 247222 -7302 247306 -7066
rect 247542 -7302 282986 -7066
rect 283222 -7302 283306 -7066
rect 283542 -7302 318986 -7066
rect 319222 -7302 319306 -7066
rect 319542 -7302 354986 -7066
rect 355222 -7302 355306 -7066
rect 355542 -7302 390986 -7066
rect 391222 -7302 391306 -7066
rect 391542 -7302 426986 -7066
rect 427222 -7302 427306 -7066
rect 427542 -7302 462986 -7066
rect 463222 -7302 463306 -7066
rect 463542 -7302 498986 -7066
rect 499222 -7302 499306 -7066
rect 499542 -7302 534986 -7066
rect 535222 -7302 535306 -7066
rect 535542 -7302 570986 -7066
rect 571222 -7302 571306 -7066
rect 571542 -7302 592062 -7066
rect 592298 -7302 592382 -7066
rect 592618 -7302 592650 -7066
rect -8726 -7386 592650 -7302
rect -8726 -7622 -8694 -7386
rect -8458 -7622 -8374 -7386
rect -8138 -7622 30986 -7386
rect 31222 -7622 31306 -7386
rect 31542 -7622 66986 -7386
rect 67222 -7622 67306 -7386
rect 67542 -7622 102986 -7386
rect 103222 -7622 103306 -7386
rect 103542 -7622 138986 -7386
rect 139222 -7622 139306 -7386
rect 139542 -7622 174986 -7386
rect 175222 -7622 175306 -7386
rect 175542 -7622 210986 -7386
rect 211222 -7622 211306 -7386
rect 211542 -7622 246986 -7386
rect 247222 -7622 247306 -7386
rect 247542 -7622 282986 -7386
rect 283222 -7622 283306 -7386
rect 283542 -7622 318986 -7386
rect 319222 -7622 319306 -7386
rect 319542 -7622 354986 -7386
rect 355222 -7622 355306 -7386
rect 355542 -7622 390986 -7386
rect 391222 -7622 391306 -7386
rect 391542 -7622 426986 -7386
rect 427222 -7622 427306 -7386
rect 427542 -7622 462986 -7386
rect 463222 -7622 463306 -7386
rect 463542 -7622 498986 -7386
rect 499222 -7622 499306 -7386
rect 499542 -7622 534986 -7386
rect 535222 -7622 535306 -7386
rect 535542 -7622 570986 -7386
rect 571222 -7622 571306 -7386
rect 571542 -7622 592062 -7386
rect 592298 -7622 592382 -7386
rect 592618 -7622 592650 -7386
rect -8726 -7654 592650 -7622
use user_proj  mprj
timestamp 1639150748
transform 1 0 4000 0 1 0
box 566 0 559438 700000
<< labels >>
rlabel metal3 s 583520 285276 584960 285516 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal3 s -960 697220 480 697460 4 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal3 s -960 644996 480 645236 4 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal3 s -960 592908 480 593148 4 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 583520 338452 584960 338692 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal3 s -960 540684 480 540924 4 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal3 s -960 488596 480 488836 4 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal3 s -960 436508 480 436748 4 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal3 s -960 384284 480 384524 4 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -960 332196 480 332436 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -960 279972 480 280212 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -960 227884 480 228124 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -960 175796 480 176036 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -960 123572 480 123812 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 583520 391628 584960 391868 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 583520 444668 584960 444908 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 583520 497844 584960 498084 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 583520 551020 584960 551260 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 583520 604060 584960 604300 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 583520 657236 584960 657476 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 583520 6476 584960 6716 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 583520 457996 584960 458236 6 io_in[10]
port 30 nsew signal input
rlabel metal3 s 583520 511172 584960 511412 6 io_in[11]
port 31 nsew signal input
rlabel metal3 s 583520 564212 584960 564452 6 io_in[12]
port 32 nsew signal input
rlabel metal3 s 583520 617388 584960 617628 6 io_in[13]
port 33 nsew signal input
rlabel metal3 s 583520 670564 584960 670804 6 io_in[14]
port 34 nsew signal input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 35 nsew signal input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 36 nsew signal input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 37 nsew signal input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 38 nsew signal input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 39 nsew signal input
rlabel metal3 s 583520 46188 584960 46428 6 io_in[1]
port 40 nsew signal input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 41 nsew signal input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 42 nsew signal input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 43 nsew signal input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 44 nsew signal input
rlabel metal3 s -960 684164 480 684404 4 io_in[24]
port 45 nsew signal input
rlabel metal3 s -960 631940 480 632180 4 io_in[25]
port 46 nsew signal input
rlabel metal3 s -960 579852 480 580092 4 io_in[26]
port 47 nsew signal input
rlabel metal3 s -960 527764 480 528004 4 io_in[27]
port 48 nsew signal input
rlabel metal3 s -960 475540 480 475780 4 io_in[28]
port 49 nsew signal input
rlabel metal3 s -960 423452 480 423692 4 io_in[29]
port 50 nsew signal input
rlabel metal3 s 583520 86036 584960 86276 6 io_in[2]
port 51 nsew signal input
rlabel metal3 s -960 371228 480 371468 4 io_in[30]
port 52 nsew signal input
rlabel metal3 s -960 319140 480 319380 4 io_in[31]
port 53 nsew signal input
rlabel metal3 s -960 267052 480 267292 4 io_in[32]
port 54 nsew signal input
rlabel metal3 s -960 214828 480 215068 4 io_in[33]
port 55 nsew signal input
rlabel metal3 s -960 162740 480 162980 4 io_in[34]
port 56 nsew signal input
rlabel metal3 s -960 110516 480 110756 4 io_in[35]
port 57 nsew signal input
rlabel metal3 s -960 71484 480 71724 4 io_in[36]
port 58 nsew signal input
rlabel metal3 s -960 32316 480 32556 4 io_in[37]
port 59 nsew signal input
rlabel metal3 s 583520 125884 584960 126124 6 io_in[3]
port 60 nsew signal input
rlabel metal3 s 583520 165732 584960 165972 6 io_in[4]
port 61 nsew signal input
rlabel metal3 s 583520 205580 584960 205820 6 io_in[5]
port 62 nsew signal input
rlabel metal3 s 583520 245428 584960 245668 6 io_in[6]
port 63 nsew signal input
rlabel metal3 s 583520 298604 584960 298844 6 io_in[7]
port 64 nsew signal input
rlabel metal3 s 583520 351780 584960 352020 6 io_in[8]
port 65 nsew signal input
rlabel metal3 s 583520 404820 584960 405060 6 io_in[9]
port 66 nsew signal input
rlabel metal3 s 583520 32996 584960 33236 6 io_oeb[0]
port 67 nsew signal tristate
rlabel metal3 s 583520 484516 584960 484756 6 io_oeb[10]
port 68 nsew signal tristate
rlabel metal3 s 583520 537692 584960 537932 6 io_oeb[11]
port 69 nsew signal tristate
rlabel metal3 s 583520 590868 584960 591108 6 io_oeb[12]
port 70 nsew signal tristate
rlabel metal3 s 583520 643908 584960 644148 6 io_oeb[13]
port 71 nsew signal tristate
rlabel metal3 s 583520 697084 584960 697324 6 io_oeb[14]
port 72 nsew signal tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 73 nsew signal tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 74 nsew signal tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 75 nsew signal tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 76 nsew signal tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 77 nsew signal tristate
rlabel metal3 s 583520 72844 584960 73084 6 io_oeb[1]
port 78 nsew signal tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 79 nsew signal tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 80 nsew signal tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 81 nsew signal tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 82 nsew signal tristate
rlabel metal3 s -960 658052 480 658292 4 io_oeb[24]
port 83 nsew signal tristate
rlabel metal3 s -960 605964 480 606204 4 io_oeb[25]
port 84 nsew signal tristate
rlabel metal3 s -960 553740 480 553980 4 io_oeb[26]
port 85 nsew signal tristate
rlabel metal3 s -960 501652 480 501892 4 io_oeb[27]
port 86 nsew signal tristate
rlabel metal3 s -960 449428 480 449668 4 io_oeb[28]
port 87 nsew signal tristate
rlabel metal3 s -960 397340 480 397580 4 io_oeb[29]
port 88 nsew signal tristate
rlabel metal3 s 583520 112692 584960 112932 6 io_oeb[2]
port 89 nsew signal tristate
rlabel metal3 s -960 345252 480 345492 4 io_oeb[30]
port 90 nsew signal tristate
rlabel metal3 s -960 293028 480 293268 4 io_oeb[31]
port 91 nsew signal tristate
rlabel metal3 s -960 240940 480 241180 4 io_oeb[32]
port 92 nsew signal tristate
rlabel metal3 s -960 188716 480 188956 4 io_oeb[33]
port 93 nsew signal tristate
rlabel metal3 s -960 136628 480 136868 4 io_oeb[34]
port 94 nsew signal tristate
rlabel metal3 s -960 84540 480 84780 4 io_oeb[35]
port 95 nsew signal tristate
rlabel metal3 s -960 45372 480 45612 4 io_oeb[36]
port 96 nsew signal tristate
rlabel metal3 s -960 6340 480 6580 4 io_oeb[37]
port 97 nsew signal tristate
rlabel metal3 s 583520 152540 584960 152780 6 io_oeb[3]
port 98 nsew signal tristate
rlabel metal3 s 583520 192388 584960 192628 6 io_oeb[4]
port 99 nsew signal tristate
rlabel metal3 s 583520 232236 584960 232476 6 io_oeb[5]
port 100 nsew signal tristate
rlabel metal3 s 583520 272084 584960 272324 6 io_oeb[6]
port 101 nsew signal tristate
rlabel metal3 s 583520 325124 584960 325364 6 io_oeb[7]
port 102 nsew signal tristate
rlabel metal3 s 583520 378300 584960 378540 6 io_oeb[8]
port 103 nsew signal tristate
rlabel metal3 s 583520 431476 584960 431716 6 io_oeb[9]
port 104 nsew signal tristate
rlabel metal3 s 583520 19668 584960 19908 6 io_out[0]
port 105 nsew signal tristate
rlabel metal3 s 583520 471324 584960 471564 6 io_out[10]
port 106 nsew signal tristate
rlabel metal3 s 583520 524364 584960 524604 6 io_out[11]
port 107 nsew signal tristate
rlabel metal3 s 583520 577540 584960 577780 6 io_out[12]
port 108 nsew signal tristate
rlabel metal3 s 583520 630716 584960 630956 6 io_out[13]
port 109 nsew signal tristate
rlabel metal3 s 583520 683756 584960 683996 6 io_out[14]
port 110 nsew signal tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 111 nsew signal tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 112 nsew signal tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 113 nsew signal tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 114 nsew signal tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 115 nsew signal tristate
rlabel metal3 s 583520 59516 584960 59756 6 io_out[1]
port 116 nsew signal tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 117 nsew signal tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 118 nsew signal tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 119 nsew signal tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 120 nsew signal tristate
rlabel metal3 s -960 671108 480 671348 4 io_out[24]
port 121 nsew signal tristate
rlabel metal3 s -960 619020 480 619260 4 io_out[25]
port 122 nsew signal tristate
rlabel metal3 s -960 566796 480 567036 4 io_out[26]
port 123 nsew signal tristate
rlabel metal3 s -960 514708 480 514948 4 io_out[27]
port 124 nsew signal tristate
rlabel metal3 s -960 462484 480 462724 4 io_out[28]
port 125 nsew signal tristate
rlabel metal3 s -960 410396 480 410636 4 io_out[29]
port 126 nsew signal tristate
rlabel metal3 s 583520 99364 584960 99604 6 io_out[2]
port 127 nsew signal tristate
rlabel metal3 s -960 358308 480 358548 4 io_out[30]
port 128 nsew signal tristate
rlabel metal3 s -960 306084 480 306324 4 io_out[31]
port 129 nsew signal tristate
rlabel metal3 s -960 253996 480 254236 4 io_out[32]
port 130 nsew signal tristate
rlabel metal3 s -960 201772 480 202012 4 io_out[33]
port 131 nsew signal tristate
rlabel metal3 s -960 149684 480 149924 4 io_out[34]
port 132 nsew signal tristate
rlabel metal3 s -960 97460 480 97700 4 io_out[35]
port 133 nsew signal tristate
rlabel metal3 s -960 58428 480 58668 4 io_out[36]
port 134 nsew signal tristate
rlabel metal3 s -960 19260 480 19500 4 io_out[37]
port 135 nsew signal tristate
rlabel metal3 s 583520 139212 584960 139452 6 io_out[3]
port 136 nsew signal tristate
rlabel metal3 s 583520 179060 584960 179300 6 io_out[4]
port 137 nsew signal tristate
rlabel metal3 s 583520 218908 584960 219148 6 io_out[5]
port 138 nsew signal tristate
rlabel metal3 s 583520 258756 584960 258996 6 io_out[6]
port 139 nsew signal tristate
rlabel metal3 s 583520 311932 584960 312172 6 io_out[7]
port 140 nsew signal tristate
rlabel metal3 s 583520 364972 584960 365212 6 io_out[8]
port 141 nsew signal tristate
rlabel metal3 s 583520 418148 584960 418388 6 io_out[9]
port 142 nsew signal tristate
rlabel metal2 s 125846 -960 125958 480 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 480506 -960 480618 480 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 484002 -960 484114 480 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 487590 -960 487702 480 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 491086 -960 491198 480 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 494674 -960 494786 480 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 498170 -960 498282 480 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 501758 -960 501870 480 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 505346 -960 505458 480 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 508842 -960 508954 480 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 512430 -960 512542 480 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 161266 -960 161378 480 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 515926 -960 516038 480 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 519514 -960 519626 480 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 523010 -960 523122 480 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 526598 -960 526710 480 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 530094 -960 530206 480 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 533682 -960 533794 480 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 537178 -960 537290 480 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 540766 -960 540878 480 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 544354 -960 544466 480 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 547850 -960 547962 480 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 164854 -960 164966 480 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 551438 -960 551550 480 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 554934 -960 555046 480 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 558522 -960 558634 480 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 562018 -960 562130 480 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 565606 -960 565718 480 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 569102 -960 569214 480 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 572690 -960 572802 480 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 576278 -960 576390 480 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 168350 -960 168462 480 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 171938 -960 172050 480 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 175434 -960 175546 480 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 179022 -960 179134 480 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 182518 -960 182630 480 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 186106 -960 186218 480 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 189694 -960 189806 480 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 193190 -960 193302 480 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 129342 -960 129454 480 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 196778 -960 196890 480 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 200274 -960 200386 480 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 203862 -960 203974 480 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 207358 -960 207470 480 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 210946 -960 211058 480 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 214442 -960 214554 480 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 218030 -960 218142 480 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 221526 -960 221638 480 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 225114 -960 225226 480 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 228702 -960 228814 480 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 132930 -960 133042 480 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 232198 -960 232310 480 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 235786 -960 235898 480 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 239282 -960 239394 480 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 242870 -960 242982 480 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 246366 -960 246478 480 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 249954 -960 250066 480 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 253450 -960 253562 480 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 257038 -960 257150 480 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 260626 -960 260738 480 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 264122 -960 264234 480 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 136426 -960 136538 480 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 267710 -960 267822 480 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 271206 -960 271318 480 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 274794 -960 274906 480 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 278290 -960 278402 480 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 281878 -960 281990 480 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 285374 -960 285486 480 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 288962 -960 289074 480 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 292550 -960 292662 480 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 296046 -960 296158 480 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 299634 -960 299746 480 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 140014 -960 140126 480 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 303130 -960 303242 480 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 306718 -960 306830 480 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 310214 -960 310326 480 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 313802 -960 313914 480 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 317298 -960 317410 480 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 320886 -960 320998 480 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 324382 -960 324494 480 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 327970 -960 328082 480 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 331558 -960 331670 480 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 335054 -960 335166 480 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 143510 -960 143622 480 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 338642 -960 338754 480 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 342138 -960 342250 480 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 345726 -960 345838 480 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 349222 -960 349334 480 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 352810 -960 352922 480 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 356306 -960 356418 480 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 359894 -960 360006 480 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 363482 -960 363594 480 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 366978 -960 367090 480 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 370566 -960 370678 480 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 147098 -960 147210 480 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 374062 -960 374174 480 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 377650 -960 377762 480 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 381146 -960 381258 480 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 384734 -960 384846 480 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 388230 -960 388342 480 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 391818 -960 391930 480 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 395314 -960 395426 480 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 398902 -960 399014 480 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 402490 -960 402602 480 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 405986 -960 406098 480 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 150594 -960 150706 480 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 409574 -960 409686 480 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 413070 -960 413182 480 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 416658 -960 416770 480 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 420154 -960 420266 480 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 423742 -960 423854 480 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 427238 -960 427350 480 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 430826 -960 430938 480 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 434414 -960 434526 480 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 437910 -960 438022 480 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 441498 -960 441610 480 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 154182 -960 154294 480 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 444994 -960 445106 480 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 448582 -960 448694 480 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 452078 -960 452190 480 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 455666 -960 455778 480 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 459162 -960 459274 480 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 462750 -960 462862 480 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 466246 -960 466358 480 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 469834 -960 469946 480 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 473422 -960 473534 480 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 476918 -960 477030 480 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 157770 -960 157882 480 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 126950 -960 127062 480 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 481702 -960 481814 480 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 485198 -960 485310 480 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 488786 -960 488898 480 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 492282 -960 492394 480 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 495870 -960 495982 480 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 499366 -960 499478 480 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 502954 -960 503066 480 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 506450 -960 506562 480 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 510038 -960 510150 480 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 513534 -960 513646 480 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 162462 -960 162574 480 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 517122 -960 517234 480 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 520710 -960 520822 480 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 524206 -960 524318 480 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 527794 -960 527906 480 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 531290 -960 531402 480 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 534878 -960 534990 480 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 538374 -960 538486 480 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 541962 -960 542074 480 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 545458 -960 545570 480 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 549046 -960 549158 480 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 166050 -960 166162 480 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 552634 -960 552746 480 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 556130 -960 556242 480 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 559718 -960 559830 480 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 563214 -960 563326 480 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 566802 -960 566914 480 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 570298 -960 570410 480 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 573886 -960 573998 480 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 169546 -960 169658 480 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 173134 -960 173246 480 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 176630 -960 176742 480 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 180218 -960 180330 480 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 183714 -960 183826 480 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 187302 -960 187414 480 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 190798 -960 190910 480 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 194386 -960 194498 480 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 130538 -960 130650 480 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 197882 -960 197994 480 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 201470 -960 201582 480 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 205058 -960 205170 480 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 208554 -960 208666 480 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 212142 -960 212254 480 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 215638 -960 215750 480 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 219226 -960 219338 480 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 222722 -960 222834 480 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 226310 -960 226422 480 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 229806 -960 229918 480 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 134126 -960 134238 480 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 233394 -960 233506 480 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 236982 -960 237094 480 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 240478 -960 240590 480 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 244066 -960 244178 480 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 247562 -960 247674 480 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 251150 -960 251262 480 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 254646 -960 254758 480 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 258234 -960 258346 480 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 261730 -960 261842 480 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 265318 -960 265430 480 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 137622 -960 137734 480 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 268814 -960 268926 480 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 272402 -960 272514 480 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 275990 -960 276102 480 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 279486 -960 279598 480 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 283074 -960 283186 480 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 286570 -960 286682 480 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 290158 -960 290270 480 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 293654 -960 293766 480 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 297242 -960 297354 480 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 300738 -960 300850 480 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 141210 -960 141322 480 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 304326 -960 304438 480 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 307914 -960 308026 480 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 311410 -960 311522 480 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 314998 -960 315110 480 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 318494 -960 318606 480 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 322082 -960 322194 480 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 325578 -960 325690 480 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 329166 -960 329278 480 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 332662 -960 332774 480 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 336250 -960 336362 480 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 144706 -960 144818 480 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 339838 -960 339950 480 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 343334 -960 343446 480 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 346922 -960 347034 480 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 350418 -960 350530 480 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 354006 -960 354118 480 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 357502 -960 357614 480 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 361090 -960 361202 480 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 364586 -960 364698 480 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 368174 -960 368286 480 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 371670 -960 371782 480 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 148294 -960 148406 480 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 375258 -960 375370 480 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 378846 -960 378958 480 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 382342 -960 382454 480 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 385930 -960 386042 480 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 389426 -960 389538 480 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 393014 -960 393126 480 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 396510 -960 396622 480 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 400098 -960 400210 480 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 403594 -960 403706 480 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 407182 -960 407294 480 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 151790 -960 151902 480 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 410770 -960 410882 480 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 414266 -960 414378 480 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 417854 -960 417966 480 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 421350 -960 421462 480 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 424938 -960 425050 480 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 428434 -960 428546 480 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 432022 -960 432134 480 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 435518 -960 435630 480 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 439106 -960 439218 480 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 442602 -960 442714 480 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 155378 -960 155490 480 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 446190 -960 446302 480 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 449778 -960 449890 480 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 453274 -960 453386 480 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 456862 -960 456974 480 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 460358 -960 460470 480 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 463946 -960 464058 480 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 467442 -960 467554 480 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 471030 -960 471142 480 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 474526 -960 474638 480 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 478114 -960 478226 480 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 158874 -960 158986 480 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 128146 -960 128258 480 8 la_oenb[0]
port 399 nsew signal input
rlabel metal2 s 482806 -960 482918 480 8 la_oenb[100]
port 400 nsew signal input
rlabel metal2 s 486394 -960 486506 480 8 la_oenb[101]
port 401 nsew signal input
rlabel metal2 s 489890 -960 490002 480 8 la_oenb[102]
port 402 nsew signal input
rlabel metal2 s 493478 -960 493590 480 8 la_oenb[103]
port 403 nsew signal input
rlabel metal2 s 497066 -960 497178 480 8 la_oenb[104]
port 404 nsew signal input
rlabel metal2 s 500562 -960 500674 480 8 la_oenb[105]
port 405 nsew signal input
rlabel metal2 s 504150 -960 504262 480 8 la_oenb[106]
port 406 nsew signal input
rlabel metal2 s 507646 -960 507758 480 8 la_oenb[107]
port 407 nsew signal input
rlabel metal2 s 511234 -960 511346 480 8 la_oenb[108]
port 408 nsew signal input
rlabel metal2 s 514730 -960 514842 480 8 la_oenb[109]
port 409 nsew signal input
rlabel metal2 s 163658 -960 163770 480 8 la_oenb[10]
port 410 nsew signal input
rlabel metal2 s 518318 -960 518430 480 8 la_oenb[110]
port 411 nsew signal input
rlabel metal2 s 521814 -960 521926 480 8 la_oenb[111]
port 412 nsew signal input
rlabel metal2 s 525402 -960 525514 480 8 la_oenb[112]
port 413 nsew signal input
rlabel metal2 s 528990 -960 529102 480 8 la_oenb[113]
port 414 nsew signal input
rlabel metal2 s 532486 -960 532598 480 8 la_oenb[114]
port 415 nsew signal input
rlabel metal2 s 536074 -960 536186 480 8 la_oenb[115]
port 416 nsew signal input
rlabel metal2 s 539570 -960 539682 480 8 la_oenb[116]
port 417 nsew signal input
rlabel metal2 s 543158 -960 543270 480 8 la_oenb[117]
port 418 nsew signal input
rlabel metal2 s 546654 -960 546766 480 8 la_oenb[118]
port 419 nsew signal input
rlabel metal2 s 550242 -960 550354 480 8 la_oenb[119]
port 420 nsew signal input
rlabel metal2 s 167154 -960 167266 480 8 la_oenb[11]
port 421 nsew signal input
rlabel metal2 s 553738 -960 553850 480 8 la_oenb[120]
port 422 nsew signal input
rlabel metal2 s 557326 -960 557438 480 8 la_oenb[121]
port 423 nsew signal input
rlabel metal2 s 560822 -960 560934 480 8 la_oenb[122]
port 424 nsew signal input
rlabel metal2 s 564410 -960 564522 480 8 la_oenb[123]
port 425 nsew signal input
rlabel metal2 s 567998 -960 568110 480 8 la_oenb[124]
port 426 nsew signal input
rlabel metal2 s 571494 -960 571606 480 8 la_oenb[125]
port 427 nsew signal input
rlabel metal2 s 575082 -960 575194 480 8 la_oenb[126]
port 428 nsew signal input
rlabel metal2 s 578578 -960 578690 480 8 la_oenb[127]
port 429 nsew signal input
rlabel metal2 s 170742 -960 170854 480 8 la_oenb[12]
port 430 nsew signal input
rlabel metal2 s 174238 -960 174350 480 8 la_oenb[13]
port 431 nsew signal input
rlabel metal2 s 177826 -960 177938 480 8 la_oenb[14]
port 432 nsew signal input
rlabel metal2 s 181414 -960 181526 480 8 la_oenb[15]
port 433 nsew signal input
rlabel metal2 s 184910 -960 185022 480 8 la_oenb[16]
port 434 nsew signal input
rlabel metal2 s 188498 -960 188610 480 8 la_oenb[17]
port 435 nsew signal input
rlabel metal2 s 191994 -960 192106 480 8 la_oenb[18]
port 436 nsew signal input
rlabel metal2 s 195582 -960 195694 480 8 la_oenb[19]
port 437 nsew signal input
rlabel metal2 s 131734 -960 131846 480 8 la_oenb[1]
port 438 nsew signal input
rlabel metal2 s 199078 -960 199190 480 8 la_oenb[20]
port 439 nsew signal input
rlabel metal2 s 202666 -960 202778 480 8 la_oenb[21]
port 440 nsew signal input
rlabel metal2 s 206162 -960 206274 480 8 la_oenb[22]
port 441 nsew signal input
rlabel metal2 s 209750 -960 209862 480 8 la_oenb[23]
port 442 nsew signal input
rlabel metal2 s 213338 -960 213450 480 8 la_oenb[24]
port 443 nsew signal input
rlabel metal2 s 216834 -960 216946 480 8 la_oenb[25]
port 444 nsew signal input
rlabel metal2 s 220422 -960 220534 480 8 la_oenb[26]
port 445 nsew signal input
rlabel metal2 s 223918 -960 224030 480 8 la_oenb[27]
port 446 nsew signal input
rlabel metal2 s 227506 -960 227618 480 8 la_oenb[28]
port 447 nsew signal input
rlabel metal2 s 231002 -960 231114 480 8 la_oenb[29]
port 448 nsew signal input
rlabel metal2 s 135230 -960 135342 480 8 la_oenb[2]
port 449 nsew signal input
rlabel metal2 s 234590 -960 234702 480 8 la_oenb[30]
port 450 nsew signal input
rlabel metal2 s 238086 -960 238198 480 8 la_oenb[31]
port 451 nsew signal input
rlabel metal2 s 241674 -960 241786 480 8 la_oenb[32]
port 452 nsew signal input
rlabel metal2 s 245170 -960 245282 480 8 la_oenb[33]
port 453 nsew signal input
rlabel metal2 s 248758 -960 248870 480 8 la_oenb[34]
port 454 nsew signal input
rlabel metal2 s 252346 -960 252458 480 8 la_oenb[35]
port 455 nsew signal input
rlabel metal2 s 255842 -960 255954 480 8 la_oenb[36]
port 456 nsew signal input
rlabel metal2 s 259430 -960 259542 480 8 la_oenb[37]
port 457 nsew signal input
rlabel metal2 s 262926 -960 263038 480 8 la_oenb[38]
port 458 nsew signal input
rlabel metal2 s 266514 -960 266626 480 8 la_oenb[39]
port 459 nsew signal input
rlabel metal2 s 138818 -960 138930 480 8 la_oenb[3]
port 460 nsew signal input
rlabel metal2 s 270010 -960 270122 480 8 la_oenb[40]
port 461 nsew signal input
rlabel metal2 s 273598 -960 273710 480 8 la_oenb[41]
port 462 nsew signal input
rlabel metal2 s 277094 -960 277206 480 8 la_oenb[42]
port 463 nsew signal input
rlabel metal2 s 280682 -960 280794 480 8 la_oenb[43]
port 464 nsew signal input
rlabel metal2 s 284270 -960 284382 480 8 la_oenb[44]
port 465 nsew signal input
rlabel metal2 s 287766 -960 287878 480 8 la_oenb[45]
port 466 nsew signal input
rlabel metal2 s 291354 -960 291466 480 8 la_oenb[46]
port 467 nsew signal input
rlabel metal2 s 294850 -960 294962 480 8 la_oenb[47]
port 468 nsew signal input
rlabel metal2 s 298438 -960 298550 480 8 la_oenb[48]
port 469 nsew signal input
rlabel metal2 s 301934 -960 302046 480 8 la_oenb[49]
port 470 nsew signal input
rlabel metal2 s 142406 -960 142518 480 8 la_oenb[4]
port 471 nsew signal input
rlabel metal2 s 305522 -960 305634 480 8 la_oenb[50]
port 472 nsew signal input
rlabel metal2 s 309018 -960 309130 480 8 la_oenb[51]
port 473 nsew signal input
rlabel metal2 s 312606 -960 312718 480 8 la_oenb[52]
port 474 nsew signal input
rlabel metal2 s 316194 -960 316306 480 8 la_oenb[53]
port 475 nsew signal input
rlabel metal2 s 319690 -960 319802 480 8 la_oenb[54]
port 476 nsew signal input
rlabel metal2 s 323278 -960 323390 480 8 la_oenb[55]
port 477 nsew signal input
rlabel metal2 s 326774 -960 326886 480 8 la_oenb[56]
port 478 nsew signal input
rlabel metal2 s 330362 -960 330474 480 8 la_oenb[57]
port 479 nsew signal input
rlabel metal2 s 333858 -960 333970 480 8 la_oenb[58]
port 480 nsew signal input
rlabel metal2 s 337446 -960 337558 480 8 la_oenb[59]
port 481 nsew signal input
rlabel metal2 s 145902 -960 146014 480 8 la_oenb[5]
port 482 nsew signal input
rlabel metal2 s 340942 -960 341054 480 8 la_oenb[60]
port 483 nsew signal input
rlabel metal2 s 344530 -960 344642 480 8 la_oenb[61]
port 484 nsew signal input
rlabel metal2 s 348026 -960 348138 480 8 la_oenb[62]
port 485 nsew signal input
rlabel metal2 s 351614 -960 351726 480 8 la_oenb[63]
port 486 nsew signal input
rlabel metal2 s 355202 -960 355314 480 8 la_oenb[64]
port 487 nsew signal input
rlabel metal2 s 358698 -960 358810 480 8 la_oenb[65]
port 488 nsew signal input
rlabel metal2 s 362286 -960 362398 480 8 la_oenb[66]
port 489 nsew signal input
rlabel metal2 s 365782 -960 365894 480 8 la_oenb[67]
port 490 nsew signal input
rlabel metal2 s 369370 -960 369482 480 8 la_oenb[68]
port 491 nsew signal input
rlabel metal2 s 372866 -960 372978 480 8 la_oenb[69]
port 492 nsew signal input
rlabel metal2 s 149490 -960 149602 480 8 la_oenb[6]
port 493 nsew signal input
rlabel metal2 s 376454 -960 376566 480 8 la_oenb[70]
port 494 nsew signal input
rlabel metal2 s 379950 -960 380062 480 8 la_oenb[71]
port 495 nsew signal input
rlabel metal2 s 383538 -960 383650 480 8 la_oenb[72]
port 496 nsew signal input
rlabel metal2 s 387126 -960 387238 480 8 la_oenb[73]
port 497 nsew signal input
rlabel metal2 s 390622 -960 390734 480 8 la_oenb[74]
port 498 nsew signal input
rlabel metal2 s 394210 -960 394322 480 8 la_oenb[75]
port 499 nsew signal input
rlabel metal2 s 397706 -960 397818 480 8 la_oenb[76]
port 500 nsew signal input
rlabel metal2 s 401294 -960 401406 480 8 la_oenb[77]
port 501 nsew signal input
rlabel metal2 s 404790 -960 404902 480 8 la_oenb[78]
port 502 nsew signal input
rlabel metal2 s 408378 -960 408490 480 8 la_oenb[79]
port 503 nsew signal input
rlabel metal2 s 152986 -960 153098 480 8 la_oenb[7]
port 504 nsew signal input
rlabel metal2 s 411874 -960 411986 480 8 la_oenb[80]
port 505 nsew signal input
rlabel metal2 s 415462 -960 415574 480 8 la_oenb[81]
port 506 nsew signal input
rlabel metal2 s 418958 -960 419070 480 8 la_oenb[82]
port 507 nsew signal input
rlabel metal2 s 422546 -960 422658 480 8 la_oenb[83]
port 508 nsew signal input
rlabel metal2 s 426134 -960 426246 480 8 la_oenb[84]
port 509 nsew signal input
rlabel metal2 s 429630 -960 429742 480 8 la_oenb[85]
port 510 nsew signal input
rlabel metal2 s 433218 -960 433330 480 8 la_oenb[86]
port 511 nsew signal input
rlabel metal2 s 436714 -960 436826 480 8 la_oenb[87]
port 512 nsew signal input
rlabel metal2 s 440302 -960 440414 480 8 la_oenb[88]
port 513 nsew signal input
rlabel metal2 s 443798 -960 443910 480 8 la_oenb[89]
port 514 nsew signal input
rlabel metal2 s 156574 -960 156686 480 8 la_oenb[8]
port 515 nsew signal input
rlabel metal2 s 447386 -960 447498 480 8 la_oenb[90]
port 516 nsew signal input
rlabel metal2 s 450882 -960 450994 480 8 la_oenb[91]
port 517 nsew signal input
rlabel metal2 s 454470 -960 454582 480 8 la_oenb[92]
port 518 nsew signal input
rlabel metal2 s 458058 -960 458170 480 8 la_oenb[93]
port 519 nsew signal input
rlabel metal2 s 461554 -960 461666 480 8 la_oenb[94]
port 520 nsew signal input
rlabel metal2 s 465142 -960 465254 480 8 la_oenb[95]
port 521 nsew signal input
rlabel metal2 s 468638 -960 468750 480 8 la_oenb[96]
port 522 nsew signal input
rlabel metal2 s 472226 -960 472338 480 8 la_oenb[97]
port 523 nsew signal input
rlabel metal2 s 475722 -960 475834 480 8 la_oenb[98]
port 524 nsew signal input
rlabel metal2 s 479310 -960 479422 480 8 la_oenb[99]
port 525 nsew signal input
rlabel metal2 s 160070 -960 160182 480 8 la_oenb[9]
port 526 nsew signal input
rlabel metal2 s 579774 -960 579886 480 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 580970 -960 581082 480 8 user_irq[0]
port 528 nsew signal tristate
rlabel metal2 s 582166 -960 582278 480 8 user_irq[1]
port 529 nsew signal tristate
rlabel metal2 s 583362 -960 583474 480 8 user_irq[2]
port 530 nsew signal tristate
rlabel metal5 s -2006 -934 585930 -314 8 vccd1
port 531 nsew power input
rlabel metal5 s -2966 2866 586890 3486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 38866 586890 39486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 74866 586890 75486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 110866 586890 111486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 146866 586890 147486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 182866 586890 183486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 218866 586890 219486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 254866 586890 255486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 290866 586890 291486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 326866 586890 327486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 362866 586890 363486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 398866 586890 399486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 434866 586890 435486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 470866 586890 471486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 506866 586890 507486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 542866 586890 543486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 578866 586890 579486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 614866 586890 615486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 650866 586890 651486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2966 686866 586890 687486 6 vccd1
port 531 nsew power input
rlabel metal5 s -2006 704250 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s -2006 -934 -1386 704870 4 vccd1
port 531 nsew power input
rlabel metal4 s 585310 -934 585930 704870 6 vccd1
port 531 nsew power input
rlabel metal4 s 1794 702000 2414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 37794 702000 38414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 73794 702000 74414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 109794 702000 110414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 145794 702000 146414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 181794 702000 182414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 217794 702000 218414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 253794 702000 254414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 289794 702000 290414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 325794 702000 326414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 361794 702000 362414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 397794 702000 398414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 433794 702000 434414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 469794 702000 470414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 505794 702000 506414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 541794 702000 542414 705830 6 vccd1
port 531 nsew power input
rlabel metal4 s 577794 -1894 578414 705830 6 vccd1
port 531 nsew power input
rlabel metal5 s -3926 -2854 587850 -2234 8 vccd2
port 532 nsew power input
rlabel metal5 s -4886 6586 588810 7206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 42586 588810 43206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 78586 588810 79206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 114586 588810 115206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 150586 588810 151206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 186586 588810 187206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 222586 588810 223206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 258586 588810 259206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 294586 588810 295206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 330586 588810 331206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 366586 588810 367206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 402586 588810 403206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 438586 588810 439206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 474586 588810 475206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 510586 588810 511206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 546586 588810 547206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 582586 588810 583206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 618586 588810 619206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 654586 588810 655206 6 vccd2
port 532 nsew power input
rlabel metal5 s -4886 690586 588810 691206 6 vccd2
port 532 nsew power input
rlabel metal5 s -3926 706170 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 -3814 6134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 41514 -3814 42134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 77514 -3814 78134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 113514 -3814 114134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 149514 -3814 150134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 185514 -3814 186134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 221514 -3814 222134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 257514 -3814 258134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 293514 -3814 294134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 329514 -3814 330134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 365514 -3814 366134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 401514 -3814 402134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 437514 -3814 438134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 473514 -3814 474134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 509514 -3814 510134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s 545514 -3814 546134 -2000 8 vccd2
port 532 nsew power input
rlabel metal4 s -3926 -2854 -3306 706790 4 vccd2
port 532 nsew power input
rlabel metal4 s 587230 -2854 587850 706790 6 vccd2
port 532 nsew power input
rlabel metal4 s 5514 702000 6134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 41514 702000 42134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 77514 702000 78134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 113514 702000 114134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 149514 702000 150134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 185514 702000 186134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 221514 702000 222134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 257514 702000 258134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 293514 702000 294134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 329514 702000 330134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 365514 702000 366134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 401514 702000 402134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 437514 702000 438134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 473514 702000 474134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 509514 702000 510134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 545514 702000 546134 707750 6 vccd2
port 532 nsew power input
rlabel metal4 s 581514 -3814 582134 707750 6 vccd2
port 532 nsew power input
rlabel metal5 s -5846 -4774 589770 -4154 8 vdda1
port 533 nsew power input
rlabel metal5 s -6806 10306 590730 10926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 46306 590730 46926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 82306 590730 82926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 118306 590730 118926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 154306 590730 154926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 190306 590730 190926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 226306 590730 226926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 262306 590730 262926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 298306 590730 298926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 334306 590730 334926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 370306 590730 370926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 406306 590730 406926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 442306 590730 442926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 478306 590730 478926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 514306 590730 514926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 550306 590730 550926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 586306 590730 586926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 622306 590730 622926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 658306 590730 658926 6 vdda1
port 533 nsew power input
rlabel metal5 s -6806 694306 590730 694926 6 vdda1
port 533 nsew power input
rlabel metal5 s -5846 708090 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 -5734 9854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 45234 -5734 45854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 81234 -5734 81854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 117234 -5734 117854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 153234 -5734 153854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 189234 -5734 189854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 225234 -5734 225854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 261234 -5734 261854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 297234 -5734 297854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 333234 -5734 333854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 369234 -5734 369854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 405234 -5734 405854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 441234 -5734 441854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 477234 -5734 477854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 513234 -5734 513854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s 549234 -5734 549854 -2000 8 vdda1
port 533 nsew power input
rlabel metal4 s -5846 -4774 -5226 708710 4 vdda1
port 533 nsew power input
rlabel metal4 s 589150 -4774 589770 708710 6 vdda1
port 533 nsew power input
rlabel metal4 s 9234 702000 9854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 45234 702000 45854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 81234 702000 81854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 117234 702000 117854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 153234 702000 153854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 189234 702000 189854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 225234 702000 225854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 261234 702000 261854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 297234 702000 297854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 333234 702000 333854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 369234 702000 369854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 405234 702000 405854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 441234 702000 441854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 477234 702000 477854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 513234 702000 513854 709670 6 vdda1
port 533 nsew power input
rlabel metal4 s 549234 702000 549854 709670 6 vdda1
port 533 nsew power input
rlabel metal5 s -7766 -6694 591690 -6074 8 vdda2
port 534 nsew power input
rlabel metal5 s -8726 14026 592650 14646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 50026 592650 50646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 86026 592650 86646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 122026 592650 122646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 158026 592650 158646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 194026 592650 194646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 230026 592650 230646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 266026 592650 266646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 302026 592650 302646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 338026 592650 338646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 374026 592650 374646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 410026 592650 410646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 446026 592650 446646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 482026 592650 482646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 518026 592650 518646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 554026 592650 554646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 590026 592650 590646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 626026 592650 626646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 662026 592650 662646 6 vdda2
port 534 nsew power input
rlabel metal5 s -8726 698026 592650 698646 6 vdda2
port 534 nsew power input
rlabel metal5 s -7766 710010 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 -7654 13574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 48954 -7654 49574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 84954 -7654 85574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 120954 -7654 121574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 156954 -7654 157574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 192954 -7654 193574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 228954 -7654 229574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 264954 -7654 265574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 300954 -7654 301574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 336954 -7654 337574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 372954 -7654 373574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 408954 -7654 409574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 444954 -7654 445574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 480954 -7654 481574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 516954 -7654 517574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s 552954 -7654 553574 -2000 8 vdda2
port 534 nsew power input
rlabel metal4 s -7766 -6694 -7146 710630 4 vdda2
port 534 nsew power input
rlabel metal4 s 591070 -6694 591690 710630 6 vdda2
port 534 nsew power input
rlabel metal4 s 12954 702000 13574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 48954 702000 49574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 84954 702000 85574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 120954 702000 121574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 156954 702000 157574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 192954 702000 193574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 228954 702000 229574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 264954 702000 265574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 300954 702000 301574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 336954 702000 337574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 372954 702000 373574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 408954 702000 409574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 444954 702000 445574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 480954 702000 481574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 516954 702000 517574 711590 6 vdda2
port 534 nsew power input
rlabel metal4 s 552954 702000 553574 711590 6 vdda2
port 534 nsew power input
rlabel metal5 s -6806 -5734 590730 -5114 8 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 28306 590730 28926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 64306 590730 64926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 100306 590730 100926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 136306 590730 136926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 172306 590730 172926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 208306 590730 208926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 244306 590730 244926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 280306 590730 280926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 316306 590730 316926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 352306 590730 352926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 388306 590730 388926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 424306 590730 424926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 460306 590730 460926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 496306 590730 496926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 532306 590730 532926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 568306 590730 568926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 604306 590730 604926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 640306 590730 640926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 676306 590730 676926 6 vssa1
port 535 nsew ground input
rlabel metal5 s -6806 709050 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 -5734 27854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 -5734 63854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 -5734 99854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 -5734 135854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 -5734 171854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 -5734 207854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 -5734 243854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 -5734 279854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 -5734 315854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 -5734 351854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 -5734 387854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 -5734 423854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 -5734 459854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 -5734 495854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 -5734 531854 -2000 8 vssa1
port 535 nsew ground input
rlabel metal4 s -6806 -5734 -6186 709670 4 vssa1
port 535 nsew ground input
rlabel metal4 s 27234 702000 27854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 63234 702000 63854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 99234 702000 99854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 135234 702000 135854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 171234 702000 171854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 207234 702000 207854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 243234 702000 243854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 279234 702000 279854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 315234 702000 315854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 351234 702000 351854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 387234 702000 387854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 423234 702000 423854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 459234 702000 459854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 495234 702000 495854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 531234 702000 531854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 567234 -5734 567854 709670 6 vssa1
port 535 nsew ground input
rlabel metal4 s 590110 -5734 590730 709670 6 vssa1
port 535 nsew ground input
rlabel metal5 s -8726 -7654 592650 -7034 8 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 32026 592650 32646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 68026 592650 68646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 104026 592650 104646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 140026 592650 140646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 176026 592650 176646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 212026 592650 212646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 248026 592650 248646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 284026 592650 284646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 320026 592650 320646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 356026 592650 356646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 392026 592650 392646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 428026 592650 428646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 464026 592650 464646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 500026 592650 500646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 536026 592650 536646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 572026 592650 572646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 608026 592650 608646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 644026 592650 644646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 680026 592650 680646 6 vssa2
port 536 nsew ground input
rlabel metal5 s -8726 710970 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 -7654 31574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 -7654 67574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 -7654 103574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 -7654 139574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 -7654 175574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 -7654 211574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 -7654 247574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 -7654 283574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 -7654 319574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 -7654 355574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 -7654 391574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 -7654 427574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 -7654 463574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 -7654 499574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 -7654 535574 -2000 8 vssa2
port 536 nsew ground input
rlabel metal4 s -8726 -7654 -8106 711590 4 vssa2
port 536 nsew ground input
rlabel metal4 s 30954 702000 31574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 66954 702000 67574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 102954 702000 103574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 138954 702000 139574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 174954 702000 175574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 210954 702000 211574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 246954 702000 247574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 282954 702000 283574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 318954 702000 319574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 354954 702000 355574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 390954 702000 391574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 426954 702000 427574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 462954 702000 463574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 498954 702000 499574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 534954 702000 535574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 570954 -7654 571574 711590 6 vssa2
port 536 nsew ground input
rlabel metal4 s 592030 -7654 592650 711590 6 vssa2
port 536 nsew ground input
rlabel metal5 s -2966 -1894 586890 -1274 8 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 20866 586890 21486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 56866 586890 57486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 92866 586890 93486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 128866 586890 129486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 164866 586890 165486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 200866 586890 201486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 236866 586890 237486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 272866 586890 273486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 308866 586890 309486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 344866 586890 345486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 380866 586890 381486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 416866 586890 417486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 452866 586890 453486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 488866 586890 489486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 524866 586890 525486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 560866 586890 561486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 596866 586890 597486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 632866 586890 633486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 668866 586890 669486 6 vssd1
port 537 nsew ground input
rlabel metal5 s -2966 705210 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s -2966 -1894 -2346 705830 4 vssd1
port 537 nsew ground input
rlabel metal4 s 19794 702000 20414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 55794 702000 56414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 91794 702000 92414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 127794 702000 128414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 163794 702000 164414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 199794 702000 200414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 235794 702000 236414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 271794 702000 272414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 307794 702000 308414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 343794 702000 344414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 379794 702000 380414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 415794 702000 416414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 451794 702000 452414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 487794 702000 488414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 523794 702000 524414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 559794 702000 560414 705830 6 vssd1
port 537 nsew ground input
rlabel metal4 s 586270 -1894 586890 705830 6 vssd1
port 537 nsew ground input
rlabel metal5 s -4886 -3814 588810 -3194 8 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 24586 588810 25206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 60586 588810 61206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 96586 588810 97206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 132586 588810 133206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 168586 588810 169206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 204586 588810 205206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 240586 588810 241206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 276586 588810 277206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 312586 588810 313206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 348586 588810 349206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 384586 588810 385206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 420586 588810 421206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 456586 588810 457206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 492586 588810 493206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 528586 588810 529206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 564586 588810 565206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 600586 588810 601206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 636586 588810 637206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 672586 588810 673206 6 vssd2
port 538 nsew ground input
rlabel metal5 s -4886 707130 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 -3814 24134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 -3814 60134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 -3814 96134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 -3814 132134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 -3814 168134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 -3814 204134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 -3814 240134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 -3814 276134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 -3814 312134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 -3814 348134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 -3814 384134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 -3814 420134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 -3814 456134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 -3814 492134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 -3814 528134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 -3814 564134 -2000 8 vssd2
port 538 nsew ground input
rlabel metal4 s -4886 -3814 -4266 707750 4 vssd2
port 538 nsew ground input
rlabel metal4 s 23514 702000 24134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 59514 702000 60134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 95514 702000 96134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 131514 702000 132134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 167514 702000 168134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 203514 702000 204134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 239514 702000 240134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 275514 702000 276134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 311514 702000 312134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 347514 702000 348134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 383514 702000 384134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 419514 702000 420134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 455514 702000 456134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 491514 702000 492134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 527514 702000 528134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 563514 702000 564134 707750 6 vssd2
port 538 nsew ground input
rlabel metal4 s 588190 -3814 588810 707750 6 vssd2
port 538 nsew ground input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 539 nsew signal input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 540 nsew signal input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 541 nsew signal tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 542 nsew signal input
rlabel metal2 s 47830 -960 47942 480 8 wbs_adr_i[10]
port 543 nsew signal input
rlabel metal2 s 51326 -960 51438 480 8 wbs_adr_i[11]
port 544 nsew signal input
rlabel metal2 s 54914 -960 55026 480 8 wbs_adr_i[12]
port 545 nsew signal input
rlabel metal2 s 58410 -960 58522 480 8 wbs_adr_i[13]
port 546 nsew signal input
rlabel metal2 s 61998 -960 62110 480 8 wbs_adr_i[14]
port 547 nsew signal input
rlabel metal2 s 65494 -960 65606 480 8 wbs_adr_i[15]
port 548 nsew signal input
rlabel metal2 s 69082 -960 69194 480 8 wbs_adr_i[16]
port 549 nsew signal input
rlabel metal2 s 72578 -960 72690 480 8 wbs_adr_i[17]
port 550 nsew signal input
rlabel metal2 s 76166 -960 76278 480 8 wbs_adr_i[18]
port 551 nsew signal input
rlabel metal2 s 79662 -960 79774 480 8 wbs_adr_i[19]
port 552 nsew signal input
rlabel metal2 s 12318 -960 12430 480 8 wbs_adr_i[1]
port 553 nsew signal input
rlabel metal2 s 83250 -960 83362 480 8 wbs_adr_i[20]
port 554 nsew signal input
rlabel metal2 s 86838 -960 86950 480 8 wbs_adr_i[21]
port 555 nsew signal input
rlabel metal2 s 90334 -960 90446 480 8 wbs_adr_i[22]
port 556 nsew signal input
rlabel metal2 s 93922 -960 94034 480 8 wbs_adr_i[23]
port 557 nsew signal input
rlabel metal2 s 97418 -960 97530 480 8 wbs_adr_i[24]
port 558 nsew signal input
rlabel metal2 s 101006 -960 101118 480 8 wbs_adr_i[25]
port 559 nsew signal input
rlabel metal2 s 104502 -960 104614 480 8 wbs_adr_i[26]
port 560 nsew signal input
rlabel metal2 s 108090 -960 108202 480 8 wbs_adr_i[27]
port 561 nsew signal input
rlabel metal2 s 111586 -960 111698 480 8 wbs_adr_i[28]
port 562 nsew signal input
rlabel metal2 s 115174 -960 115286 480 8 wbs_adr_i[29]
port 563 nsew signal input
rlabel metal2 s 17010 -960 17122 480 8 wbs_adr_i[2]
port 564 nsew signal input
rlabel metal2 s 118762 -960 118874 480 8 wbs_adr_i[30]
port 565 nsew signal input
rlabel metal2 s 122258 -960 122370 480 8 wbs_adr_i[31]
port 566 nsew signal input
rlabel metal2 s 21794 -960 21906 480 8 wbs_adr_i[3]
port 567 nsew signal input
rlabel metal2 s 26486 -960 26598 480 8 wbs_adr_i[4]
port 568 nsew signal input
rlabel metal2 s 30074 -960 30186 480 8 wbs_adr_i[5]
port 569 nsew signal input
rlabel metal2 s 33570 -960 33682 480 8 wbs_adr_i[6]
port 570 nsew signal input
rlabel metal2 s 37158 -960 37270 480 8 wbs_adr_i[7]
port 571 nsew signal input
rlabel metal2 s 40654 -960 40766 480 8 wbs_adr_i[8]
port 572 nsew signal input
rlabel metal2 s 44242 -960 44354 480 8 wbs_adr_i[9]
port 573 nsew signal input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 574 nsew signal input
rlabel metal2 s 8730 -960 8842 480 8 wbs_dat_i[0]
port 575 nsew signal input
rlabel metal2 s 48934 -960 49046 480 8 wbs_dat_i[10]
port 576 nsew signal input
rlabel metal2 s 52522 -960 52634 480 8 wbs_dat_i[11]
port 577 nsew signal input
rlabel metal2 s 56018 -960 56130 480 8 wbs_dat_i[12]
port 578 nsew signal input
rlabel metal2 s 59606 -960 59718 480 8 wbs_dat_i[13]
port 579 nsew signal input
rlabel metal2 s 63194 -960 63306 480 8 wbs_dat_i[14]
port 580 nsew signal input
rlabel metal2 s 66690 -960 66802 480 8 wbs_dat_i[15]
port 581 nsew signal input
rlabel metal2 s 70278 -960 70390 480 8 wbs_dat_i[16]
port 582 nsew signal input
rlabel metal2 s 73774 -960 73886 480 8 wbs_dat_i[17]
port 583 nsew signal input
rlabel metal2 s 77362 -960 77474 480 8 wbs_dat_i[18]
port 584 nsew signal input
rlabel metal2 s 80858 -960 80970 480 8 wbs_dat_i[19]
port 585 nsew signal input
rlabel metal2 s 13514 -960 13626 480 8 wbs_dat_i[1]
port 586 nsew signal input
rlabel metal2 s 84446 -960 84558 480 8 wbs_dat_i[20]
port 587 nsew signal input
rlabel metal2 s 87942 -960 88054 480 8 wbs_dat_i[21]
port 588 nsew signal input
rlabel metal2 s 91530 -960 91642 480 8 wbs_dat_i[22]
port 589 nsew signal input
rlabel metal2 s 95118 -960 95230 480 8 wbs_dat_i[23]
port 590 nsew signal input
rlabel metal2 s 98614 -960 98726 480 8 wbs_dat_i[24]
port 591 nsew signal input
rlabel metal2 s 102202 -960 102314 480 8 wbs_dat_i[25]
port 592 nsew signal input
rlabel metal2 s 105698 -960 105810 480 8 wbs_dat_i[26]
port 593 nsew signal input
rlabel metal2 s 109286 -960 109398 480 8 wbs_dat_i[27]
port 594 nsew signal input
rlabel metal2 s 112782 -960 112894 480 8 wbs_dat_i[28]
port 595 nsew signal input
rlabel metal2 s 116370 -960 116482 480 8 wbs_dat_i[29]
port 596 nsew signal input
rlabel metal2 s 18206 -960 18318 480 8 wbs_dat_i[2]
port 597 nsew signal input
rlabel metal2 s 119866 -960 119978 480 8 wbs_dat_i[30]
port 598 nsew signal input
rlabel metal2 s 123454 -960 123566 480 8 wbs_dat_i[31]
port 599 nsew signal input
rlabel metal2 s 22990 -960 23102 480 8 wbs_dat_i[3]
port 600 nsew signal input
rlabel metal2 s 27682 -960 27794 480 8 wbs_dat_i[4]
port 601 nsew signal input
rlabel metal2 s 31270 -960 31382 480 8 wbs_dat_i[5]
port 602 nsew signal input
rlabel metal2 s 34766 -960 34878 480 8 wbs_dat_i[6]
port 603 nsew signal input
rlabel metal2 s 38354 -960 38466 480 8 wbs_dat_i[7]
port 604 nsew signal input
rlabel metal2 s 41850 -960 41962 480 8 wbs_dat_i[8]
port 605 nsew signal input
rlabel metal2 s 45438 -960 45550 480 8 wbs_dat_i[9]
port 606 nsew signal input
rlabel metal2 s 9926 -960 10038 480 8 wbs_dat_o[0]
port 607 nsew signal tristate
rlabel metal2 s 50130 -960 50242 480 8 wbs_dat_o[10]
port 608 nsew signal tristate
rlabel metal2 s 53718 -960 53830 480 8 wbs_dat_o[11]
port 609 nsew signal tristate
rlabel metal2 s 57214 -960 57326 480 8 wbs_dat_o[12]
port 610 nsew signal tristate
rlabel metal2 s 60802 -960 60914 480 8 wbs_dat_o[13]
port 611 nsew signal tristate
rlabel metal2 s 64298 -960 64410 480 8 wbs_dat_o[14]
port 612 nsew signal tristate
rlabel metal2 s 67886 -960 67998 480 8 wbs_dat_o[15]
port 613 nsew signal tristate
rlabel metal2 s 71474 -960 71586 480 8 wbs_dat_o[16]
port 614 nsew signal tristate
rlabel metal2 s 74970 -960 75082 480 8 wbs_dat_o[17]
port 615 nsew signal tristate
rlabel metal2 s 78558 -960 78670 480 8 wbs_dat_o[18]
port 616 nsew signal tristate
rlabel metal2 s 82054 -960 82166 480 8 wbs_dat_o[19]
port 617 nsew signal tristate
rlabel metal2 s 14710 -960 14822 480 8 wbs_dat_o[1]
port 618 nsew signal tristate
rlabel metal2 s 85642 -960 85754 480 8 wbs_dat_o[20]
port 619 nsew signal tristate
rlabel metal2 s 89138 -960 89250 480 8 wbs_dat_o[21]
port 620 nsew signal tristate
rlabel metal2 s 92726 -960 92838 480 8 wbs_dat_o[22]
port 621 nsew signal tristate
rlabel metal2 s 96222 -960 96334 480 8 wbs_dat_o[23]
port 622 nsew signal tristate
rlabel metal2 s 99810 -960 99922 480 8 wbs_dat_o[24]
port 623 nsew signal tristate
rlabel metal2 s 103306 -960 103418 480 8 wbs_dat_o[25]
port 624 nsew signal tristate
rlabel metal2 s 106894 -960 107006 480 8 wbs_dat_o[26]
port 625 nsew signal tristate
rlabel metal2 s 110482 -960 110594 480 8 wbs_dat_o[27]
port 626 nsew signal tristate
rlabel metal2 s 113978 -960 114090 480 8 wbs_dat_o[28]
port 627 nsew signal tristate
rlabel metal2 s 117566 -960 117678 480 8 wbs_dat_o[29]
port 628 nsew signal tristate
rlabel metal2 s 19402 -960 19514 480 8 wbs_dat_o[2]
port 629 nsew signal tristate
rlabel metal2 s 121062 -960 121174 480 8 wbs_dat_o[30]
port 630 nsew signal tristate
rlabel metal2 s 124650 -960 124762 480 8 wbs_dat_o[31]
port 631 nsew signal tristate
rlabel metal2 s 24186 -960 24298 480 8 wbs_dat_o[3]
port 632 nsew signal tristate
rlabel metal2 s 28878 -960 28990 480 8 wbs_dat_o[4]
port 633 nsew signal tristate
rlabel metal2 s 32374 -960 32486 480 8 wbs_dat_o[5]
port 634 nsew signal tristate
rlabel metal2 s 35962 -960 36074 480 8 wbs_dat_o[6]
port 635 nsew signal tristate
rlabel metal2 s 39550 -960 39662 480 8 wbs_dat_o[7]
port 636 nsew signal tristate
rlabel metal2 s 43046 -960 43158 480 8 wbs_dat_o[8]
port 637 nsew signal tristate
rlabel metal2 s 46634 -960 46746 480 8 wbs_dat_o[9]
port 638 nsew signal tristate
rlabel metal2 s 11122 -960 11234 480 8 wbs_sel_i[0]
port 639 nsew signal input
rlabel metal2 s 15906 -960 16018 480 8 wbs_sel_i[1]
port 640 nsew signal input
rlabel metal2 s 20598 -960 20710 480 8 wbs_sel_i[2]
port 641 nsew signal input
rlabel metal2 s 25290 -960 25402 480 8 wbs_sel_i[3]
port 642 nsew signal input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 643 nsew signal input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 644 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
